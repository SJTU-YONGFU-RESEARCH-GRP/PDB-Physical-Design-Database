module ibex_core (alert_major_o,
    alert_minor_o,
    clk_i,
    core_sleep_o,
    data_err_i,
    data_gnt_i,
    data_req_o,
    data_rvalid_i,
    data_we_o,
    debug_req_i,
    fetch_enable_i,
    instr_err_i,
    instr_gnt_i,
    instr_req_o,
    instr_rvalid_i,
    irq_external_i,
    irq_nm_i,
    irq_software_i,
    irq_timer_i,
    rst_ni,
    test_en_i,
    boot_addr_i,
    data_addr_o,
    data_be_o,
    data_rdata_i,
    data_wdata_o,
    hart_id_i,
    instr_addr_o,
    instr_rdata_i,
    irq_fast_i);
 output alert_major_o;
 output alert_minor_o;
 input clk_i;
 output core_sleep_o;
 input data_err_i;
 input data_gnt_i;
 output data_req_o;
 input data_rvalid_i;
 output data_we_o;
 input debug_req_i;
 input fetch_enable_i;
 input instr_err_i;
 input instr_gnt_i;
 output instr_req_o;
 input instr_rvalid_i;
 input irq_external_i;
 input irq_nm_i;
 input irq_software_i;
 input irq_timer_i;
 input rst_ni;
 input test_en_i;
 input [31:0] boot_addr_i;
 output [31:0] data_addr_o;
 output [3:0] data_be_o;
 input [31:0] data_rdata_i;
 output [31:0] data_wdata_o;
 input [31:0] hart_id_i;
 output [31:0] instr_addr_o;
 input [31:0] instr_rdata_i;
 input [14:0] irq_fast_i;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire clknet_leaf_23_clk_i_regs;
 wire clknet_leaf_22_clk_i_regs;
 wire clknet_leaf_21_clk_i_regs;
 wire clknet_leaf_20_clk_i_regs;
 wire _01670_;
 wire clknet_leaf_19_clk_i_regs;
 wire _01672_;
 wire clknet_leaf_18_clk_i_regs;
 wire _01674_;
 wire clknet_leaf_17_clk_i_regs;
 wire clknet_leaf_16_clk_i_regs;
 wire clknet_leaf_15_clk_i_regs;
 wire clknet_leaf_14_clk_i_regs;
 wire _01679_;
 wire _01680_;
 wire clknet_leaf_13_clk_i_regs;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire clknet_leaf_12_clk_i_regs;
 wire clknet_leaf_11_clk_i_regs;
 wire _01687_;
 wire _01688_;
 wire clknet_leaf_10_clk_i_regs;
 wire _01690_;
 wire clknet_leaf_9_clk_i_regs;
 wire clknet_leaf_8_clk_i_regs;
 wire _01693_;
 wire clknet_leaf_7_clk_i_regs;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire clknet_leaf_6_clk_i_regs;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire clknet_leaf_5_clk_i_regs;
 wire clknet_leaf_4_clk_i_regs;
 wire clknet_leaf_3_clk_i_regs;
 wire clknet_leaf_2_clk_i_regs;
 wire clknet_leaf_1_clk_i_regs;
 wire clknet_leaf_0_clk_i_regs;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire clknet_1_0__leaf_clk_i;
 wire clknet_0_clk_i;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire net475;
 wire _01719_;
 wire _01720_;
 wire net474;
 wire net473;
 wire net472;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire net471;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire net470;
 wire _01737_;
 wire _01738_;
 wire net469;
 wire net468;
 wire net467;
 wire _01742_;
 wire _01743_;
 wire net466;
 wire net465;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire net464;
 wire _01750_;
 wire _01751_;
 wire net463;
 wire net462;
 wire net461;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire net460;
 wire net459;
 wire _01761_;
 wire _01762_;
 wire net458;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire net457;
 wire _01773_;
 wire net456;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire net455;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire net454;
 wire net453;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire net452;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire net451;
 wire net450;
 wire net449;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire net448;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire net447;
 wire _01847_;
 wire _01848_;
 wire net446;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire net445;
 wire _01882_;
 wire _01883_;
 wire net444;
 wire net443;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire net442;
 wire net441;
 wire _01896_;
 wire net440;
 wire _01898_;
 wire net439;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire net438;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire net437;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire net436;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire net435;
 wire _01921_;
 wire net434;
 wire _01923_;
 wire net433;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire net432;
 wire net431;
 wire net430;
 wire net429;
 wire net428;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire net427;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire net426;
 wire net425;
 wire net424;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire net423;
 wire _01968_;
 wire net422;
 wire _01970_;
 wire net421;
 wire _01972_;
 wire net420;
 wire net419;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire net418;
 wire _01980_;
 wire net417;
 wire _01982_;
 wire net416;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire net415;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire net414;
 wire net413;
 wire net412;
 wire _02002_;
 wire _02003_;
 wire net411;
 wire _02005_;
 wire _02006_;
 wire net410;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire net409;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire net408;
 wire net407;
 wire net406;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire net405;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire net404;
 wire _02032_;
 wire net403;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire net402;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire net401;
 wire net400;
 wire _02061_;
 wire net399;
 wire net398;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire net397;
 wire _02083_;
 wire net396;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire net395;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire net394;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire net393;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire net392;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire net391;
 wire _02125_;
 wire net390;
 wire net389;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire net388;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire net387;
 wire net386;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire net385;
 wire net384;
 wire _02228_;
 wire net383;
 wire net382;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire net381;
 wire net380;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire net379;
 wire _02252_;
 wire _02253_;
 wire net378;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire net377;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire net376;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire net375;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire net374;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire net373;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire net372;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire net371;
 wire net370;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire net369;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire net368;
 wire _02419_;
 wire net367;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire net366;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire net365;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire net364;
 wire _02467_;
 wire _02468_;
 wire net363;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire net362;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire net361;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire net360;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire net359;
 wire net358;
 wire _02516_;
 wire _02517_;
 wire net357;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire net356;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire net355;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire net354;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire net353;
 wire _02621_;
 wire _02622_;
 wire net352;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire net351;
 wire net350;
 wire net349;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire net348;
 wire _02655_;
 wire _02656_;
 wire net347;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire net346;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire net345;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire net344;
 wire _02725_;
 wire net343;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire net342;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire net341;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire net340;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire net339;
 wire net338;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire net337;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire net336;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire net335;
 wire net334;
 wire _02935_;
 wire _02936_;
 wire net333;
 wire net332;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire net331;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire net330;
 wire _03082_;
 wire _03083_;
 wire net329;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire net328;
 wire _03096_;
 wire _03097_;
 wire net327;
 wire _03099_;
 wire _03100_;
 wire net326;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire net325;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire net324;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire net323;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire net322;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire net321;
 wire _03216_;
 wire net320;
 wire _03218_;
 wire net319;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire net318;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire net317;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire net316;
 wire _03312_;
 wire _03313_;
 wire net315;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire net314;
 wire _03350_;
 wire _03351_;
 wire net313;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire net312;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire net311;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire net310;
 wire _03483_;
 wire net309;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire net308;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire net307;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire net306;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire net305;
 wire net304;
 wire _03698_;
 wire _03699_;
 wire net303;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire net302;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire net301;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire net300;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire net299;
 wire _03821_;
 wire net298;
 wire _03823_;
 wire net297;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire net296;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire net295;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire net294;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire net293;
 wire _03933_;
 wire net292;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire net291;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire net290;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire net289;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire net288;
 wire net287;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire net286;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire net285;
 wire net284;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire net283;
 wire _04083_;
 wire net282;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire net281;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire net280;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire net279;
 wire net278;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire net277;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire net276;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire net275;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire net274;
 wire net273;
 wire net272;
 wire net271;
 wire _04344_;
 wire net270;
 wire net269;
 wire net268;
 wire _04348_;
 wire net267;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire net266;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire net265;
 wire _04429_;
 wire net264;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire net263;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire net262;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire net261;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire net260;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire net259;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire net258;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire net257;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire net256;
 wire _04810_;
 wire net255;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire net254;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire net253;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire net252;
 wire net251;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire net250;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire net249;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire net248;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire net247;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire net246;
 wire _05218_;
 wire net245;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire net244;
 wire _05263_;
 wire _05264_;
 wire net243;
 wire _05266_;
 wire net242;
 wire _05268_;
 wire net241;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire net240;
 wire _05274_;
 wire net239;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire net238;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire net237;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire net236;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire net235;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire net234;
 wire _05357_;
 wire _05358_;
 wire net233;
 wire _05360_;
 wire _05361_;
 wire net232;
 wire _05363_;
 wire _05364_;
 wire net231;
 wire _05366_;
 wire _05367_;
 wire net230;
 wire _05369_;
 wire _05370_;
 wire net229;
 wire _05372_;
 wire _05373_;
 wire net228;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire net227;
 wire net226;
 wire _05381_;
 wire net225;
 wire _05383_;
 wire net224;
 wire _05385_;
 wire _05386_;
 wire net223;
 wire _05388_;
 wire _05389_;
 wire net222;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire net221;
 wire _05395_;
 wire _05396_;
 wire net220;
 wire _05398_;
 wire _05399_;
 wire net219;
 wire _05401_;
 wire _05402_;
 wire net218;
 wire _05404_;
 wire _05405_;
 wire net217;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire net216;
 wire _05412_;
 wire _05413_;
 wire net215;
 wire _05415_;
 wire _05416_;
 wire net214;
 wire _05418_;
 wire _05419_;
 wire net213;
 wire _05421_;
 wire _05422_;
 wire net212;
 wire _05424_;
 wire _05425_;
 wire net211;
 wire _05427_;
 wire net210;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire net209;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire net208;
 wire _05439_;
 wire net207;
 wire _05441_;
 wire net206;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire net205;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire net204;
 wire _05465_;
 wire net203;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire net202;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire net201;
 wire _05508_;
 wire net200;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire net199;
 wire _05534_;
 wire net198;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire net197;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire net196;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire net195;
 wire _05574_;
 wire net194;
 wire _05576_;
 wire _05577_;
 wire net193;
 wire _05579_;
 wire net192;
 wire _05581_;
 wire net191;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire net190;
 wire _05604_;
 wire net189;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire net188;
 wire _05642_;
 wire _05643_;
 wire net187;
 wire _05645_;
 wire net186;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire net185;
 wire _05670_;
 wire net184;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire net183;
 wire _05708_;
 wire _05709_;
 wire net182;
 wire _05711_;
 wire net181;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire net180;
 wire _05737_;
 wire net179;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire net178;
 wire _05772_;
 wire _05773_;
 wire net177;
 wire _05775_;
 wire net176;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire net175;
 wire _05795_;
 wire _05796_;
 wire net174;
 wire _05798_;
 wire net173;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire net172;
 wire _05806_;
 wire net171;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire net170;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire net169;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire net168;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire net167;
 wire _05844_;
 wire net166;
 wire net165;
 wire _05847_;
 wire net164;
 wire _05849_;
 wire net163;
 wire net162;
 wire _05852_;
 wire net161;
 wire _05854_;
 wire net160;
 wire _05856_;
 wire net159;
 wire net158;
 wire _05859_;
 wire net157;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire net156;
 wire _05865_;
 wire _05866_;
 wire net155;
 wire _05868_;
 wire net154;
 wire _05870_;
 wire _05871_;
 wire net153;
 wire net152;
 wire _05874_;
 wire _05875_;
 wire net151;
 wire net150;
 wire _05878_;
 wire net149;
 wire net148;
 wire _05881_;
 wire _05882_;
 wire net147;
 wire net146;
 wire net145;
 wire net144;
 wire net143;
 wire net142;
 wire net141;
 wire net140;
 wire net139;
 wire net138;
 wire net137;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire net136;
 wire _05898_;
 wire net135;
 wire net134;
 wire net133;
 wire net132;
 wire net131;
 wire net130;
 wire net129;
 wire net128;
 wire _05907_;
 wire _05908_;
 wire net127;
 wire net126;
 wire _05911_;
 wire net125;
 wire _05913_;
 wire net124;
 wire _05915_;
 wire net123;
 wire net122;
 wire _05918_;
 wire _05919_;
 wire net121;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire net120;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire net119;
 wire net118;
 wire _05935_;
 wire _05936_;
 wire net117;
 wire _05938_;
 wire net116;
 wire _05940_;
 wire net115;
 wire _05942_;
 wire net114;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire net113;
 wire _05950_;
 wire net112;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire net111;
 wire net110;
 wire _05960_;
 wire _05961_;
 wire net109;
 wire _05963_;
 wire _05964_;
 wire net108;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire net107;
 wire net106;
 wire _05978_;
 wire _05979_;
 wire net105;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire net104;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire net103;
 wire net102;
 wire _05994_;
 wire _05995_;
 wire net101;
 wire _05997_;
 wire net100;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire net99;
 wire net98;
 wire _06009_;
 wire _06010_;
 wire net97;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire net96;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire net95;
 wire _06028_;
 wire _06029_;
 wire net94;
 wire _06031_;
 wire net93;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire net92;
 wire _06055_;
 wire net91;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire net90;
 wire _06091_;
 wire _06092_;
 wire net89;
 wire _06094_;
 wire net88;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire net87;
 wire _06114_;
 wire _06115_;
 wire net86;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire net85;
 wire _06123_;
 wire net84;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire net83;
 wire net82;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire net81;
 wire _06163_;
 wire _06164_;
 wire net80;
 wire _06166_;
 wire net79;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire net78;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire net77;
 wire _06191_;
 wire net76;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire net75;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire net74;
 wire _06230_;
 wire net73;
 wire _06232_;
 wire _06233_;
 wire net72;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire net71;
 wire _06239_;
 wire net70;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire net69;
 wire _06264_;
 wire net68;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire net67;
 wire _06302_;
 wire _06303_;
 wire net66;
 wire _06305_;
 wire net65;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire net64;
 wire _06330_;
 wire net63;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire net62;
 wire _06368_;
 wire _06369_;
 wire net61;
 wire _06371_;
 wire net60;
 wire _06373_;
 wire net59;
 wire _06375_;
 wire net58;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire net57;
 wire _06400_;
 wire net56;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire net55;
 wire _06440_;
 wire _06441_;
 wire net54;
 wire _06443_;
 wire net53;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire net52;
 wire _06467_;
 wire net51;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire net50;
 wire _06505_;
 wire _06506_;
 wire net49;
 wire _06508_;
 wire net48;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire net47;
 wire _06533_;
 wire net46;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire net45;
 wire net44;
 wire _06572_;
 wire _06573_;
 wire net43;
 wire _06575_;
 wire net42;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire net41;
 wire net40;
 wire _06587_;
 wire _06588_;
 wire net39;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire net38;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire net37;
 wire net36;
 wire _06606_;
 wire _06607_;
 wire net35;
 wire _06609_;
 wire net34;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire net33;
 wire net32;
 wire _06619_;
 wire _06620_;
 wire net31;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire net30;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire net1142;
 wire net1141;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire net1140;
 wire net1139;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire net1138;
 wire net1137;
 wire net1136;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire net1135;
 wire net1134;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire net1133;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire net1132;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire net1131;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire net1130;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire net1129;
 wire _06757_;
 wire net1128;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire net1127;
 wire net1126;
 wire net1125;
 wire net1124;
 wire _06770_;
 wire net1123;
 wire _06772_;
 wire net1122;
 wire _06774_;
 wire net1121;
 wire _06776_;
 wire net1120;
 wire _06778_;
 wire net1119;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire net1118;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire net1117;
 wire net1116;
 wire _06814_;
 wire net1115;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire net1114;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire net1113;
 wire _06826_;
 wire net1112;
 wire _06828_;
 wire net1111;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire net1110;
 wire net1109;
 wire _06836_;
 wire _06837_;
 wire net1108;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire net1107;
 wire net1106;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire net1105;
 wire _06864_;
 wire _06865_;
 wire net1104;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire net1103;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire net1102;
 wire _06895_;
 wire _06896_;
 wire net1101;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire net1100;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire net1099;
 wire _07029_;
 wire net1098;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire net1097;
 wire net1096;
 wire net1095;
 wire _07284_;
 wire net1094;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire net1093;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire net1092;
 wire net1091;
 wire net1090;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire net1089;
 wire _07346_;
 wire _07347_;
 wire net1088;
 wire _07349_;
 wire net1087;
 wire _07351_;
 wire _07352_;
 wire net1086;
 wire net1085;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire net1084;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire net1083;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire net1082;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire net1081;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire net1080;
 wire _07432_;
 wire _07433_;
 wire net1079;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire net1078;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire net1077;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire net1076;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire net1075;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire net1074;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire net1073;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire net1072;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire net1071;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire net1070;
 wire net1030;
 wire net1029;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire net1016;
 wire _07728_;
 wire _07729_;
 wire net1015;
 wire net1014;
 wire net1013;
 wire _07733_;
 wire net1012;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire net1011;
 wire net1010;
 wire net1009;
 wire _07759_;
 wire _07760_;
 wire net1008;
 wire net1007;
 wire net1006;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire net1005;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire net1004;
 wire _07783_;
 wire net1003;
 wire _07785_;
 wire _07786_;
 wire net1002;
 wire net1001;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire net1000;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire net999;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire net998;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire net997;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire net996;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire net995;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire net994;
 wire _08100_;
 wire net993;
 wire net992;
 wire net991;
 wire _08104_;
 wire net990;
 wire _08106_;
 wire _08107_;
 wire net989;
 wire _08109_;
 wire net988;
 wire _08111_;
 wire net987;
 wire net986;
 wire net985;
 wire net984;
 wire net983;
 wire _08117_;
 wire _08118_;
 wire net982;
 wire net981;
 wire _08121_;
 wire net980;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire net979;
 wire net978;
 wire net977;
 wire net976;
 wire net975;
 wire net974;
 wire net973;
 wire net972;
 wire net971;
 wire net970;
 wire net969;
 wire net968;
 wire _08138_;
 wire _08139_;
 wire net967;
 wire net966;
 wire _08142_;
 wire _08143_;
 wire net965;
 wire net964;
 wire net963;
 wire net962;
 wire net961;
 wire net960;
 wire net959;
 wire net958;
 wire _08152_;
 wire net957;
 wire net956;
 wire net955;
 wire net954;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire net953;
 wire net952;
 wire net951;
 wire net950;
 wire net949;
 wire net948;
 wire net947;
 wire net946;
 wire net945;
 wire net944;
 wire net943;
 wire net942;
 wire net941;
 wire _08179_;
 wire net940;
 wire net939;
 wire net938;
 wire net937;
 wire net936;
 wire net935;
 wire net934;
 wire _08187_;
 wire net933;
 wire net932;
 wire _08190_;
 wire net931;
 wire net930;
 wire net929;
 wire _08194_;
 wire _08195_;
 wire net928;
 wire net927;
 wire net926;
 wire net925;
 wire _08200_;
 wire net924;
 wire _08202_;
 wire net923;
 wire net922;
 wire _08205_;
 wire _08206_;
 wire net921;
 wire _08208_;
 wire net920;
 wire net919;
 wire _08211_;
 wire net918;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire net917;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire net916;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire net915;
 wire net914;
 wire net913;
 wire net912;
 wire _08277_;
 wire net911;
 wire net910;
 wire _08280_;
 wire net909;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire net908;
 wire net907;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire net906;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire net905;
 wire net904;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire net903;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire net902;
 wire _08309_;
 wire net901;
 wire net900;
 wire net899;
 wire net898;
 wire _08314_;
 wire net897;
 wire net896;
 wire _08317_;
 wire net895;
 wire net894;
 wire _08320_;
 wire _08321_;
 wire net893;
 wire _08323_;
 wire _08324_;
 wire net892;
 wire net891;
 wire net890;
 wire _08328_;
 wire net889;
 wire _08330_;
 wire _08331_;
 wire net888;
 wire _08333_;
 wire _08334_;
 wire net887;
 wire net886;
 wire net885;
 wire net884;
 wire _08339_;
 wire net883;
 wire net882;
 wire _08342_;
 wire net881;
 wire _08344_;
 wire net880;
 wire net879;
 wire net878;
 wire net877;
 wire _08349_;
 wire _08350_;
 wire net876;
 wire net875;
 wire _08353_;
 wire net874;
 wire net873;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire net872;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire net871;
 wire _08370_;
 wire net870;
 wire _08372_;
 wire net869;
 wire _08374_;
 wire _08375_;
 wire net868;
 wire _08377_;
 wire net867;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire net866;
 wire _08431_;
 wire net865;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire net864;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire net863;
 wire net862;
 wire _08453_;
 wire net861;
 wire net860;
 wire _08456_;
 wire _08457_;
 wire net859;
 wire net858;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire net857;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire net856;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire net855;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire net854;
 wire _08497_;
 wire _08498_;
 wire net853;
 wire _08500_;
 wire net852;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire net851;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire net850;
 wire _08512_;
 wire net849;
 wire net848;
 wire _08515_;
 wire net847;
 wire net846;
 wire _08518_;
 wire net845;
 wire _08520_;
 wire net844;
 wire _08522_;
 wire net843;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire net842;
 wire net841;
 wire _08529_;
 wire net840;
 wire _08531_;
 wire _08532_;
 wire net839;
 wire _08534_;
 wire net838;
 wire _08536_;
 wire net837;
 wire net836;
 wire _08539_;
 wire net835;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire net834;
 wire net833;
 wire _08554_;
 wire net832;
 wire net831;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire net830;
 wire _08561_;
 wire net829;
 wire _08563_;
 wire _08564_;
 wire net828;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire net827;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire net826;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire net825;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire net824;
 wire _08592_;
 wire _08593_;
 wire net823;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire net822;
 wire net821;
 wire _08605_;
 wire _08606_;
 wire net820;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire net819;
 wire _08612_;
 wire _08613_;
 wire net818;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire net817;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire net816;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire net815;
 wire _08646_;
 wire _08647_;
 wire net814;
 wire net813;
 wire net812;
 wire net811;
 wire net810;
 wire net809;
 wire net808;
 wire net807;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire net806;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire net805;
 wire net804;
 wire net803;
 wire _08666_;
 wire net802;
 wire net801;
 wire _08669_;
 wire _08670_;
 wire net800;
 wire net799;
 wire _08673_;
 wire net798;
 wire _08675_;
 wire net797;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire net796;
 wire net795;
 wire net794;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire net793;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire net792;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire net791;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire net790;
 wire net789;
 wire _08716_;
 wire net788;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire net787;
 wire _08723_;
 wire _08724_;
 wire net786;
 wire _08726_;
 wire _08727_;
 wire net785;
 wire net784;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire net783;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire net782;
 wire _08745_;
 wire _08746_;
 wire net781;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire net780;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire net779;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire net778;
 wire net777;
 wire net776;
 wire _08769_;
 wire _08770_;
 wire net775;
 wire _08772_;
 wire _08773_;
 wire net774;
 wire net773;
 wire _08776_;
 wire net772;
 wire _08778_;
 wire net771;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire net770;
 wire net769;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire net768;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire net767;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire net766;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire net765;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire net764;
 wire _08823_;
 wire _08824_;
 wire net763;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire net762;
 wire net761;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire net760;
 wire net759;
 wire net758;
 wire net757;
 wire _08861_;
 wire net756;
 wire net755;
 wire _08864_;
 wire _08865_;
 wire net754;
 wire _08867_;
 wire net753;
 wire net752;
 wire _08870_;
 wire net751;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire net750;
 wire net749;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire net748;
 wire _08900_;
 wire _08901_;
 wire net747;
 wire net746;
 wire net745;
 wire net744;
 wire _08906_;
 wire _08907_;
 wire net743;
 wire _08909_;
 wire _08910_;
 wire net742;
 wire _08912_;
 wire _08913_;
 wire net741;
 wire _08915_;
 wire _08916_;
 wire net740;
 wire net739;
 wire net738;
 wire _08920_;
 wire net737;
 wire net736;
 wire _08923_;
 wire _08924_;
 wire net735;
 wire _08926_;
 wire net734;
 wire net733;
 wire net732;
 wire net731;
 wire _08931_;
 wire _08932_;
 wire net730;
 wire net729;
 wire _08935_;
 wire net728;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire net727;
 wire net726;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire net725;
 wire net724;
 wire _08970_;
 wire net723;
 wire net722;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire net721;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire net1576;
 wire net719;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire net1577;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire net717;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire net716;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire net715;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire net714;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire net713;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire net712;
 wire _09132_;
 wire _09133_;
 wire net711;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire net710;
 wire _09142_;
 wire net709;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire net708;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire net707;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire net706;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire net705;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire net704;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire net703;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire net702;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire net701;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire net700;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire net699;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire net698;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire net697;
 wire net696;
 wire _09455_;
 wire net695;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire net694;
 wire _09494_;
 wire net693;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire net692;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire net691;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire net690;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire net689;
 wire _09579_;
 wire net688;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire net687;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire net686;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire net685;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire net684;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire net683;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire net682;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire net681;
 wire _09828_;
 wire _09829_;
 wire net680;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire net679;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire net678;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire net677;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire net676;
 wire net675;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire net674;
 wire net673;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire net672;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire net671;
 wire net670;
 wire net669;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire net668;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire net667;
 wire net666;
 wire _10133_;
 wire net665;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire net664;
 wire net663;
 wire net662;
 wire _10141_;
 wire _10142_;
 wire net661;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire net660;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire net659;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire net658;
 wire _10175_;
 wire _10176_;
 wire net657;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire net656;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire net655;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire net654;
 wire net653;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire net652;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire net1578;
 wire _10499_;
 wire _10500_;
 wire net650;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire net649;
 wire _10564_;
 wire _10565_;
 wire net648;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire net647;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire net646;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire net645;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire net644;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire net643;
 wire net642;
 wire net641;
 wire net640;
 wire _10815_;
 wire net639;
 wire net638;
 wire net637;
 wire net636;
 wire _10820_;
 wire net635;
 wire net634;
 wire _10823_;
 wire _10824_;
 wire net633;
 wire _10826_;
 wire net632;
 wire net631;
 wire net630;
 wire net629;
 wire net628;
 wire net627;
 wire net626;
 wire net625;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire net623;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire net622;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire net621;
 wire _10854_;
 wire net620;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire net619;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire net618;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire net617;
 wire _10917_;
 wire _10918_;
 wire net616;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire net615;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire net614;
 wire net613;
 wire net612;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire net611;
 wire net610;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire net609;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire net608;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire net607;
 wire _11042_;
 wire _11043_;
 wire net606;
 wire net605;
 wire net604;
 wire net603;
 wire net602;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire net601;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire net599;
 wire _11061_;
 wire net598;
 wire net597;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire net595;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire net590;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire net585;
 wire net583;
 wire _11118_;
 wire net582;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire net581;
 wire net580;
 wire net579;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire net578;
 wire _11146_;
 wire net577;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire net576;
 wire net575;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire net574;
 wire _11206_;
 wire _11207_;
 wire net573;
 wire _11209_;
 wire net572;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire net571;
 wire net570;
 wire _11217_;
 wire _11218_;
 wire net569;
 wire net568;
 wire net567;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire net566;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire net565;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire net564;
 wire _11251_;
 wire _11252_;
 wire net563;
 wire _11254_;
 wire _11255_;
 wire net562;
 wire net561;
 wire net560;
 wire _11259_;
 wire _11260_;
 wire net559;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire net558;
 wire _11266_;
 wire _11267_;
 wire net557;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire net556;
 wire _11279_;
 wire _11280_;
 wire net555;
 wire _11282_;
 wire net554;
 wire net553;
 wire net552;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire net551;
 wire _11290_;
 wire net550;
 wire net549;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire net548;
 wire net547;
 wire net546;
 wire _11299_;
 wire net545;
 wire net544;
 wire _11302_;
 wire net543;
 wire net542;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire net541;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire net540;
 wire _11316_;
 wire net539;
 wire net538;
 wire net537;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire net536;
 wire _11324_;
 wire _11325_;
 wire net535;
 wire net534;
 wire _11328_;
 wire net533;
 wire _11330_;
 wire _11331_;
 wire net532;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire net531;
 wire net530;
 wire net529;
 wire net528;
 wire net527;
 wire _11345_;
 wire _11346_;
 wire net526;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire net525;
 wire net524;
 wire _11353_;
 wire _11354_;
 wire net523;
 wire _11356_;
 wire _11357_;
 wire net522;
 wire net521;
 wire _11360_;
 wire net520;
 wire net519;
 wire net518;
 wire net517;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire net516;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire net515;
 wire net514;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire net513;
 wire _11386_;
 wire net512;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire net511;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire net510;
 wire _11400_;
 wire _11401_;
 wire net509;
 wire _11403_;
 wire net508;
 wire net507;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire net506;
 wire _11418_;
 wire net505;
 wire net504;
 wire _11421_;
 wire _11422_;
 wire net503;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire net502;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire net501;
 wire net500;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire net499;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire net498;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire net497;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire net496;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire net495;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire net494;
 wire net493;
 wire _11475_;
 wire _11476_;
 wire net492;
 wire net491;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire net490;
 wire _11507_;
 wire net489;
 wire _11509_;
 wire _11510_;
 wire net488;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire net487;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire net486;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire net485;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire net484;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire net483;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire net482;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire net481;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire net480;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire net479;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire net1474;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire net477;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire net476;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire delaynet_1_core_clock;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire delaynet_0_core_clock;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire clknet_3_7_0_clk;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire clknet_3_6_0_clk;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire clknet_3_5_0_clk;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire clknet_3_4_0_clk;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire clknet_3_3_0_clk;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire clknet_3_2_0_clk;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire clknet_3_1_0_clk;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire clknet_3_0_0_clk;
 wire _11835_;
 wire clknet_0_clk;
 wire clknet_leaf_81_clk;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire clknet_leaf_80_clk;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire clknet_leaf_79_clk;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire clknet_leaf_78_clk;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire clknet_leaf_77_clk;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire clknet_leaf_76_clk;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire clknet_leaf_75_clk;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire clknet_leaf_74_clk;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire clknet_leaf_73_clk;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire clknet_leaf_72_clk;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_70_clk;
 wire _12143_;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_68_clk;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire clknet_leaf_67_clk;
 wire _12158_;
 wire clknet_leaf_66_clk;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire clknet_leaf_65_clk;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire clknet_leaf_64_clk;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire clknet_leaf_63_clk;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire clknet_leaf_62_clk;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire clknet_leaf_61_clk;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_58_clk;
 wire _12252_;
 wire clknet_leaf_57_clk;
 wire _12254_;
 wire _12255_;
 wire clknet_leaf_56_clk;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire clknet_leaf_55_clk;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire clknet_leaf_54_clk;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire clknet_leaf_53_clk;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire clknet_leaf_52_clk;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire clknet_leaf_51_clk;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire clknet_leaf_50_clk;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_48_clk;
 wire _12455_;
 wire clknet_leaf_47_clk;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_45_clk;
 wire _12462_;
 wire _12463_;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_43_clk;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire clknet_leaf_42_clk;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire clknet_leaf_41_clk;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_39_clk;
 wire _12497_;
 wire _12498_;
 wire clknet_leaf_38_clk;
 wire _12500_;
 wire _12501_;
 wire clknet_leaf_37_clk;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire clknet_leaf_36_clk;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire clknet_leaf_35_clk;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire clknet_leaf_34_clk;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_31_clk;
 wire _12538_;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_29_clk;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire clknet_leaf_28_clk;
 wire _12553_;
 wire _12554_;
 wire clknet_leaf_27_clk;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire clknet_leaf_26_clk;
 wire _12573_;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_24_clk;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_22_clk;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire clknet_leaf_21_clk;
 wire _12622_;
 wire clknet_leaf_20_clk;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire clknet_leaf_19_clk;
 wire _12634_;
 wire clknet_leaf_18_clk;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_16_clk;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire clknet_leaf_15_clk;
 wire _12660_;
 wire clknet_leaf_14_clk;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire clknet_leaf_13_clk;
 wire _12672_;
 wire clknet_leaf_12_clk;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire clknet_leaf_11_clk;
 wire _12687_;
 wire _12688_;
 wire clknet_leaf_10_clk;
 wire _12690_;
 wire clknet_leaf_9_clk;
 wire _12692_;
 wire clknet_leaf_8_clk;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_6_clk;
 wire _12721_;
 wire clknet_leaf_5_clk;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire clknet_leaf_4_clk;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire clknet_leaf_3_clk;
 wire _12760_;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_1_clk;
 wire _12763_;
 wire _12764_;
 wire clknet_leaf_0_clk;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire clknet_3_7__leaf_clk_i_regs;
 wire _12771_;
 wire clknet_3_6__leaf_clk_i_regs;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire clknet_3_5__leaf_clk_i_regs;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire clknet_3_4__leaf_clk_i_regs;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire clknet_3_3__leaf_clk_i_regs;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire clknet_3_2__leaf_clk_i_regs;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire clknet_3_1__leaf_clk_i_regs;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire clknet_3_0__leaf_clk_i_regs;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire clknet_0_clk_i_regs;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire clknet_leaf_99_clk_i_regs;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire clknet_leaf_98_clk_i_regs;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire clknet_leaf_97_clk_i_regs;
 wire clknet_leaf_96_clk_i_regs;
 wire _12893_;
 wire _12894_;
 wire clknet_leaf_95_clk_i_regs;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire clknet_leaf_94_clk_i_regs;
 wire clknet_leaf_93_clk_i_regs;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire clknet_leaf_92_clk_i_regs;
 wire _12925_;
 wire clknet_leaf_91_clk_i_regs;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire clknet_leaf_90_clk_i_regs;
 wire _12937_;
 wire clknet_leaf_89_clk_i_regs;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire clknet_leaf_88_clk_i_regs;
 wire clknet_leaf_87_clk_i_regs;
 wire clknet_leaf_86_clk_i_regs;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire clknet_leaf_85_clk_i_regs;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire clknet_leaf_84_clk_i_regs;
 wire _12976_;
 wire _12977_;
 wire clknet_leaf_83_clk_i_regs;
 wire _12979_;
 wire clknet_leaf_82_clk_i_regs;
 wire _12981_;
 wire _12982_;
 wire clknet_leaf_81_clk_i_regs;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire clknet_leaf_80_clk_i_regs;
 wire clknet_leaf_79_clk_i_regs;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire clknet_leaf_78_clk_i_regs;
 wire _13000_;
 wire clknet_leaf_77_clk_i_regs;
 wire _13002_;
 wire _13003_;
 wire clknet_leaf_76_clk_i_regs;
 wire clknet_leaf_75_clk_i_regs;
 wire clknet_leaf_74_clk_i_regs;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire clknet_leaf_73_clk_i_regs;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire clknet_leaf_72_clk_i_regs;
 wire clknet_leaf_71_clk_i_regs;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire clknet_leaf_70_clk_i_regs;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire clknet_leaf_69_clk_i_regs;
 wire clknet_leaf_68_clk_i_regs;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire clknet_leaf_67_clk_i_regs;
 wire _13090_;
 wire _13091_;
 wire clknet_leaf_66_clk_i_regs;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire clknet_leaf_65_clk_i_regs;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire clknet_leaf_64_clk_i_regs;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire clknet_leaf_63_clk_i_regs;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire clknet_leaf_62_clk_i_regs;
 wire clknet_leaf_61_clk_i_regs;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire clknet_leaf_60_clk_i_regs;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire clknet_leaf_59_clk_i_regs;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire clknet_leaf_58_clk_i_regs;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire clknet_leaf_57_clk_i_regs;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire clknet_leaf_56_clk_i_regs;
 wire clknet_leaf_55_clk_i_regs;
 wire clknet_leaf_54_clk_i_regs;
 wire _13255_;
 wire clknet_leaf_53_clk_i_regs;
 wire _13257_;
 wire clknet_leaf_52_clk_i_regs;
 wire clknet_leaf_51_clk_i_regs;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire clknet_leaf_50_clk_i_regs;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire clknet_leaf_49_clk_i_regs;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire clknet_leaf_48_clk_i_regs;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire clknet_leaf_47_clk_i_regs;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire clknet_leaf_46_clk_i_regs;
 wire _13337_;
 wire _13338_;
 wire clknet_leaf_45_clk_i_regs;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire clknet_leaf_44_clk_i_regs;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire clknet_leaf_43_clk_i_regs;
 wire clknet_leaf_42_clk_i_regs;
 wire _13357_;
 wire _13358_;
 wire clknet_leaf_41_clk_i_regs;
 wire clknet_leaf_40_clk_i_regs;
 wire _13361_;
 wire _13362_;
 wire clknet_leaf_39_clk_i_regs;
 wire clknet_leaf_38_clk_i_regs;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire clknet_leaf_37_clk_i_regs;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire clknet_leaf_36_clk_i_regs;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire clknet_leaf_35_clk_i_regs;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire clknet_leaf_34_clk_i_regs;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire clknet_leaf_33_clk_i_regs;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire clknet_leaf_32_clk_i_regs;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire clknet_leaf_31_clk_i_regs;
 wire _13423_;
 wire _13424_;
 wire clknet_leaf_30_clk_i_regs;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire clknet_leaf_29_clk_i_regs;
 wire _13472_;
 wire clknet_leaf_28_clk_i_regs;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire clknet_leaf_27_clk_i_regs;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire clknet_leaf_26_clk_i_regs;
 wire _13490_;
 wire clknet_leaf_25_clk_i_regs;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire clknet_leaf_24_clk_i_regs;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire net29;
 wire clk_i_regs;
 wire net20;
 wire net19;
 wire net18;
 wire net17;
 wire net16;
 wire net15;
 wire net14;
 wire net13;
 wire net12;
 wire net11;
 wire net10;
 wire net9;
 wire net8;
 wire net7;
 wire net6;
 wire net5;
 wire net4;
 wire net3;
 wire net2;
 wire net1;
 wire net28;
 wire net27;
 wire net26;
 wire net25;
 wire net24;
 wire net23;
 wire net22;
 wire net21;
 wire clk;
 wire core_busy_d;
 wire core_busy_q;
 wire \core_clock_gate_i.en_latch ;
 wire \cs_registers_i.csr_depc_o[10] ;
 wire \cs_registers_i.csr_depc_o[11] ;
 wire \cs_registers_i.csr_depc_o[12] ;
 wire \cs_registers_i.csr_depc_o[13] ;
 wire \cs_registers_i.csr_depc_o[14] ;
 wire \cs_registers_i.csr_depc_o[15] ;
 wire \cs_registers_i.csr_depc_o[16] ;
 wire \cs_registers_i.csr_depc_o[17] ;
 wire \cs_registers_i.csr_depc_o[18] ;
 wire \cs_registers_i.csr_depc_o[19] ;
 wire \cs_registers_i.csr_depc_o[1] ;
 wire \cs_registers_i.csr_depc_o[20] ;
 wire \cs_registers_i.csr_depc_o[21] ;
 wire \cs_registers_i.csr_depc_o[22] ;
 wire \cs_registers_i.csr_depc_o[23] ;
 wire \cs_registers_i.csr_depc_o[24] ;
 wire \cs_registers_i.csr_depc_o[25] ;
 wire \cs_registers_i.csr_depc_o[26] ;
 wire \cs_registers_i.csr_depc_o[27] ;
 wire \cs_registers_i.csr_depc_o[28] ;
 wire \cs_registers_i.csr_depc_o[29] ;
 wire \cs_registers_i.csr_depc_o[2] ;
 wire \cs_registers_i.csr_depc_o[30] ;
 wire \cs_registers_i.csr_depc_o[31] ;
 wire \cs_registers_i.csr_depc_o[3] ;
 wire \cs_registers_i.csr_depc_o[4] ;
 wire \cs_registers_i.csr_depc_o[5] ;
 wire \cs_registers_i.csr_depc_o[6] ;
 wire \cs_registers_i.csr_depc_o[7] ;
 wire \cs_registers_i.csr_depc_o[8] ;
 wire \cs_registers_i.csr_depc_o[9] ;
 wire \cs_registers_i.csr_mepc_o[0] ;
 wire \cs_registers_i.csr_mepc_o[10] ;
 wire \cs_registers_i.csr_mepc_o[11] ;
 wire \cs_registers_i.csr_mepc_o[12] ;
 wire \cs_registers_i.csr_mepc_o[13] ;
 wire \cs_registers_i.csr_mepc_o[14] ;
 wire \cs_registers_i.csr_mepc_o[15] ;
 wire \cs_registers_i.csr_mepc_o[16] ;
 wire \cs_registers_i.csr_mepc_o[17] ;
 wire \cs_registers_i.csr_mepc_o[18] ;
 wire \cs_registers_i.csr_mepc_o[19] ;
 wire \cs_registers_i.csr_mepc_o[1] ;
 wire \cs_registers_i.csr_mepc_o[20] ;
 wire \cs_registers_i.csr_mepc_o[21] ;
 wire \cs_registers_i.csr_mepc_o[22] ;
 wire \cs_registers_i.csr_mepc_o[23] ;
 wire \cs_registers_i.csr_mepc_o[24] ;
 wire \cs_registers_i.csr_mepc_o[25] ;
 wire \cs_registers_i.csr_mepc_o[26] ;
 wire \cs_registers_i.csr_mepc_o[27] ;
 wire \cs_registers_i.csr_mepc_o[28] ;
 wire \cs_registers_i.csr_mepc_o[29] ;
 wire \cs_registers_i.csr_mepc_o[2] ;
 wire \cs_registers_i.csr_mepc_o[30] ;
 wire \cs_registers_i.csr_mepc_o[31] ;
 wire \cs_registers_i.csr_mepc_o[3] ;
 wire \cs_registers_i.csr_mepc_o[4] ;
 wire \cs_registers_i.csr_mepc_o[5] ;
 wire \cs_registers_i.csr_mepc_o[6] ;
 wire \cs_registers_i.csr_mepc_o[7] ;
 wire \cs_registers_i.csr_mepc_o[8] ;
 wire \cs_registers_i.csr_mepc_o[9] ;
 wire \cs_registers_i.csr_mstatus_mie_o ;
 wire \cs_registers_i.csr_mstatus_tw_o ;
 wire \cs_registers_i.csr_mtvec_o[10] ;
 wire \cs_registers_i.csr_mtvec_o[11] ;
 wire \cs_registers_i.csr_mtvec_o[12] ;
 wire \cs_registers_i.csr_mtvec_o[13] ;
 wire \cs_registers_i.csr_mtvec_o[14] ;
 wire \cs_registers_i.csr_mtvec_o[15] ;
 wire \cs_registers_i.csr_mtvec_o[16] ;
 wire \cs_registers_i.csr_mtvec_o[17] ;
 wire \cs_registers_i.csr_mtvec_o[18] ;
 wire \cs_registers_i.csr_mtvec_o[19] ;
 wire \cs_registers_i.csr_mtvec_o[20] ;
 wire \cs_registers_i.csr_mtvec_o[21] ;
 wire \cs_registers_i.csr_mtvec_o[22] ;
 wire \cs_registers_i.csr_mtvec_o[23] ;
 wire \cs_registers_i.csr_mtvec_o[24] ;
 wire \cs_registers_i.csr_mtvec_o[25] ;
 wire \cs_registers_i.csr_mtvec_o[26] ;
 wire \cs_registers_i.csr_mtvec_o[27] ;
 wire \cs_registers_i.csr_mtvec_o[28] ;
 wire \cs_registers_i.csr_mtvec_o[29] ;
 wire \cs_registers_i.csr_mtvec_o[30] ;
 wire \cs_registers_i.csr_mtvec_o[31] ;
 wire \cs_registers_i.csr_mtvec_o[8] ;
 wire \cs_registers_i.csr_mtvec_o[9] ;
 wire \cs_registers_i.dcsr_q[0] ;
 wire \cs_registers_i.dcsr_q[11] ;
 wire \cs_registers_i.dcsr_q[12] ;
 wire \cs_registers_i.dcsr_q[13] ;
 wire \cs_registers_i.dcsr_q[15] ;
 wire \cs_registers_i.dcsr_q[1] ;
 wire \cs_registers_i.dcsr_q[2] ;
 wire \cs_registers_i.dcsr_q[6] ;
 wire \cs_registers_i.dcsr_q[7] ;
 wire \cs_registers_i.dcsr_q[8] ;
 wire \cs_registers_i.debug_mode_i ;
 wire \cs_registers_i.dscratch0_q[0] ;
 wire \cs_registers_i.dscratch0_q[10] ;
 wire \cs_registers_i.dscratch0_q[11] ;
 wire \cs_registers_i.dscratch0_q[12] ;
 wire \cs_registers_i.dscratch0_q[13] ;
 wire \cs_registers_i.dscratch0_q[14] ;
 wire \cs_registers_i.dscratch0_q[15] ;
 wire \cs_registers_i.dscratch0_q[16] ;
 wire \cs_registers_i.dscratch0_q[17] ;
 wire \cs_registers_i.dscratch0_q[18] ;
 wire \cs_registers_i.dscratch0_q[19] ;
 wire \cs_registers_i.dscratch0_q[1] ;
 wire \cs_registers_i.dscratch0_q[20] ;
 wire \cs_registers_i.dscratch0_q[21] ;
 wire \cs_registers_i.dscratch0_q[22] ;
 wire \cs_registers_i.dscratch0_q[23] ;
 wire \cs_registers_i.dscratch0_q[24] ;
 wire \cs_registers_i.dscratch0_q[25] ;
 wire \cs_registers_i.dscratch0_q[26] ;
 wire \cs_registers_i.dscratch0_q[27] ;
 wire \cs_registers_i.dscratch0_q[28] ;
 wire \cs_registers_i.dscratch0_q[29] ;
 wire \cs_registers_i.dscratch0_q[2] ;
 wire \cs_registers_i.dscratch0_q[30] ;
 wire \cs_registers_i.dscratch0_q[31] ;
 wire \cs_registers_i.dscratch0_q[3] ;
 wire \cs_registers_i.dscratch0_q[4] ;
 wire \cs_registers_i.dscratch0_q[5] ;
 wire \cs_registers_i.dscratch0_q[6] ;
 wire \cs_registers_i.dscratch0_q[7] ;
 wire \cs_registers_i.dscratch0_q[8] ;
 wire \cs_registers_i.dscratch0_q[9] ;
 wire \cs_registers_i.dscratch1_q[0] ;
 wire \cs_registers_i.dscratch1_q[10] ;
 wire \cs_registers_i.dscratch1_q[11] ;
 wire \cs_registers_i.dscratch1_q[12] ;
 wire \cs_registers_i.dscratch1_q[13] ;
 wire \cs_registers_i.dscratch1_q[14] ;
 wire \cs_registers_i.dscratch1_q[15] ;
 wire \cs_registers_i.dscratch1_q[16] ;
 wire \cs_registers_i.dscratch1_q[17] ;
 wire \cs_registers_i.dscratch1_q[18] ;
 wire \cs_registers_i.dscratch1_q[19] ;
 wire \cs_registers_i.dscratch1_q[1] ;
 wire \cs_registers_i.dscratch1_q[20] ;
 wire \cs_registers_i.dscratch1_q[21] ;
 wire \cs_registers_i.dscratch1_q[22] ;
 wire \cs_registers_i.dscratch1_q[23] ;
 wire \cs_registers_i.dscratch1_q[24] ;
 wire \cs_registers_i.dscratch1_q[25] ;
 wire \cs_registers_i.dscratch1_q[26] ;
 wire \cs_registers_i.dscratch1_q[27] ;
 wire \cs_registers_i.dscratch1_q[28] ;
 wire \cs_registers_i.dscratch1_q[29] ;
 wire \cs_registers_i.dscratch1_q[2] ;
 wire \cs_registers_i.dscratch1_q[30] ;
 wire \cs_registers_i.dscratch1_q[31] ;
 wire \cs_registers_i.dscratch1_q[3] ;
 wire \cs_registers_i.dscratch1_q[4] ;
 wire \cs_registers_i.dscratch1_q[5] ;
 wire \cs_registers_i.dscratch1_q[6] ;
 wire \cs_registers_i.dscratch1_q[7] ;
 wire \cs_registers_i.dscratch1_q[8] ;
 wire \cs_registers_i.dscratch1_q[9] ;
 wire \cs_registers_i.mcause_q[0] ;
 wire \cs_registers_i.mcause_q[1] ;
 wire \cs_registers_i.mcause_q[2] ;
 wire \cs_registers_i.mcause_q[3] ;
 wire \cs_registers_i.mcause_q[4] ;
 wire \cs_registers_i.mcause_q[5] ;
 wire \cs_registers_i.mcountinhibit[0] ;
 wire \cs_registers_i.mcountinhibit[2] ;
 wire \cs_registers_i.mcycle_counter_i.counter[0] ;
 wire \cs_registers_i.mcycle_counter_i.counter[10] ;
 wire \cs_registers_i.mcycle_counter_i.counter[11] ;
 wire \cs_registers_i.mcycle_counter_i.counter[12] ;
 wire \cs_registers_i.mcycle_counter_i.counter[13] ;
 wire \cs_registers_i.mcycle_counter_i.counter[14] ;
 wire \cs_registers_i.mcycle_counter_i.counter[15] ;
 wire \cs_registers_i.mcycle_counter_i.counter[16] ;
 wire \cs_registers_i.mcycle_counter_i.counter[17] ;
 wire \cs_registers_i.mcycle_counter_i.counter[18] ;
 wire \cs_registers_i.mcycle_counter_i.counter[19] ;
 wire \cs_registers_i.mcycle_counter_i.counter[1] ;
 wire \cs_registers_i.mcycle_counter_i.counter[20] ;
 wire \cs_registers_i.mcycle_counter_i.counter[21] ;
 wire \cs_registers_i.mcycle_counter_i.counter[22] ;
 wire \cs_registers_i.mcycle_counter_i.counter[23] ;
 wire \cs_registers_i.mcycle_counter_i.counter[24] ;
 wire \cs_registers_i.mcycle_counter_i.counter[25] ;
 wire \cs_registers_i.mcycle_counter_i.counter[26] ;
 wire \cs_registers_i.mcycle_counter_i.counter[27] ;
 wire \cs_registers_i.mcycle_counter_i.counter[28] ;
 wire \cs_registers_i.mcycle_counter_i.counter[29] ;
 wire \cs_registers_i.mcycle_counter_i.counter[2] ;
 wire \cs_registers_i.mcycle_counter_i.counter[30] ;
 wire \cs_registers_i.mcycle_counter_i.counter[31] ;
 wire \cs_registers_i.mcycle_counter_i.counter[32] ;
 wire \cs_registers_i.mcycle_counter_i.counter[33] ;
 wire \cs_registers_i.mcycle_counter_i.counter[34] ;
 wire \cs_registers_i.mcycle_counter_i.counter[35] ;
 wire \cs_registers_i.mcycle_counter_i.counter[36] ;
 wire \cs_registers_i.mcycle_counter_i.counter[37] ;
 wire \cs_registers_i.mcycle_counter_i.counter[38] ;
 wire \cs_registers_i.mcycle_counter_i.counter[39] ;
 wire \cs_registers_i.mcycle_counter_i.counter[3] ;
 wire \cs_registers_i.mcycle_counter_i.counter[40] ;
 wire \cs_registers_i.mcycle_counter_i.counter[41] ;
 wire \cs_registers_i.mcycle_counter_i.counter[42] ;
 wire \cs_registers_i.mcycle_counter_i.counter[43] ;
 wire \cs_registers_i.mcycle_counter_i.counter[44] ;
 wire \cs_registers_i.mcycle_counter_i.counter[45] ;
 wire \cs_registers_i.mcycle_counter_i.counter[46] ;
 wire \cs_registers_i.mcycle_counter_i.counter[47] ;
 wire \cs_registers_i.mcycle_counter_i.counter[48] ;
 wire \cs_registers_i.mcycle_counter_i.counter[49] ;
 wire \cs_registers_i.mcycle_counter_i.counter[4] ;
 wire \cs_registers_i.mcycle_counter_i.counter[50] ;
 wire \cs_registers_i.mcycle_counter_i.counter[51] ;
 wire \cs_registers_i.mcycle_counter_i.counter[52] ;
 wire \cs_registers_i.mcycle_counter_i.counter[53] ;
 wire \cs_registers_i.mcycle_counter_i.counter[54] ;
 wire \cs_registers_i.mcycle_counter_i.counter[55] ;
 wire \cs_registers_i.mcycle_counter_i.counter[56] ;
 wire \cs_registers_i.mcycle_counter_i.counter[57] ;
 wire \cs_registers_i.mcycle_counter_i.counter[58] ;
 wire \cs_registers_i.mcycle_counter_i.counter[59] ;
 wire \cs_registers_i.mcycle_counter_i.counter[5] ;
 wire \cs_registers_i.mcycle_counter_i.counter[60] ;
 wire \cs_registers_i.mcycle_counter_i.counter[61] ;
 wire \cs_registers_i.mcycle_counter_i.counter[62] ;
 wire \cs_registers_i.mcycle_counter_i.counter[63] ;
 wire \cs_registers_i.mcycle_counter_i.counter[6] ;
 wire \cs_registers_i.mcycle_counter_i.counter[7] ;
 wire \cs_registers_i.mcycle_counter_i.counter[8] ;
 wire \cs_registers_i.mcycle_counter_i.counter[9] ;
 wire \cs_registers_i.mhpmcounter[2][0] ;
 wire \cs_registers_i.mhpmcounter[2][10] ;
 wire \cs_registers_i.mhpmcounter[2][11] ;
 wire \cs_registers_i.mhpmcounter[2][12] ;
 wire \cs_registers_i.mhpmcounter[2][13] ;
 wire \cs_registers_i.mhpmcounter[2][14] ;
 wire \cs_registers_i.mhpmcounter[2][15] ;
 wire \cs_registers_i.mhpmcounter[2][16] ;
 wire \cs_registers_i.mhpmcounter[2][17] ;
 wire \cs_registers_i.mhpmcounter[2][18] ;
 wire \cs_registers_i.mhpmcounter[2][19] ;
 wire \cs_registers_i.mhpmcounter[2][1] ;
 wire \cs_registers_i.mhpmcounter[2][20] ;
 wire \cs_registers_i.mhpmcounter[2][21] ;
 wire \cs_registers_i.mhpmcounter[2][22] ;
 wire \cs_registers_i.mhpmcounter[2][23] ;
 wire \cs_registers_i.mhpmcounter[2][24] ;
 wire \cs_registers_i.mhpmcounter[2][25] ;
 wire \cs_registers_i.mhpmcounter[2][26] ;
 wire \cs_registers_i.mhpmcounter[2][27] ;
 wire \cs_registers_i.mhpmcounter[2][28] ;
 wire \cs_registers_i.mhpmcounter[2][29] ;
 wire \cs_registers_i.mhpmcounter[2][2] ;
 wire \cs_registers_i.mhpmcounter[2][30] ;
 wire \cs_registers_i.mhpmcounter[2][31] ;
 wire \cs_registers_i.mhpmcounter[2][32] ;
 wire \cs_registers_i.mhpmcounter[2][33] ;
 wire \cs_registers_i.mhpmcounter[2][34] ;
 wire \cs_registers_i.mhpmcounter[2][35] ;
 wire \cs_registers_i.mhpmcounter[2][36] ;
 wire \cs_registers_i.mhpmcounter[2][37] ;
 wire \cs_registers_i.mhpmcounter[2][38] ;
 wire \cs_registers_i.mhpmcounter[2][39] ;
 wire \cs_registers_i.mhpmcounter[2][3] ;
 wire \cs_registers_i.mhpmcounter[2][40] ;
 wire \cs_registers_i.mhpmcounter[2][41] ;
 wire \cs_registers_i.mhpmcounter[2][42] ;
 wire \cs_registers_i.mhpmcounter[2][43] ;
 wire \cs_registers_i.mhpmcounter[2][44] ;
 wire \cs_registers_i.mhpmcounter[2][45] ;
 wire \cs_registers_i.mhpmcounter[2][46] ;
 wire \cs_registers_i.mhpmcounter[2][47] ;
 wire \cs_registers_i.mhpmcounter[2][48] ;
 wire \cs_registers_i.mhpmcounter[2][49] ;
 wire \cs_registers_i.mhpmcounter[2][4] ;
 wire \cs_registers_i.mhpmcounter[2][50] ;
 wire \cs_registers_i.mhpmcounter[2][51] ;
 wire \cs_registers_i.mhpmcounter[2][52] ;
 wire \cs_registers_i.mhpmcounter[2][53] ;
 wire \cs_registers_i.mhpmcounter[2][54] ;
 wire \cs_registers_i.mhpmcounter[2][55] ;
 wire \cs_registers_i.mhpmcounter[2][56] ;
 wire \cs_registers_i.mhpmcounter[2][57] ;
 wire \cs_registers_i.mhpmcounter[2][58] ;
 wire \cs_registers_i.mhpmcounter[2][59] ;
 wire \cs_registers_i.mhpmcounter[2][5] ;
 wire \cs_registers_i.mhpmcounter[2][60] ;
 wire \cs_registers_i.mhpmcounter[2][61] ;
 wire \cs_registers_i.mhpmcounter[2][62] ;
 wire \cs_registers_i.mhpmcounter[2][63] ;
 wire \cs_registers_i.mhpmcounter[2][6] ;
 wire \cs_registers_i.mhpmcounter[2][7] ;
 wire \cs_registers_i.mhpmcounter[2][8] ;
 wire \cs_registers_i.mhpmcounter[2][9] ;
 wire \cs_registers_i.mie_q[0] ;
 wire \cs_registers_i.mie_q[10] ;
 wire \cs_registers_i.mie_q[11] ;
 wire \cs_registers_i.mie_q[12] ;
 wire \cs_registers_i.mie_q[13] ;
 wire \cs_registers_i.mie_q[14] ;
 wire \cs_registers_i.mie_q[15] ;
 wire \cs_registers_i.mie_q[16] ;
 wire \cs_registers_i.mie_q[17] ;
 wire \cs_registers_i.mie_q[1] ;
 wire \cs_registers_i.mie_q[2] ;
 wire \cs_registers_i.mie_q[3] ;
 wire \cs_registers_i.mie_q[4] ;
 wire \cs_registers_i.mie_q[5] ;
 wire \cs_registers_i.mie_q[6] ;
 wire \cs_registers_i.mie_q[7] ;
 wire \cs_registers_i.mie_q[8] ;
 wire \cs_registers_i.mie_q[9] ;
 wire \cs_registers_i.mscratch_q[0] ;
 wire \cs_registers_i.mscratch_q[10] ;
 wire \cs_registers_i.mscratch_q[11] ;
 wire \cs_registers_i.mscratch_q[12] ;
 wire \cs_registers_i.mscratch_q[13] ;
 wire \cs_registers_i.mscratch_q[14] ;
 wire \cs_registers_i.mscratch_q[15] ;
 wire \cs_registers_i.mscratch_q[16] ;
 wire \cs_registers_i.mscratch_q[17] ;
 wire \cs_registers_i.mscratch_q[18] ;
 wire \cs_registers_i.mscratch_q[19] ;
 wire \cs_registers_i.mscratch_q[1] ;
 wire \cs_registers_i.mscratch_q[20] ;
 wire \cs_registers_i.mscratch_q[21] ;
 wire \cs_registers_i.mscratch_q[22] ;
 wire \cs_registers_i.mscratch_q[23] ;
 wire \cs_registers_i.mscratch_q[24] ;
 wire \cs_registers_i.mscratch_q[25] ;
 wire \cs_registers_i.mscratch_q[26] ;
 wire \cs_registers_i.mscratch_q[27] ;
 wire \cs_registers_i.mscratch_q[28] ;
 wire \cs_registers_i.mscratch_q[29] ;
 wire \cs_registers_i.mscratch_q[2] ;
 wire \cs_registers_i.mscratch_q[30] ;
 wire \cs_registers_i.mscratch_q[31] ;
 wire \cs_registers_i.mscratch_q[3] ;
 wire \cs_registers_i.mscratch_q[4] ;
 wire \cs_registers_i.mscratch_q[5] ;
 wire \cs_registers_i.mscratch_q[6] ;
 wire \cs_registers_i.mscratch_q[7] ;
 wire \cs_registers_i.mscratch_q[8] ;
 wire \cs_registers_i.mscratch_q[9] ;
 wire \cs_registers_i.mstack_cause_q[0] ;
 wire \cs_registers_i.mstack_cause_q[1] ;
 wire \cs_registers_i.mstack_cause_q[2] ;
 wire \cs_registers_i.mstack_cause_q[3] ;
 wire \cs_registers_i.mstack_cause_q[4] ;
 wire \cs_registers_i.mstack_cause_q[5] ;
 wire \cs_registers_i.mstack_d[0] ;
 wire \cs_registers_i.mstack_d[1] ;
 wire \cs_registers_i.mstack_d[2] ;
 wire \cs_registers_i.mstack_epc_q[0] ;
 wire \cs_registers_i.mstack_epc_q[10] ;
 wire \cs_registers_i.mstack_epc_q[11] ;
 wire \cs_registers_i.mstack_epc_q[12] ;
 wire \cs_registers_i.mstack_epc_q[13] ;
 wire \cs_registers_i.mstack_epc_q[14] ;
 wire \cs_registers_i.mstack_epc_q[15] ;
 wire \cs_registers_i.mstack_epc_q[16] ;
 wire \cs_registers_i.mstack_epc_q[17] ;
 wire \cs_registers_i.mstack_epc_q[18] ;
 wire \cs_registers_i.mstack_epc_q[19] ;
 wire \cs_registers_i.mstack_epc_q[1] ;
 wire \cs_registers_i.mstack_epc_q[20] ;
 wire \cs_registers_i.mstack_epc_q[21] ;
 wire \cs_registers_i.mstack_epc_q[22] ;
 wire \cs_registers_i.mstack_epc_q[23] ;
 wire \cs_registers_i.mstack_epc_q[24] ;
 wire \cs_registers_i.mstack_epc_q[25] ;
 wire \cs_registers_i.mstack_epc_q[26] ;
 wire \cs_registers_i.mstack_epc_q[27] ;
 wire \cs_registers_i.mstack_epc_q[28] ;
 wire \cs_registers_i.mstack_epc_q[29] ;
 wire \cs_registers_i.mstack_epc_q[2] ;
 wire \cs_registers_i.mstack_epc_q[30] ;
 wire \cs_registers_i.mstack_epc_q[31] ;
 wire \cs_registers_i.mstack_epc_q[3] ;
 wire \cs_registers_i.mstack_epc_q[4] ;
 wire \cs_registers_i.mstack_epc_q[5] ;
 wire \cs_registers_i.mstack_epc_q[6] ;
 wire \cs_registers_i.mstack_epc_q[7] ;
 wire \cs_registers_i.mstack_epc_q[8] ;
 wire \cs_registers_i.mstack_epc_q[9] ;
 wire \cs_registers_i.mstack_q[0] ;
 wire \cs_registers_i.mstack_q[1] ;
 wire \cs_registers_i.mstack_q[2] ;
 wire \cs_registers_i.mstatus_q[1] ;
 wire \cs_registers_i.mtval_q[0] ;
 wire \cs_registers_i.mtval_q[10] ;
 wire \cs_registers_i.mtval_q[11] ;
 wire \cs_registers_i.mtval_q[12] ;
 wire \cs_registers_i.mtval_q[13] ;
 wire \cs_registers_i.mtval_q[14] ;
 wire \cs_registers_i.mtval_q[15] ;
 wire \cs_registers_i.mtval_q[16] ;
 wire \cs_registers_i.mtval_q[17] ;
 wire \cs_registers_i.mtval_q[18] ;
 wire \cs_registers_i.mtval_q[19] ;
 wire \cs_registers_i.mtval_q[1] ;
 wire \cs_registers_i.mtval_q[20] ;
 wire \cs_registers_i.mtval_q[21] ;
 wire \cs_registers_i.mtval_q[22] ;
 wire \cs_registers_i.mtval_q[23] ;
 wire \cs_registers_i.mtval_q[24] ;
 wire \cs_registers_i.mtval_q[25] ;
 wire \cs_registers_i.mtval_q[26] ;
 wire \cs_registers_i.mtval_q[27] ;
 wire \cs_registers_i.mtval_q[28] ;
 wire \cs_registers_i.mtval_q[29] ;
 wire \cs_registers_i.mtval_q[2] ;
 wire \cs_registers_i.mtval_q[30] ;
 wire \cs_registers_i.mtval_q[31] ;
 wire \cs_registers_i.mtval_q[3] ;
 wire \cs_registers_i.mtval_q[4] ;
 wire \cs_registers_i.mtval_q[5] ;
 wire \cs_registers_i.mtval_q[6] ;
 wire \cs_registers_i.mtval_q[7] ;
 wire \cs_registers_i.mtval_q[8] ;
 wire \cs_registers_i.mtval_q[9] ;
 wire \cs_registers_i.nmi_mode_i ;
 wire \cs_registers_i.pc_id_i[10] ;
 wire \cs_registers_i.pc_id_i[11] ;
 wire \cs_registers_i.pc_id_i[12] ;
 wire \cs_registers_i.pc_id_i[13] ;
 wire \cs_registers_i.pc_id_i[14] ;
 wire \cs_registers_i.pc_id_i[15] ;
 wire \cs_registers_i.pc_id_i[16] ;
 wire \cs_registers_i.pc_id_i[17] ;
 wire \cs_registers_i.pc_id_i[18] ;
 wire \cs_registers_i.pc_id_i[19] ;
 wire \cs_registers_i.pc_id_i[1] ;
 wire \cs_registers_i.pc_id_i[20] ;
 wire \cs_registers_i.pc_id_i[21] ;
 wire \cs_registers_i.pc_id_i[22] ;
 wire \cs_registers_i.pc_id_i[23] ;
 wire \cs_registers_i.pc_id_i[24] ;
 wire \cs_registers_i.pc_id_i[25] ;
 wire \cs_registers_i.pc_id_i[26] ;
 wire \cs_registers_i.pc_id_i[27] ;
 wire \cs_registers_i.pc_id_i[28] ;
 wire \cs_registers_i.pc_id_i[29] ;
 wire \cs_registers_i.pc_id_i[2] ;
 wire \cs_registers_i.pc_id_i[30] ;
 wire \cs_registers_i.pc_id_i[31] ;
 wire \cs_registers_i.pc_id_i[3] ;
 wire \cs_registers_i.pc_id_i[4] ;
 wire \cs_registers_i.pc_id_i[5] ;
 wire \cs_registers_i.pc_id_i[6] ;
 wire \cs_registers_i.pc_id_i[7] ;
 wire \cs_registers_i.pc_id_i[8] ;
 wire \cs_registers_i.pc_id_i[9] ;
 wire \cs_registers_i.pc_if_i[10] ;
 wire \cs_registers_i.pc_if_i[11] ;
 wire \cs_registers_i.pc_if_i[12] ;
 wire \cs_registers_i.pc_if_i[13] ;
 wire \cs_registers_i.pc_if_i[14] ;
 wire \cs_registers_i.pc_if_i[15] ;
 wire \cs_registers_i.pc_if_i[16] ;
 wire \cs_registers_i.pc_if_i[17] ;
 wire \cs_registers_i.pc_if_i[18] ;
 wire \cs_registers_i.pc_if_i[19] ;
 wire \cs_registers_i.pc_if_i[1] ;
 wire \cs_registers_i.pc_if_i[20] ;
 wire \cs_registers_i.pc_if_i[21] ;
 wire \cs_registers_i.pc_if_i[22] ;
 wire \cs_registers_i.pc_if_i[23] ;
 wire \cs_registers_i.pc_if_i[24] ;
 wire \cs_registers_i.pc_if_i[25] ;
 wire \cs_registers_i.pc_if_i[26] ;
 wire \cs_registers_i.pc_if_i[27] ;
 wire \cs_registers_i.pc_if_i[28] ;
 wire \cs_registers_i.pc_if_i[29] ;
 wire \cs_registers_i.pc_if_i[2] ;
 wire \cs_registers_i.pc_if_i[30] ;
 wire \cs_registers_i.pc_if_i[31] ;
 wire \cs_registers_i.pc_if_i[3] ;
 wire \cs_registers_i.pc_if_i[4] ;
 wire \cs_registers_i.pc_if_i[5] ;
 wire \cs_registers_i.pc_if_i[6] ;
 wire \cs_registers_i.pc_if_i[7] ;
 wire \cs_registers_i.pc_if_i[8] ;
 wire \cs_registers_i.pc_if_i[9] ;
 wire \cs_registers_i.priv_lvl_q[0] ;
 wire \cs_registers_i.priv_lvl_q[1] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[0] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[10] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[11] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[12] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[13] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[14] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[15] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[16] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[17] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[18] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[19] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[1] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[20] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[21] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[22] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[23] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[24] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[25] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[26] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[27] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[28] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[29] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[2] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[30] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[31] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[32] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[33] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[34] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[35] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[36] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[37] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[38] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[39] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[3] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[40] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[41] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[42] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[43] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[44] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[45] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[46] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[47] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[48] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[49] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[4] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[50] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[51] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[52] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[53] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[54] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[55] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[56] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[57] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[58] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[59] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[5] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[60] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[61] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[62] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[63] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[6] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[7] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[8] ;
 wire \ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[9] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_by_zero_q ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[3] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[4] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_valid ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[0] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[2] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[0] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[10] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[11] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[12] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[13] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[14] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[15] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[16] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[17] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[18] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[19] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[1] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[20] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[21] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[22] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[23] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[24] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[25] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[26] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[27] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[28] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[29] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[2] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[30] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[3] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[4] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[5] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[6] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[7] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[8] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[9] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[0] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[10] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[11] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[12] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[13] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[14] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[15] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[16] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[17] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[18] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[19] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[1] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[20] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[21] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[22] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[23] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[24] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[25] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[26] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[27] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[28] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[29] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[2] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[30] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[31] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[3] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[4] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[5] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[6] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[7] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[8] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ;
 wire fetch_enable_q;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[0] ;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[1] ;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[2] ;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[3] ;
 wire \gen_regfile_ff.register_file_i.raddr_a_i[4] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[0] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[1] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[2] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[3] ;
 wire \gen_regfile_ff.register_file_i.raddr_b_i[4] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1000] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1001] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1002] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1003] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1004] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1005] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1006] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1007] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1008] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1009] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[100] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1010] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1011] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1012] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1013] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1014] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1015] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1016] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1017] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1018] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1019] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[101] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1020] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1021] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1022] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[1023] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[102] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[103] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[104] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[105] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[106] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[107] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[108] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[109] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[110] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[111] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[112] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[113] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[114] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[115] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[116] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[117] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[118] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[119] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[120] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[121] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[122] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[123] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[124] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[125] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[126] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[127] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[128] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[129] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[130] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[131] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[132] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[133] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[134] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[135] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[136] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[137] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[138] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[139] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[140] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[141] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[142] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[143] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[144] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[145] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[146] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[147] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[148] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[149] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[150] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[151] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[152] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[153] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[154] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[155] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[156] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[157] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[158] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[159] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[160] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[161] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[162] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[163] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[164] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[165] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[166] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[167] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[168] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[169] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[170] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[171] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[172] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[173] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[174] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[175] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[176] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[177] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[178] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[179] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[180] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[181] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[182] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[183] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[184] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[185] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[186] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[187] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[188] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[189] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[190] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[191] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[192] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[193] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[194] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[195] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[196] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[197] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[198] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[199] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[200] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[201] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[202] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[203] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[204] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[205] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[206] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[207] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[208] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[209] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[210] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[211] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[212] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[213] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[214] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[215] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[216] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[217] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[218] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[219] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[220] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[221] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[222] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[223] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[224] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[225] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[226] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[227] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[228] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[229] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[230] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[231] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[232] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[233] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[234] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[235] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[236] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[237] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[238] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[239] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[240] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[241] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[242] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[243] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[244] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[245] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[246] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[247] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[248] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[249] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[250] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[251] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[252] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[253] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[254] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[255] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[256] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[257] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[258] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[259] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[260] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[261] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[262] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[263] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[264] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[265] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[266] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[267] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[268] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[269] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[270] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[271] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[272] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[273] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[274] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[275] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[276] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[277] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[278] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[279] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[280] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[281] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[282] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[283] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[284] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[285] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[286] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[287] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[288] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[289] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[290] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[291] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[292] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[293] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[294] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[295] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[296] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[297] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[298] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[299] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[300] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[301] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[302] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[303] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[304] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[305] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[306] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[307] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[308] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[309] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[310] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[311] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[312] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[313] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[314] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[315] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[316] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[317] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[318] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[319] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[320] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[321] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[322] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[323] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[324] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[325] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[326] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[327] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[328] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[329] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[32] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[330] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[331] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[332] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[333] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[334] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[335] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[336] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[337] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[338] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[339] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[33] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[340] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[341] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[342] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[343] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[344] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[345] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[346] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[347] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[348] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[349] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[34] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[350] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[351] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[352] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[353] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[354] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[355] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[356] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[357] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[358] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[359] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[35] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[360] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[361] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[362] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[363] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[364] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[365] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[366] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[367] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[368] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[369] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[36] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[370] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[371] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[372] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[373] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[374] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[375] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[376] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[377] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[378] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[379] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[37] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[380] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[381] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[382] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[383] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[384] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[385] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[386] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[387] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[388] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[389] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[38] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[390] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[391] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[392] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[393] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[394] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[395] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[396] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[397] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[398] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[399] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[39] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[400] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[401] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[402] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[403] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[404] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[405] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[406] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[407] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[408] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[409] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[40] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[410] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[411] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[412] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[413] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[414] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[415] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[416] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[417] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[418] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[419] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[41] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[420] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[421] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[422] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[423] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[424] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[425] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[426] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[427] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[428] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[429] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[42] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[430] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[431] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[432] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[433] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[434] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[435] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[436] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[437] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[438] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[439] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[43] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[440] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[441] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[442] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[443] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[444] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[445] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[446] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[447] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[448] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[449] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[44] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[450] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[451] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[452] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[453] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[454] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[455] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[456] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[457] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[458] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[459] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[45] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[460] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[461] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[462] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[463] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[464] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[465] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[466] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[467] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[468] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[469] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[46] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[470] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[471] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[472] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[473] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[474] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[475] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[476] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[477] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[478] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[479] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[47] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[480] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[481] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[482] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[483] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[484] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[485] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[486] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[487] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[488] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[489] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[48] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[490] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[491] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[492] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[493] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[494] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[495] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[496] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[497] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[498] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[499] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[49] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[500] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[501] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[502] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[503] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[504] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[505] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[506] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[507] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[508] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[509] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[50] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[510] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[511] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[512] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[513] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[514] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[515] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[516] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[517] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[518] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[519] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[51] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[520] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[521] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[522] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[523] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[524] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[525] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[526] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[527] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[528] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[529] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[52] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[530] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[531] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[532] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[533] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[534] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[535] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[536] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[537] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[538] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[539] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[53] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[540] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[541] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[542] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[543] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[544] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[545] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[546] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[547] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[548] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[549] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[54] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[550] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[551] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[552] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[553] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[554] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[555] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[556] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[557] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[558] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[559] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[55] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[560] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[561] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[562] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[563] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[564] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[565] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[566] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[567] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[568] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[569] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[56] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[570] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[571] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[572] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[573] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[574] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[575] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[576] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[577] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[578] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[579] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[57] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[580] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[581] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[582] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[583] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[584] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[585] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[586] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[587] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[588] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[589] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[58] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[590] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[591] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[592] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[593] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[594] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[595] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[596] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[597] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[598] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[599] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[59] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[600] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[601] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[602] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[603] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[604] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[605] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[606] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[607] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[608] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[609] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[60] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[610] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[611] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[612] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[613] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[614] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[615] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[616] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[617] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[618] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[619] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[61] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[620] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[621] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[622] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[623] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[624] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[625] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[626] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[627] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[628] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[629] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[62] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[630] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[631] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[632] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[633] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[634] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[635] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[636] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[637] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[638] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[639] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[63] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[640] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[641] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[642] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[643] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[644] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[645] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[646] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[647] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[648] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[649] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[64] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[650] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[651] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[652] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[653] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[654] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[655] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[656] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[657] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[658] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[659] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[65] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[660] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[661] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[662] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[663] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[664] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[665] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[666] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[667] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[668] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[669] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[66] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[670] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[671] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[672] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[673] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[674] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[675] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[676] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[677] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[678] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[679] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[67] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[680] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[681] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[682] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[683] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[684] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[685] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[686] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[687] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[688] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[689] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[68] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[690] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[691] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[692] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[693] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[694] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[695] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[696] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[697] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[698] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[699] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[69] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[700] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[701] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[702] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[703] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[704] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[705] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[706] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[707] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[708] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[709] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[70] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[710] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[711] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[712] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[713] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[714] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[715] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[716] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[717] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[718] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[719] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[71] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[720] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[721] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[722] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[723] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[724] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[725] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[726] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[727] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[728] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[729] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[72] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[730] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[731] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[732] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[733] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[734] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[735] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[736] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[737] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[738] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[739] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[73] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[740] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[741] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[742] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[743] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[744] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[745] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[746] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[747] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[748] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[749] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[74] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[750] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[751] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[752] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[753] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[754] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[755] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[756] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[757] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[758] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[759] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[75] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[760] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[761] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[762] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[763] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[764] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[765] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[766] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[767] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[768] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[769] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[76] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[770] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[771] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[772] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[773] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[774] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[775] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[776] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[777] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[778] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[779] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[77] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[780] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[781] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[782] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[783] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[784] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[785] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[786] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[787] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[788] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[789] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[78] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[790] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[791] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[792] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[793] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[794] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[795] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[796] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[797] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[798] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[799] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[79] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[800] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[801] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[802] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[803] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[804] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[805] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[806] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[807] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[808] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[809] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[80] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[810] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[811] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[812] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[813] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[814] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[815] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[816] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[817] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[818] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[819] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[81] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[820] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[821] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[822] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[823] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[824] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[825] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[826] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[827] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[828] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[829] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[82] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[830] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[831] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[832] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[833] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[834] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[835] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[836] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[837] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[838] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[839] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[83] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[840] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[841] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[842] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[843] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[844] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[845] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[846] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[847] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[848] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[849] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[84] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[850] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[851] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[852] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[853] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[854] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[855] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[856] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[857] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[858] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[859] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[85] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[860] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[861] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[862] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[863] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[864] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[865] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[866] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[867] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[868] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[869] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[86] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[870] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[871] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[872] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[873] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[874] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[875] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[876] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[877] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[878] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[879] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[87] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[880] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[881] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[882] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[883] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[884] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[885] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[886] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[887] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[888] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[889] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[88] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[890] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[891] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[892] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[893] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[894] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[895] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[896] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[897] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[898] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[899] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[89] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[900] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[901] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[902] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[903] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[904] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[905] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[906] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[907] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[908] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[909] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[90] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[910] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[911] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[912] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[913] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[914] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[915] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[916] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[917] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[918] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[919] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[91] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[920] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[921] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[922] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[923] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[924] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[925] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[926] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[927] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[928] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[929] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[92] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[930] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[931] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[932] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[933] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[934] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[935] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[936] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[937] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[938] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[939] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[93] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[940] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[941] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[942] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[943] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[944] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[945] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[946] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[947] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[948] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[949] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[94] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[950] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[951] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[952] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[953] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[954] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[955] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[956] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[957] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[958] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[959] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[95] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[960] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[961] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[962] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[963] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[964] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[965] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[966] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[967] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[968] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[969] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[96] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[970] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[971] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[972] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[973] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[974] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[975] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[976] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[977] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[978] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[979] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[97] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[980] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[981] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[982] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[983] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[984] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[985] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[986] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[987] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[988] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[989] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[98] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[990] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[991] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[992] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[993] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[994] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[995] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[996] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[997] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[998] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[999] ;
 wire \gen_regfile_ff.register_file_i.rf_reg[99] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[0] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[1] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[2] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[3] ;
 wire \gen_regfile_ff.register_file_i.waddr_a_i[4] ;
 wire \id_stage_i.branch_set ;
 wire \id_stage_i.branch_set_d ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs[0] ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs[1] ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs[2] ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs[3] ;
 wire \id_stage_i.controller_i.exc_req_d ;
 wire \id_stage_i.controller_i.exc_req_q ;
 wire \id_stage_i.controller_i.illegal_insn_d ;
 wire \id_stage_i.controller_i.illegal_insn_q ;
 wire \id_stage_i.controller_i.instr_compressed_i[0] ;
 wire \id_stage_i.controller_i.instr_compressed_i[10] ;
 wire \id_stage_i.controller_i.instr_compressed_i[11] ;
 wire \id_stage_i.controller_i.instr_compressed_i[12] ;
 wire \id_stage_i.controller_i.instr_compressed_i[13] ;
 wire \id_stage_i.controller_i.instr_compressed_i[14] ;
 wire \id_stage_i.controller_i.instr_compressed_i[15] ;
 wire \id_stage_i.controller_i.instr_compressed_i[1] ;
 wire \id_stage_i.controller_i.instr_compressed_i[2] ;
 wire \id_stage_i.controller_i.instr_compressed_i[3] ;
 wire \id_stage_i.controller_i.instr_compressed_i[4] ;
 wire \id_stage_i.controller_i.instr_compressed_i[5] ;
 wire \id_stage_i.controller_i.instr_compressed_i[6] ;
 wire \id_stage_i.controller_i.instr_compressed_i[7] ;
 wire \id_stage_i.controller_i.instr_compressed_i[8] ;
 wire \id_stage_i.controller_i.instr_compressed_i[9] ;
 wire \id_stage_i.controller_i.instr_fetch_err_i ;
 wire \id_stage_i.controller_i.instr_fetch_err_plus2_i ;
 wire \id_stage_i.controller_i.instr_i[0] ;
 wire \id_stage_i.controller_i.instr_i[12] ;
 wire \id_stage_i.controller_i.instr_i[13] ;
 wire \id_stage_i.controller_i.instr_i[14] ;
 wire \id_stage_i.controller_i.instr_i[1] ;
 wire \id_stage_i.controller_i.instr_i[25] ;
 wire \id_stage_i.controller_i.instr_i[26] ;
 wire \id_stage_i.controller_i.instr_i[27] ;
 wire \id_stage_i.controller_i.instr_i[28] ;
 wire \id_stage_i.controller_i.instr_i[29] ;
 wire \id_stage_i.controller_i.instr_i[2] ;
 wire \id_stage_i.controller_i.instr_i[30] ;
 wire \id_stage_i.controller_i.instr_i[31] ;
 wire \id_stage_i.controller_i.instr_i[3] ;
 wire \id_stage_i.controller_i.instr_i[4] ;
 wire \id_stage_i.controller_i.instr_i[5] ;
 wire \id_stage_i.controller_i.instr_i[6] ;
 wire \id_stage_i.controller_i.instr_is_compressed_i ;
 wire \id_stage_i.controller_i.instr_valid_i ;
 wire \id_stage_i.controller_i.load_err_d ;
 wire \id_stage_i.controller_i.load_err_q ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[0] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[10] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[11] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[12] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[13] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[14] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[15] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[16] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[17] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[18] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[19] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[1] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[20] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[21] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[22] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[23] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[24] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[25] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[26] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[27] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[28] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[29] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[2] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[30] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[31] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[3] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[4] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[5] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[6] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[7] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[8] ;
 wire \id_stage_i.controller_i.lsu_addr_last_i[9] ;
 wire \id_stage_i.controller_i.store_err_d ;
 wire \id_stage_i.controller_i.store_err_q ;
 wire \id_stage_i.decoder_i.illegal_c_insn_i ;
 wire \id_stage_i.id_fsm_q ;
 wire \if_stage_i.compressed_decoder_i.illegal_instr_o ;
 wire \if_stage_i.compressed_decoder_i.instr_i[0] ;
 wire net593;
 wire net592;
 wire net584;
 wire net600;
 wire net596;
 wire net594;
 wire net624;
 wire net589;
 wire net588;
 wire \if_stage_i.compressed_decoder_i.instr_i[4] ;
 wire net591;
 wire \if_stage_i.compressed_decoder_i.instr_i[6] ;
 wire net587;
 wire net586;
 wire \if_stage_i.compressed_decoder_i.instr_i[9] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[0] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[10] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[11] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[12] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[13] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[14] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[15] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[16] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[17] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[18] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[19] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[1] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[20] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[21] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[22] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[23] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[24] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[25] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[26] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[27] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[28] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[29] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[2] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[30] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[31] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[3] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[4] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[5] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[6] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[7] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[8] ;
 wire \if_stage_i.compressed_decoder_i.instr_o[9] ;
 wire \if_stage_i.compressed_decoder_i.is_compressed_o ;
 wire \if_stage_i.fetch_err ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[10] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[11] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[12] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[13] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[14] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[15] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[16] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[17] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[18] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[19] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[20] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[21] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[22] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[23] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[24] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[25] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[26] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[27] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[28] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[29] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[30] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[31] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[4] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[5] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[6] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[7] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[8] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[9] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_d[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_d[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[10] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[11] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[12] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[13] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[14] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[15] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[16] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[17] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[18] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[19] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[20] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[21] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[22] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[23] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[24] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[25] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[26] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[27] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[28] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[29] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[30] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[31] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[4] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[5] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[6] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[7] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[8] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[9] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[10] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[11] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[12] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[13] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[14] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[15] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[16] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[17] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[18] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[19] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[20] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[21] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[22] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[23] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[24] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[25] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[26] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[27] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[28] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[29] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[30] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[31] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[32] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[33] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[34] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[35] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[36] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[37] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[38] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[39] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[40] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[41] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[42] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[43] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[44] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[45] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[46] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[47] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[48] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[49] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[4] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[50] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[51] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[52] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[53] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[54] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[55] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[56] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[57] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[58] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[59] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[5] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[60] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[61] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[62] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[63] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[6] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[7] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[8] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[9] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ;
 wire \if_stage_i.instr_valid_id_d ;
 wire \load_store_unit_i.data_sign_ext_q ;
 wire \load_store_unit_i.data_type_q[1] ;
 wire \load_store_unit_i.data_type_q[2] ;
 wire \load_store_unit_i.data_we_q ;
 wire \load_store_unit_i.handle_misaligned_q ;
 wire \load_store_unit_i.ls_fsm_cs[0] ;
 wire \load_store_unit_i.ls_fsm_cs[1] ;
 wire \load_store_unit_i.ls_fsm_cs[2] ;
 wire \load_store_unit_i.lsu_err_q ;
 wire \load_store_unit_i.rdata_offset_q[0] ;
 wire \load_store_unit_i.rdata_offset_q[1] ;
 wire \load_store_unit_i.rdata_q[10] ;
 wire \load_store_unit_i.rdata_q[11] ;
 wire \load_store_unit_i.rdata_q[12] ;
 wire \load_store_unit_i.rdata_q[13] ;
 wire \load_store_unit_i.rdata_q[14] ;
 wire \load_store_unit_i.rdata_q[15] ;
 wire \load_store_unit_i.rdata_q[16] ;
 wire \load_store_unit_i.rdata_q[17] ;
 wire \load_store_unit_i.rdata_q[18] ;
 wire \load_store_unit_i.rdata_q[19] ;
 wire \load_store_unit_i.rdata_q[20] ;
 wire \load_store_unit_i.rdata_q[21] ;
 wire \load_store_unit_i.rdata_q[22] ;
 wire \load_store_unit_i.rdata_q[23] ;
 wire \load_store_unit_i.rdata_q[24] ;
 wire \load_store_unit_i.rdata_q[25] ;
 wire \load_store_unit_i.rdata_q[26] ;
 wire \load_store_unit_i.rdata_q[27] ;
 wire \load_store_unit_i.rdata_q[28] ;
 wire \load_store_unit_i.rdata_q[29] ;
 wire \load_store_unit_i.rdata_q[30] ;
 wire \load_store_unit_i.rdata_q[31] ;
 wire \load_store_unit_i.rdata_q[8] ;
 wire \load_store_unit_i.rdata_q[9] ;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1270;
 wire net1271;
 wire net1273;
 wire net1274;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1300;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1243;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1272;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1335;
 wire net1336;
 wire net1413;
 wire net1414;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1510;
 wire net1511;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1529;
 wire net1530;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1547;
 wire net1548;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1564;
 wire net1565;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1575;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;

 sky130_fd_sc_hd__nand2_1 _13505_ (.A(_06633_),
    .B(_06634_),
    .Y(_01505_));
 sky130_fd_sc_hd__inv_1 _13506_ (.A(_11156_),
    .Y(_06635_));
 sky130_fd_sc_hd__nor3_1 _13507_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .B(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .C(_11158_),
    .Y(_06636_));
 sky130_fd_sc_hd__a21oi_1 _13508_ (.A1(_06635_),
    .A2(_06636_),
    .B1(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .Y(_06637_));
 sky130_fd_sc_hd__o21ai_0 _13509_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .A2(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .B1(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .Y(_06638_));
 sky130_fd_sc_hd__nor4b_1 _13510_ (.A(_10946_),
    .B(_11162_),
    .C(_11201_),
    .D_N(_06638_),
    .Y(_06639_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1295 ();
 sky130_fd_sc_hd__nand2_1 _13513_ (.A(_08107_),
    .B(_11155_),
    .Y(_06642_));
 sky130_fd_sc_hd__a21oi_1 _13514_ (.A1(_11158_),
    .A2(_11200_),
    .B1(_06642_),
    .Y(_06643_));
 sky130_fd_sc_hd__o21ai_0 _13515_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .A2(_11158_),
    .B1(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .Y(_06644_));
 sky130_fd_sc_hd__and3_1 _13516_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .B(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .C(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .X(_06645_));
 sky130_fd_sc_hd__a21oi_1 _13517_ (.A1(_08104_),
    .A2(_06644_),
    .B1(_06645_),
    .Y(_06646_));
 sky130_fd_sc_hd__nand2_1 _13518_ (.A(_11007_),
    .B(_11030_),
    .Y(_06647_));
 sky130_fd_sc_hd__or4b_1 _13519_ (.A(_08104_),
    .B(_06647_),
    .C(\cs_registers_i.debug_mode_i ),
    .D_N(_11162_),
    .X(_06648_));
 sky130_fd_sc_hd__o21ai_1 _13520_ (.A1(_12466_),
    .A2(_11002_),
    .B1(_11158_),
    .Y(_06649_));
 sky130_fd_sc_hd__and2_0 _13521_ (.A(_10946_),
    .B(_06649_),
    .X(_06650_));
 sky130_fd_sc_hd__o21ai_1 _13522_ (.A1(_11143_),
    .A2(_10996_),
    .B1(_06650_),
    .Y(_06651_));
 sky130_fd_sc_hd__o2111ai_1 _13523_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .A2(_06646_),
    .B1(_06648_),
    .C1(_06651_),
    .D1(_11009_),
    .Y(_06652_));
 sky130_fd_sc_hd__o32a_1 _13524_ (.A1(_11008_),
    .A2(_06637_),
    .A3(_06639_),
    .B1(_06643_),
    .B2(_06652_),
    .X(_01506_));
 sky130_fd_sc_hd__or2_0 _13525_ (.A(\cs_registers_i.debug_mode_i ),
    .B(_11157_),
    .X(_06653_));
 sky130_fd_sc_hd__nand4_1 _13526_ (.A(_08107_),
    .B(_11156_),
    .C(_06653_),
    .D(_11200_),
    .Y(_06654_));
 sky130_fd_sc_hd__o21ai_0 _13527_ (.A1(_11154_),
    .A2(_06635_),
    .B1(_11143_),
    .Y(_06655_));
 sky130_fd_sc_hd__nor2b_1 _13528_ (.A(_10996_),
    .B_N(_06650_),
    .Y(_06656_));
 sky130_fd_sc_hd__nor2_1 _13529_ (.A(_11037_),
    .B(_11155_),
    .Y(_06657_));
 sky130_fd_sc_hd__a31oi_1 _13530_ (.A1(_11036_),
    .A2(_11156_),
    .A3(_06653_),
    .B1(_11162_),
    .Y(_06658_));
 sky130_fd_sc_hd__o21ai_0 _13531_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .A2(_06658_),
    .B1(_06648_),
    .Y(_06659_));
 sky130_fd_sc_hd__a211oi_1 _13532_ (.A1(_06655_),
    .A2(_06656_),
    .B1(_06657_),
    .C1(_06659_),
    .Y(_06660_));
 sky130_fd_sc_hd__nand2_1 _13533_ (.A(_06654_),
    .B(_06660_),
    .Y(_01507_));
 sky130_fd_sc_hd__a31oi_1 _13534_ (.A1(_11155_),
    .A2(_11158_),
    .A3(_11200_),
    .B1(_11037_),
    .Y(_06661_));
 sky130_fd_sc_hd__nor3_1 _13535_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .B(_08106_),
    .C(_11158_),
    .Y(_06662_));
 sky130_fd_sc_hd__a21oi_1 _13536_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .A2(_11161_),
    .B1(_06662_),
    .Y(_06663_));
 sky130_fd_sc_hd__o21ai_0 _13537_ (.A1(_10944_),
    .A2(_11008_),
    .B1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .Y(_06664_));
 sky130_fd_sc_hd__o21ai_0 _13538_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .A2(_06663_),
    .B1(_06664_),
    .Y(_06665_));
 sky130_fd_sc_hd__nor2_1 _13539_ (.A(_11003_),
    .B(_06651_),
    .Y(_06666_));
 sky130_fd_sc_hd__o311a_1 _13540_ (.A1(_06661_),
    .A2(_06665_),
    .A3(_06666_),
    .B1(_06638_),
    .C1(_06648_),
    .X(_01508_));
 sky130_fd_sc_hd__nand2_1 _13541_ (.A(_11155_),
    .B(_11200_),
    .Y(_06667_));
 sky130_fd_sc_hd__nand2b_1 _13542_ (.A_N(_11003_),
    .B(_06649_),
    .Y(_06668_));
 sky130_fd_sc_hd__a22oi_1 _13543_ (.A1(_11036_),
    .A2(_11158_),
    .B1(_06668_),
    .B2(_10946_),
    .Y(_06669_));
 sky130_fd_sc_hd__a21oi_1 _13544_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .A2(_06667_),
    .B1(_06669_),
    .Y(_01509_));
 sky130_fd_sc_hd__nand4_1 _13545_ (.A(_10946_),
    .B(_10935_),
    .C(_10995_),
    .D(_11142_),
    .Y(_06670_));
 sky130_fd_sc_hd__nand2_1 _13546_ (.A(\cs_registers_i.debug_mode_i ),
    .B(_06670_),
    .Y(_06671_));
 sky130_fd_sc_hd__nand2_1 _13547_ (.A(_11010_),
    .B(_06671_),
    .Y(_01510_));
 sky130_fd_sc_hd__nand2_1 _13548_ (.A(_11034_),
    .B(_12711_),
    .Y(_06672_));
 sky130_fd_sc_hd__o21ai_0 _13549_ (.A1(_11032_),
    .A2(_12455_),
    .B1(_06672_),
    .Y(_01511_));
 sky130_fd_sc_hd__nand2_1 _13550_ (.A(_08443_),
    .B(_08440_),
    .Y(_06673_));
 sky130_fd_sc_hd__nor2_1 _13551_ (.A(_06673_),
    .B(_11197_),
    .Y(_06674_));
 sky130_fd_sc_hd__nand3_1 _13552_ (.A(_08214_),
    .B(_11193_),
    .C(_06674_),
    .Y(_06675_));
 sky130_fd_sc_hd__a21oi_1 _13553_ (.A1(_08269_),
    .A2(_06675_),
    .B1(\id_stage_i.id_fsm_q ),
    .Y(_06676_));
 sky130_fd_sc_hd__a2111oi_0 _13554_ (.A1(_10849_),
    .A2(_11195_),
    .B1(_11197_),
    .C1(_08109_),
    .D1(_11194_),
    .Y(_06677_));
 sky130_fd_sc_hd__nor2_1 _13555_ (.A(_06676_),
    .B(_06677_),
    .Y(_01512_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1293 ();
 sky130_fd_sc_hd__nor2_1 _13558_ (.A(_08948_),
    .B(_03369_),
    .Y(_06680_));
 sky130_fd_sc_hd__a21oi_1 _13559_ (.A1(_10968_),
    .A2(_03369_),
    .B1(_06680_),
    .Y(_06681_));
 sky130_fd_sc_hd__nand2_1 _13560_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[0] ),
    .B(_10952_),
    .Y(_06682_));
 sky130_fd_sc_hd__o21ai_0 _13561_ (.A1(_10952_),
    .A2(_06681_),
    .B1(_06682_),
    .Y(_01513_));
 sky130_fd_sc_hd__mux2i_1 _13562_ (.A0(_09413_),
    .A1(net151),
    .S(_03369_),
    .Y(_06683_));
 sky130_fd_sc_hd__nand2_1 _13563_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[10] ),
    .B(_10952_),
    .Y(_06684_));
 sky130_fd_sc_hd__o21ai_0 _13564_ (.A1(_10952_),
    .A2(_06683_),
    .B1(_06684_),
    .Y(_01514_));
 sky130_fd_sc_hd__nand2b_4 _13565_ (.A_N(_03378_),
    .B(_10721_),
    .Y(_06685_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1290 ();
 sky130_fd_sc_hd__nand2_1 _13569_ (.A(net307),
    .B(net301),
    .Y(_06689_));
 sky130_fd_sc_hd__o21ai_0 _13570_ (.A1(net152),
    .A2(_06685_),
    .B1(_06689_),
    .Y(_06690_));
 sky130_fd_sc_hd__nand2_1 _13571_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[11] ),
    .B(_10952_),
    .Y(_06691_));
 sky130_fd_sc_hd__o21ai_0 _13572_ (.A1(_10952_),
    .A2(_06690_),
    .B1(_06691_),
    .Y(_01515_));
 sky130_fd_sc_hd__mux2i_1 _13573_ (.A0(net153),
    .A1(_09524_),
    .S(_06685_),
    .Y(_06692_));
 sky130_fd_sc_hd__nand2_1 _13574_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[12] ),
    .B(_10952_),
    .Y(_06693_));
 sky130_fd_sc_hd__o21ai_0 _13575_ (.A1(_10952_),
    .A2(_06692_),
    .B1(_06693_),
    .Y(_01516_));
 sky130_fd_sc_hd__nand2_1 _13576_ (.A(_09486_),
    .B(net1207),
    .Y(_06694_));
 sky130_fd_sc_hd__o21ai_0 _13577_ (.A1(net154),
    .A2(_06685_),
    .B1(_06694_),
    .Y(_06695_));
 sky130_fd_sc_hd__nand2_1 _13578_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[13] ),
    .B(_10952_),
    .Y(_06696_));
 sky130_fd_sc_hd__o21ai_0 _13579_ (.A1(_10952_),
    .A2(_06695_),
    .B1(_06696_),
    .Y(_01517_));
 sky130_fd_sc_hd__mux2i_1 _13580_ (.A0(net155),
    .A1(_09606_),
    .S(_06685_),
    .Y(_06697_));
 sky130_fd_sc_hd__nand2_1 _13581_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[14] ),
    .B(_10952_),
    .Y(_06698_));
 sky130_fd_sc_hd__o21ai_0 _13582_ (.A1(_10952_),
    .A2(_06697_),
    .B1(_06698_),
    .Y(_01518_));
 sky130_fd_sc_hd__mux2i_1 _13583_ (.A0(net721),
    .A1(net979),
    .S(_06685_),
    .Y(_06699_));
 sky130_fd_sc_hd__nand2_1 _13584_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[15] ),
    .B(_10952_),
    .Y(_06700_));
 sky130_fd_sc_hd__o21ai_0 _13585_ (.A1(_10952_),
    .A2(_06699_),
    .B1(_06700_),
    .Y(_01519_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1288 ();
 sky130_fd_sc_hd__nand2_1 _13588_ (.A(_09856_),
    .B(net1207),
    .Y(_06703_));
 sky130_fd_sc_hd__o21ai_0 _13589_ (.A1(net157),
    .A2(_06685_),
    .B1(_06703_),
    .Y(_06704_));
 sky130_fd_sc_hd__nand2_1 _13590_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[16] ),
    .B(_10952_),
    .Y(_06705_));
 sky130_fd_sc_hd__o21ai_0 _13591_ (.A1(_10952_),
    .A2(_06704_),
    .B1(_06705_),
    .Y(_01520_));
 sky130_fd_sc_hd__nor2_1 _13592_ (.A(_09784_),
    .B(_03369_),
    .Y(_06706_));
 sky130_fd_sc_hd__nor2_1 _13593_ (.A(net158),
    .B(net1207),
    .Y(_06707_));
 sky130_fd_sc_hd__nand2_1 _13594_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[17] ),
    .B(_10952_),
    .Y(_06708_));
 sky130_fd_sc_hd__o31ai_1 _13595_ (.A1(_10952_),
    .A2(_06706_),
    .A3(_06707_),
    .B1(_06708_),
    .Y(_01521_));
 sky130_fd_sc_hd__nand2_1 _13596_ (.A(net305),
    .B(net1207),
    .Y(_06709_));
 sky130_fd_sc_hd__o21ai_0 _13597_ (.A1(net159),
    .A2(_06685_),
    .B1(_06709_),
    .Y(_06710_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1287 ();
 sky130_fd_sc_hd__nand2_1 _13599_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[18] ),
    .B(_10952_),
    .Y(_06712_));
 sky130_fd_sc_hd__o21ai_0 _13600_ (.A1(_10952_),
    .A2(_06710_),
    .B1(_06712_),
    .Y(_01522_));
 sky130_fd_sc_hd__nand2_1 _13601_ (.A(net304),
    .B(net1207),
    .Y(_06713_));
 sky130_fd_sc_hd__o21ai_0 _13602_ (.A1(net160),
    .A2(_06685_),
    .B1(_06713_),
    .Y(_06714_));
 sky130_fd_sc_hd__nand2_1 _13603_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[19] ),
    .B(_10952_),
    .Y(_06715_));
 sky130_fd_sc_hd__o21ai_0 _13604_ (.A1(_10952_),
    .A2(_06714_),
    .B1(_06715_),
    .Y(_01523_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1286 ();
 sky130_fd_sc_hd__nor2_1 _13606_ (.A(net699),
    .B(_03369_),
    .Y(_06717_));
 sky130_fd_sc_hd__a21oi_1 _13607_ (.A1(net287),
    .A2(_03369_),
    .B1(_06717_),
    .Y(_06718_));
 sky130_fd_sc_hd__nand2_1 _13608_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[1] ),
    .B(_10952_),
    .Y(_06719_));
 sky130_fd_sc_hd__o21ai_0 _13609_ (.A1(_10952_),
    .A2(_06718_),
    .B1(_06719_),
    .Y(_01524_));
 sky130_fd_sc_hd__mux2i_1 _13610_ (.A0(net1007),
    .A1(_10040_),
    .S(_06685_),
    .Y(_06720_));
 sky130_fd_sc_hd__nand2_1 _13611_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[20] ),
    .B(_10952_),
    .Y(_06721_));
 sky130_fd_sc_hd__o21ai_0 _13612_ (.A1(_10952_),
    .A2(_06720_),
    .B1(_06721_),
    .Y(_01525_));
 sky130_fd_sc_hd__mux2i_1 _13613_ (.A0(net162),
    .A1(_10110_),
    .S(_06685_),
    .Y(_06722_));
 sky130_fd_sc_hd__nand2_1 _13614_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[21] ),
    .B(_10952_),
    .Y(_06723_));
 sky130_fd_sc_hd__o21ai_0 _13615_ (.A1(_10952_),
    .A2(_06722_),
    .B1(_06723_),
    .Y(_01526_));
 sky130_fd_sc_hd__mux2i_1 _13616_ (.A0(net1547),
    .A1(_10202_),
    .S(_06685_),
    .Y(_06724_));
 sky130_fd_sc_hd__nand2_1 _13617_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[22] ),
    .B(_10952_),
    .Y(_06725_));
 sky130_fd_sc_hd__o21ai_0 _13618_ (.A1(_10952_),
    .A2(_06724_),
    .B1(_06725_),
    .Y(_01527_));
 sky130_fd_sc_hd__mux2i_1 _13619_ (.A0(net1245),
    .A1(_10259_),
    .S(_06685_),
    .Y(_06726_));
 sky130_fd_sc_hd__nand2_1 _13620_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[23] ),
    .B(_10952_),
    .Y(_06727_));
 sky130_fd_sc_hd__o21ai_0 _13621_ (.A1(_10952_),
    .A2(_06726_),
    .B1(_06727_),
    .Y(_01528_));
 sky130_fd_sc_hd__nor2_1 _13622_ (.A(net1212),
    .B(_03369_),
    .Y(_06728_));
 sky130_fd_sc_hd__a21oi_1 _13623_ (.A1(net775),
    .A2(_03369_),
    .B1(_06728_),
    .Y(_06729_));
 sky130_fd_sc_hd__nand2_1 _13624_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[24] ),
    .B(_10952_),
    .Y(_06730_));
 sky130_fd_sc_hd__o21ai_0 _13625_ (.A1(_10952_),
    .A2(_06729_),
    .B1(_06730_),
    .Y(_01529_));
 sky130_fd_sc_hd__nor2_1 _13626_ (.A(_10407_),
    .B(net1207),
    .Y(_06731_));
 sky130_fd_sc_hd__a21oi_1 _13627_ (.A1(_10332_),
    .A2(net1207),
    .B1(_06731_),
    .Y(_06732_));
 sky130_fd_sc_hd__nand2_1 _13628_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[25] ),
    .B(_10952_),
    .Y(_06733_));
 sky130_fd_sc_hd__o21ai_0 _13629_ (.A1(_10952_),
    .A2(_06732_),
    .B1(_06733_),
    .Y(_01530_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1285 ();
 sky130_fd_sc_hd__nor2_1 _13631_ (.A(net1042),
    .B(net301),
    .Y(_06735_));
 sky130_fd_sc_hd__a21oi_1 _13632_ (.A1(_10437_),
    .A2(net301),
    .B1(_06735_),
    .Y(_06736_));
 sky130_fd_sc_hd__nand2_1 _13633_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[26] ),
    .B(_10952_),
    .Y(_06737_));
 sky130_fd_sc_hd__o21ai_0 _13634_ (.A1(_10952_),
    .A2(_06736_),
    .B1(_06737_),
    .Y(_01531_));
 sky130_fd_sc_hd__mux2i_1 _13635_ (.A0(net168),
    .A1(_10522_),
    .S(_06685_),
    .Y(_06738_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1284 ();
 sky130_fd_sc_hd__nand2_1 _13637_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[27] ),
    .B(_10952_),
    .Y(_06740_));
 sky130_fd_sc_hd__o21ai_0 _13638_ (.A1(_10952_),
    .A2(_06738_),
    .B1(_06740_),
    .Y(_01532_));
 sky130_fd_sc_hd__nor2_1 _13639_ (.A(_10620_),
    .B(_03369_),
    .Y(_06741_));
 sky130_fd_sc_hd__a21oi_1 _13640_ (.A1(net169),
    .A2(_03369_),
    .B1(_06741_),
    .Y(_06742_));
 sky130_fd_sc_hd__nand2_1 _13641_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[28] ),
    .B(_10952_),
    .Y(_06743_));
 sky130_fd_sc_hd__o21ai_0 _13642_ (.A1(_10952_),
    .A2(_06742_),
    .B1(_06743_),
    .Y(_01533_));
 sky130_fd_sc_hd__nor2_1 _13643_ (.A(_10665_),
    .B(net1207),
    .Y(_06744_));
 sky130_fd_sc_hd__a21oi_1 _13644_ (.A1(_10590_),
    .A2(net1207),
    .B1(_06744_),
    .Y(_06745_));
 sky130_fd_sc_hd__nand2_1 _13645_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[29] ),
    .B(_10952_),
    .Y(_06746_));
 sky130_fd_sc_hd__o21ai_0 _13646_ (.A1(_10952_),
    .A2(_06745_),
    .B1(_06746_),
    .Y(_01534_));
 sky130_fd_sc_hd__nor2_1 _13647_ (.A(_10974_),
    .B(net301),
    .Y(_06747_));
 sky130_fd_sc_hd__a21oi_1 _13648_ (.A1(_08795_),
    .A2(net301),
    .B1(_06747_),
    .Y(_06748_));
 sky130_fd_sc_hd__nand2_1 _13649_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[2] ),
    .B(_10952_),
    .Y(_06749_));
 sky130_fd_sc_hd__o21ai_0 _13650_ (.A1(_10952_),
    .A2(_06748_),
    .B1(_06749_),
    .Y(_01535_));
 sky130_fd_sc_hd__nor2_1 _13651_ (.A(_10809_),
    .B(net301),
    .Y(_06750_));
 sky130_fd_sc_hd__a21oi_1 _13652_ (.A1(_10792_),
    .A2(net301),
    .B1(_06750_),
    .Y(_06751_));
 sky130_fd_sc_hd__nand2_1 _13653_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[30] ),
    .B(_10952_),
    .Y(_06752_));
 sky130_fd_sc_hd__o21ai_0 _13654_ (.A1(_10952_),
    .A2(_06751_),
    .B1(_06752_),
    .Y(_01536_));
 sky130_fd_sc_hd__o21ai_0 _13655_ (.A1(net481),
    .A2(_03378_),
    .B1(_10721_),
    .Y(_06753_));
 sky130_fd_sc_hd__nand2_1 _13656_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[31] ),
    .B(_10952_),
    .Y(_06754_));
 sky130_fd_sc_hd__o21ai_0 _13657_ (.A1(_10952_),
    .A2(_06753_),
    .B1(_06754_),
    .Y(_01537_));
 sky130_fd_sc_hd__or3_4 _13658_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .C(_08377_),
    .X(_06755_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1283 ();
 sky130_fd_sc_hd__or3_4 _13660_ (.A(net445),
    .B(_08100_),
    .C(_08290_),
    .X(_06757_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1282 ();
 sky130_fd_sc_hd__nor3_1 _13662_ (.A(_06757_),
    .B(_13358_),
    .C(_06685_),
    .Y(_06759_));
 sky130_fd_sc_hd__a21oi_1 _13663_ (.A1(_13358_),
    .A2(_06685_),
    .B1(_06759_),
    .Y(_06760_));
 sky130_fd_sc_hd__a21oi_1 _13664_ (.A1(_06757_),
    .A2(_13358_),
    .B1(_08502_),
    .Y(_06761_));
 sky130_fd_sc_hd__o21ai_0 _13665_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_by_zero_q ),
    .A2(_06760_),
    .B1(_06761_),
    .Y(_06762_));
 sky130_fd_sc_hd__o21ai_0 _13666_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .A2(_06755_),
    .B1(_06762_),
    .Y(_06763_));
 sky130_fd_sc_hd__nand2_1 _13667_ (.A(net442),
    .B(_06763_),
    .Y(_06764_));
 sky130_fd_sc_hd__and3_4 _13668_ (.A(_08269_),
    .B(net313),
    .C(_06764_),
    .X(_06765_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1278 ();
 sky130_fd_sc_hd__nor3_4 _13673_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .C(_08377_),
    .Y(_06770_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1277 ();
 sky130_fd_sc_hd__nand2_2 _13675_ (.A(_06757_),
    .B(_06770_),
    .Y(_06772_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1276 ();
 sky130_fd_sc_hd__nor2_8 _13677_ (.A(net445),
    .B(_03724_),
    .Y(_06774_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1275 ();
 sky130_fd_sc_hd__a21oi_1 _13679_ (.A1(_13350_),
    .A2(_13469_),
    .B1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[0] ),
    .Y(_06776_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1274 ();
 sky130_fd_sc_hd__nand2_1 _13681_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[32] ),
    .B(_13468_),
    .Y(_06778_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1273 ();
 sky130_fd_sc_hd__nand2_1 _13683_ (.A(net288),
    .B(_13488_),
    .Y(_06780_));
 sky130_fd_sc_hd__nand2_1 _13684_ (.A(_06778_),
    .B(_06780_),
    .Y(_06781_));
 sky130_fd_sc_hd__nor2_1 _13685_ (.A(_06774_),
    .B(_06781_),
    .Y(_06782_));
 sky130_fd_sc_hd__a21oi_1 _13686_ (.A1(_06774_),
    .A2(_06776_),
    .B1(_06782_),
    .Y(_06783_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1272 ();
 sky130_fd_sc_hd__xnor2_1 _13688_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .B(_13350_),
    .Y(_06785_));
 sky130_fd_sc_hd__mux4_1 _13689_ (.A0(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[7] ),
    .A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[4] ),
    .A2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[5] ),
    .A3(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[6] ),
    .S0(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .S1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .X(_06786_));
 sky130_fd_sc_hd__mux4_1 _13690_ (.A0(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[3] ),
    .A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[0] ),
    .A2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[1] ),
    .A3(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[2] ),
    .S0(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .S1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .X(_06787_));
 sky130_fd_sc_hd__xnor2_4 _13691_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .B(_13344_),
    .Y(_06788_));
 sky130_fd_sc_hd__mux2i_1 _13692_ (.A0(_06786_),
    .A1(_06787_),
    .S(_06788_),
    .Y(_06789_));
 sky130_fd_sc_hd__mux4_1 _13693_ (.A0(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[11] ),
    .A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[8] ),
    .A2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[9] ),
    .A3(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[10] ),
    .S0(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .S1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .X(_06790_));
 sky130_fd_sc_hd__mux4_1 _13694_ (.A0(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[15] ),
    .A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[12] ),
    .A2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[13] ),
    .A3(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[14] ),
    .S0(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .S1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .X(_06791_));
 sky130_fd_sc_hd__nor2b_1 _13695_ (.A(_06788_),
    .B_N(_06791_),
    .Y(_06792_));
 sky130_fd_sc_hd__a211oi_1 _13696_ (.A1(_06788_),
    .A2(_06790_),
    .B1(_06792_),
    .C1(_13351_),
    .Y(_06793_));
 sky130_fd_sc_hd__a21oi_1 _13697_ (.A1(_13351_),
    .A2(_06789_),
    .B1(_06793_),
    .Y(_06794_));
 sky130_fd_sc_hd__mux4_1 _13698_ (.A0(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[23] ),
    .A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[20] ),
    .A2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[21] ),
    .A3(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[22] ),
    .S0(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .S1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .X(_06795_));
 sky130_fd_sc_hd__mux4_1 _13699_ (.A0(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[19] ),
    .A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[16] ),
    .A2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[17] ),
    .A3(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[18] ),
    .S0(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .S1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .X(_06796_));
 sky130_fd_sc_hd__mux2i_1 _13700_ (.A0(_06795_),
    .A1(_06796_),
    .S(_06788_),
    .Y(_06797_));
 sky130_fd_sc_hd__mux4_1 _13701_ (.A0(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[27] ),
    .A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[24] ),
    .A2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[25] ),
    .A3(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[26] ),
    .S0(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .S1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .X(_06798_));
 sky130_fd_sc_hd__mux4_1 _13702_ (.A0(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ),
    .A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[28] ),
    .A2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[29] ),
    .A3(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[30] ),
    .S0(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .S1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .X(_06799_));
 sky130_fd_sc_hd__nor2b_1 _13703_ (.A(_06788_),
    .B_N(_06799_),
    .Y(_06800_));
 sky130_fd_sc_hd__a211oi_1 _13704_ (.A1(_06788_),
    .A2(_06798_),
    .B1(_06800_),
    .C1(_13351_),
    .Y(_06801_));
 sky130_fd_sc_hd__a211oi_1 _13705_ (.A1(_13351_),
    .A2(_06797_),
    .B1(_06785_),
    .C1(_06801_),
    .Y(_06802_));
 sky130_fd_sc_hd__a21oi_1 _13706_ (.A1(_06785_),
    .A2(_06794_),
    .B1(_06802_),
    .Y(_06803_));
 sky130_fd_sc_hd__a211oi_1 _13707_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .A2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ),
    .B1(_03724_),
    .C1(_06770_),
    .Y(_06804_));
 sky130_fd_sc_hd__o21ai_0 _13708_ (.A1(_10810_),
    .A2(_06803_),
    .B1(_06804_),
    .Y(_06805_));
 sky130_fd_sc_hd__a221o_1 _13709_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net288),
    .B1(_06783_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .C1(_06805_),
    .X(_06806_));
 sky130_fd_sc_hd__o311ai_0 _13710_ (.A1(net496),
    .A2(_03724_),
    .A3(_06772_),
    .B1(_06806_),
    .C1(_01728_),
    .Y(_06807_));
 sky130_fd_sc_hd__nand3_4 _13711_ (.A(_08269_),
    .B(net313),
    .C(_06764_),
    .Y(_06808_));
 sky130_fd_sc_hd__nor2_4 _13712_ (.A(_01698_),
    .B(_06808_),
    .Y(_06809_));
 sky130_fd_sc_hd__nor2_1 _13713_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[32] ),
    .B(_06809_),
    .Y(_06810_));
 sky130_fd_sc_hd__a21oi_1 _13714_ (.A1(_06765_),
    .A2(_06807_),
    .B1(_06810_),
    .Y(_01538_));
 sky130_fd_sc_hd__nor2_1 _13715_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[33] ),
    .B(_06809_),
    .Y(_06811_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1270 ();
 sky130_fd_sc_hd__a221oi_1 _13718_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(_10970_),
    .B1(_06781_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(_06770_),
    .Y(_06814_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1269 ();
 sky130_fd_sc_hd__nor2_1 _13720_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[33] ),
    .B(_13488_),
    .Y(_06816_));
 sky130_fd_sc_hd__a21oi_1 _13721_ (.A1(net276),
    .A2(_13488_),
    .B1(_06816_),
    .Y(_06817_));
 sky130_fd_sc_hd__or3_4 _13722_ (.A(net445),
    .B(_08100_),
    .C(net739),
    .X(_06818_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1268 ();
 sky130_fd_sc_hd__a311o_1 _13724_ (.A1(_10820_),
    .A2(_10823_),
    .A3(_13469_),
    .B1(_06818_),
    .C1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[1] ),
    .X(_06820_));
 sky130_fd_sc_hd__o211ai_1 _13725_ (.A1(_13333_),
    .A2(_06817_),
    .B1(_06820_),
    .C1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06821_));
 sky130_fd_sc_hd__nand2_1 _13726_ (.A(_06814_),
    .B(_06821_),
    .Y(_06822_));
 sky130_fd_sc_hd__o21ai_0 _13727_ (.A1(net560),
    .A2(_06772_),
    .B1(_06822_),
    .Y(_06823_));
 sky130_fd_sc_hd__nand2_1 _13728_ (.A(_13335_),
    .B(_06823_),
    .Y(_06824_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1267 ();
 sky130_fd_sc_hd__a21oi_1 _13730_ (.A1(_05282_),
    .A2(_06824_),
    .B1(_06808_),
    .Y(_06826_));
 sky130_fd_sc_hd__nor2_1 _13731_ (.A(_06811_),
    .B(_06826_),
    .Y(_01539_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1266 ();
 sky130_fd_sc_hd__nor2_8 _13733_ (.A(_13333_),
    .B(_06755_),
    .Y(_06828_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1265 ();
 sky130_fd_sc_hd__a221oi_1 _13735_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net171),
    .B1(_06817_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(_06770_),
    .Y(_06830_));
 sky130_fd_sc_hd__nor2_1 _13736_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[34] ),
    .B(_13488_),
    .Y(_06831_));
 sky130_fd_sc_hd__a21oi_1 _13737_ (.A1(_10974_),
    .A2(_13488_),
    .B1(_06831_),
    .Y(_06832_));
 sky130_fd_sc_hd__nand2b_4 _13738_ (.A_N(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .Y(_06833_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1263 ();
 sky130_fd_sc_hd__nor2_1 _13741_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[2] ),
    .B(_06818_),
    .Y(_06836_));
 sky130_fd_sc_hd__o21ai_1 _13742_ (.A1(_06833_),
    .A2(_01652_),
    .B1(_06836_),
    .Y(_06837_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1262 ();
 sky130_fd_sc_hd__o211ai_1 _13744_ (.A1(_06774_),
    .A2(_06832_),
    .B1(_06837_),
    .C1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06839_));
 sky130_fd_sc_hd__a22oi_1 _13745_ (.A1(net751),
    .A2(_06828_),
    .B1(_06830_),
    .B2(_06839_),
    .Y(_06840_));
 sky130_fd_sc_hd__o21ai_0 _13746_ (.A1(_03724_),
    .A2(_06840_),
    .B1(_05304_),
    .Y(_06841_));
 sky130_fd_sc_hd__nor2_1 _13747_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[34] ),
    .B(_06809_),
    .Y(_06842_));
 sky130_fd_sc_hd__a21oi_1 _13748_ (.A1(_06765_),
    .A2(_06841_),
    .B1(_06842_),
    .Y(_01540_));
 sky130_fd_sc_hd__a221oi_1 _13749_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net174),
    .B1(_06832_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(_06770_),
    .Y(_06843_));
 sky130_fd_sc_hd__nand2_2 _13750_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_06844_));
 sky130_fd_sc_hd__nor2_1 _13751_ (.A(_06844_),
    .B(_01652_),
    .Y(_06845_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1260 ();
 sky130_fd_sc_hd__mux2i_4 _13754_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[35] ),
    .A1(net174),
    .S(_13488_),
    .Y(_06848_));
 sky130_fd_sc_hd__nand2_1 _13755_ (.A(_06818_),
    .B(_06848_),
    .Y(_06849_));
 sky130_fd_sc_hd__o311ai_4 _13756_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[3] ),
    .A2(_06818_),
    .A3(_06845_),
    .B1(_06849_),
    .C1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06850_));
 sky130_fd_sc_hd__a22oi_1 _13757_ (.A1(net839),
    .A2(_06828_),
    .B1(_06843_),
    .B2(_06850_),
    .Y(_06851_));
 sky130_fd_sc_hd__o21ai_0 _13758_ (.A1(_03724_),
    .A2(_06851_),
    .B1(_05346_),
    .Y(_06852_));
 sky130_fd_sc_hd__nor2_1 _13759_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[35] ),
    .B(_06809_),
    .Y(_06853_));
 sky130_fd_sc_hd__a21oi_1 _13760_ (.A1(_06765_),
    .A2(_06852_),
    .B1(_06853_),
    .Y(_01541_));
 sky130_fd_sc_hd__nor2_1 _13761_ (.A(_10810_),
    .B(_06848_),
    .Y(_06854_));
 sky130_fd_sc_hd__a211oi_1 _13762_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net175),
    .B1(_06770_),
    .C1(_06854_),
    .Y(_06855_));
 sky130_fd_sc_hd__nor2_1 _13763_ (.A(_13345_),
    .B(_01657_),
    .Y(_06856_));
 sky130_fd_sc_hd__mux2i_2 _13764_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[36] ),
    .A1(net175),
    .S(_13488_),
    .Y(_06857_));
 sky130_fd_sc_hd__nand2_1 _13765_ (.A(_06818_),
    .B(_06857_),
    .Y(_06858_));
 sky130_fd_sc_hd__o311ai_2 _13766_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[4] ),
    .A2(_06818_),
    .A3(_06856_),
    .B1(_06858_),
    .C1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06859_));
 sky130_fd_sc_hd__a22oi_1 _13767_ (.A1(net1458),
    .A2(_06828_),
    .B1(_06855_),
    .B2(_06859_),
    .Y(_06860_));
 sky130_fd_sc_hd__o21ai_0 _13768_ (.A1(_03724_),
    .A2(_06860_),
    .B1(_02098_),
    .Y(_06861_));
 sky130_fd_sc_hd__nor2_1 _13769_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[36] ),
    .B(_06809_),
    .Y(_06862_));
 sky130_fd_sc_hd__a21oi_1 _13770_ (.A1(_06765_),
    .A2(_06861_),
    .B1(_06862_),
    .Y(_01542_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1259 ();
 sky130_fd_sc_hd__nand2_1 _13772_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[37] ),
    .B(_06808_),
    .Y(_06864_));
 sky130_fd_sc_hd__nor2_1 _13773_ (.A(_13335_),
    .B(_02172_),
    .Y(_06865_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1258 ();
 sky130_fd_sc_hd__nor2_1 _13775_ (.A(_10810_),
    .B(_06857_),
    .Y(_06867_));
 sky130_fd_sc_hd__a211oi_1 _13776_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net1062),
    .B1(_06770_),
    .C1(_06867_),
    .Y(_06868_));
 sky130_fd_sc_hd__nand2b_2 _13777_ (.A_N(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_06869_));
 sky130_fd_sc_hd__nor2_1 _13778_ (.A(_06869_),
    .B(_01657_),
    .Y(_06870_));
 sky130_fd_sc_hd__mux2i_2 _13779_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[37] ),
    .A1(net176),
    .S(_13488_),
    .Y(_06871_));
 sky130_fd_sc_hd__nand2_1 _13780_ (.A(_06818_),
    .B(_06871_),
    .Y(_06872_));
 sky130_fd_sc_hd__o311ai_2 _13781_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[5] ),
    .A2(_06757_),
    .A3(_06870_),
    .B1(_06872_),
    .C1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06873_));
 sky130_fd_sc_hd__a221oi_1 _13782_ (.A1(net797),
    .A2(_06828_),
    .B1(_06868_),
    .B2(_06873_),
    .C1(_03724_),
    .Y(_06874_));
 sky130_fd_sc_hd__o21ai_0 _13783_ (.A1(_06865_),
    .A2(_06874_),
    .B1(_06765_),
    .Y(_06875_));
 sky130_fd_sc_hd__nand2_1 _13784_ (.A(_06864_),
    .B(_06875_),
    .Y(_01543_));
 sky130_fd_sc_hd__nand2_1 _13785_ (.A(_08693_),
    .B(net301),
    .Y(_06876_));
 sky130_fd_sc_hd__o21ai_0 _13786_ (.A1(net174),
    .A2(_06685_),
    .B1(_06876_),
    .Y(_06877_));
 sky130_fd_sc_hd__nand2_1 _13787_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[3] ),
    .B(_10952_),
    .Y(_06878_));
 sky130_fd_sc_hd__o21ai_0 _13788_ (.A1(_10952_),
    .A2(_06877_),
    .B1(_06878_),
    .Y(_01544_));
 sky130_fd_sc_hd__o221a_1 _13789_ (.A1(_08502_),
    .A2(_09159_),
    .B1(_06871_),
    .B2(_10810_),
    .C1(_06755_),
    .X(_06879_));
 sky130_fd_sc_hd__nor2_1 _13790_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[38] ),
    .B(_13488_),
    .Y(_06880_));
 sky130_fd_sc_hd__a21oi_1 _13791_ (.A1(_09159_),
    .A2(_13488_),
    .B1(_06880_),
    .Y(_06881_));
 sky130_fd_sc_hd__nor2_1 _13792_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[6] ),
    .B(_06818_),
    .Y(_06882_));
 sky130_fd_sc_hd__o21ai_1 _13793_ (.A1(_06833_),
    .A2(_01657_),
    .B1(_06882_),
    .Y(_06883_));
 sky130_fd_sc_hd__o211ai_1 _13794_ (.A1(_06774_),
    .A2(_06881_),
    .B1(_06883_),
    .C1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06884_));
 sky130_fd_sc_hd__a22oi_1 _13795_ (.A1(net573),
    .A2(_06828_),
    .B1(_06879_),
    .B2(_06884_),
    .Y(_06885_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1257 ();
 sky130_fd_sc_hd__o22ai_1 _13797_ (.A1(_02284_),
    .A2(_02345_),
    .B1(_06885_),
    .B2(_03724_),
    .Y(_06887_));
 sky130_fd_sc_hd__nor2_1 _13798_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[38] ),
    .B(_06809_),
    .Y(_06888_));
 sky130_fd_sc_hd__a21oi_1 _13799_ (.A1(_06765_),
    .A2(_06887_),
    .B1(_06888_),
    .Y(_01545_));
 sky130_fd_sc_hd__nand2_1 _13800_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[39] ),
    .B(_13468_),
    .Y(_06889_));
 sky130_fd_sc_hd__o21ai_0 _13801_ (.A1(net1023),
    .A2(_13468_),
    .B1(_06889_),
    .Y(_06890_));
 sky130_fd_sc_hd__o21ai_0 _13802_ (.A1(_13333_),
    .A2(_06890_),
    .B1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06891_));
 sky130_fd_sc_hd__nor2_1 _13803_ (.A(_06844_),
    .B(_01657_),
    .Y(_06892_));
 sky130_fd_sc_hd__nor3_1 _13804_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[7] ),
    .B(_06757_),
    .C(_06892_),
    .Y(_06893_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1256 ();
 sky130_fd_sc_hd__a221oi_1 _13806_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net178),
    .B1(_06881_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(_06770_),
    .Y(_06895_));
 sky130_fd_sc_hd__o21ai_0 _13807_ (.A1(_06891_),
    .A2(_06893_),
    .B1(_06895_),
    .Y(_06896_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1255 ();
 sky130_fd_sc_hd__a21oi_1 _13809_ (.A1(net768),
    .A2(_06828_),
    .B1(_03724_),
    .Y(_06898_));
 sky130_fd_sc_hd__nor2_1 _13810_ (.A(_13335_),
    .B(_02453_),
    .Y(_06899_));
 sky130_fd_sc_hd__a21oi_1 _13811_ (.A1(_06896_),
    .A2(_06898_),
    .B1(_06899_),
    .Y(_06900_));
 sky130_fd_sc_hd__nand2_1 _13812_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[39] ),
    .B(_06808_),
    .Y(_06901_));
 sky130_fd_sc_hd__o21ai_0 _13813_ (.A1(_06808_),
    .A2(_06900_),
    .B1(_06901_),
    .Y(_01546_));
 sky130_fd_sc_hd__nand2_1 _13814_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[40] ),
    .B(_13468_),
    .Y(_06902_));
 sky130_fd_sc_hd__o21ai_0 _13815_ (.A1(_09303_),
    .A2(_13468_),
    .B1(_06902_),
    .Y(_06903_));
 sky130_fd_sc_hd__o21ai_0 _13816_ (.A1(_13333_),
    .A2(_06903_),
    .B1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06904_));
 sky130_fd_sc_hd__nor2_1 _13817_ (.A(_13345_),
    .B(_13475_),
    .Y(_06905_));
 sky130_fd_sc_hd__nor3_2 _13818_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[8] ),
    .B(_06757_),
    .C(_06905_),
    .Y(_06906_));
 sky130_fd_sc_hd__a221oi_1 _13819_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net179),
    .B1(_06890_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(_06770_),
    .Y(_06907_));
 sky130_fd_sc_hd__o21ai_1 _13820_ (.A1(_06904_),
    .A2(_06906_),
    .B1(_06907_),
    .Y(_06908_));
 sky130_fd_sc_hd__a21oi_1 _13821_ (.A1(_09184_),
    .A2(_06828_),
    .B1(_03724_),
    .Y(_06909_));
 sky130_fd_sc_hd__nor2_1 _13822_ (.A(_13335_),
    .B(_02540_),
    .Y(_06910_));
 sky130_fd_sc_hd__a21oi_1 _13823_ (.A1(_06908_),
    .A2(_06909_),
    .B1(_06910_),
    .Y(_06911_));
 sky130_fd_sc_hd__nand2_1 _13824_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[40] ),
    .B(_06808_),
    .Y(_06912_));
 sky130_fd_sc_hd__o21ai_0 _13825_ (.A1(_06808_),
    .A2(_06911_),
    .B1(_06912_),
    .Y(_01547_));
 sky130_fd_sc_hd__nand2_1 _13826_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[41] ),
    .B(_13468_),
    .Y(_06913_));
 sky130_fd_sc_hd__nand2_1 _13827_ (.A(net180),
    .B(_13488_),
    .Y(_06914_));
 sky130_fd_sc_hd__nand2_1 _13828_ (.A(_06913_),
    .B(_06914_),
    .Y(_06915_));
 sky130_fd_sc_hd__o21ai_0 _13829_ (.A1(_13333_),
    .A2(_06915_),
    .B1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06916_));
 sky130_fd_sc_hd__nor2_1 _13830_ (.A(_06869_),
    .B(_13475_),
    .Y(_06917_));
 sky130_fd_sc_hd__nor3_1 _13831_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ),
    .B(_06757_),
    .C(_06917_),
    .Y(_06918_));
 sky130_fd_sc_hd__a221oi_1 _13832_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net180),
    .B1(_06903_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(_06770_),
    .Y(_06919_));
 sky130_fd_sc_hd__o21ai_0 _13833_ (.A1(_06916_),
    .A2(_06918_),
    .B1(_06919_),
    .Y(_06920_));
 sky130_fd_sc_hd__a21oi_1 _13834_ (.A1(net1121),
    .A2(_06828_),
    .B1(_03724_),
    .Y(_06921_));
 sky130_fd_sc_hd__a21oi_1 _13835_ (.A1(_06920_),
    .A2(_06921_),
    .B1(_02643_),
    .Y(_06922_));
 sky130_fd_sc_hd__nand2_1 _13836_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[41] ),
    .B(_06808_),
    .Y(_06923_));
 sky130_fd_sc_hd__o21ai_0 _13837_ (.A1(_06808_),
    .A2(_06922_),
    .B1(_06923_),
    .Y(_01548_));
 sky130_fd_sc_hd__nand2_1 _13838_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[42] ),
    .B(_13468_),
    .Y(_06924_));
 sky130_fd_sc_hd__nand2_1 _13839_ (.A(net151),
    .B(_13488_),
    .Y(_06925_));
 sky130_fd_sc_hd__nand2_1 _13840_ (.A(_06924_),
    .B(_06925_),
    .Y(_06926_));
 sky130_fd_sc_hd__o21ai_0 _13841_ (.A1(_13333_),
    .A2(_06926_),
    .B1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06927_));
 sky130_fd_sc_hd__nor2_1 _13842_ (.A(_06833_),
    .B(_13475_),
    .Y(_06928_));
 sky130_fd_sc_hd__nor3_1 _13843_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[10] ),
    .B(_06757_),
    .C(_06928_),
    .Y(_06929_));
 sky130_fd_sc_hd__a221oi_1 _13844_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net151),
    .B1(_06915_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(_06770_),
    .Y(_06930_));
 sky130_fd_sc_hd__o21ai_0 _13845_ (.A1(_06927_),
    .A2(_06929_),
    .B1(_06930_),
    .Y(_06931_));
 sky130_fd_sc_hd__a21oi_1 _13846_ (.A1(_09380_),
    .A2(_06828_),
    .B1(_03724_),
    .Y(_06932_));
 sky130_fd_sc_hd__a22oi_1 _13847_ (.A1(_03724_),
    .A2(_02753_),
    .B1(_06931_),
    .B2(_06932_),
    .Y(_06933_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1254 ();
 sky130_fd_sc_hd__nand2_1 _13849_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[42] ),
    .B(_06808_),
    .Y(_06935_));
 sky130_fd_sc_hd__o21ai_0 _13850_ (.A1(_06808_),
    .A2(_06933_),
    .B1(_06935_),
    .Y(_01549_));
 sky130_fd_sc_hd__nor2_1 _13851_ (.A(_13335_),
    .B(_02829_),
    .Y(_06936_));
 sky130_fd_sc_hd__a221oi_1 _13852_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net152),
    .B1(_06926_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(_06770_),
    .Y(_06937_));
 sky130_fd_sc_hd__nor2_1 _13853_ (.A(_13475_),
    .B(_06844_),
    .Y(_06938_));
 sky130_fd_sc_hd__mux2i_2 _13854_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[43] ),
    .A1(net152),
    .S(_13488_),
    .Y(_06939_));
 sky130_fd_sc_hd__nand2_1 _13855_ (.A(_06818_),
    .B(_06939_),
    .Y(_06940_));
 sky130_fd_sc_hd__o311ai_2 _13856_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[11] ),
    .A2(_06757_),
    .A3(_06938_),
    .B1(_06940_),
    .C1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06941_));
 sky130_fd_sc_hd__o21ai_0 _13857_ (.A1(net1188),
    .A2(_06772_),
    .B1(_13335_),
    .Y(_06942_));
 sky130_fd_sc_hd__a21oi_1 _13858_ (.A1(_06937_),
    .A2(_06941_),
    .B1(_06942_),
    .Y(_06943_));
 sky130_fd_sc_hd__nor2_1 _13859_ (.A(_06936_),
    .B(_06943_),
    .Y(_06944_));
 sky130_fd_sc_hd__nand2_1 _13860_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[43] ),
    .B(_06808_),
    .Y(_06945_));
 sky130_fd_sc_hd__o21ai_0 _13861_ (.A1(_06808_),
    .A2(_06944_),
    .B1(_06945_),
    .Y(_01550_));
 sky130_fd_sc_hd__nand2_1 _13862_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[44] ),
    .B(_06808_),
    .Y(_06946_));
 sky130_fd_sc_hd__nor2_1 _13863_ (.A(_13335_),
    .B(_02969_),
    .Y(_06947_));
 sky130_fd_sc_hd__nor2_1 _13864_ (.A(_10810_),
    .B(_06939_),
    .Y(_06948_));
 sky130_fd_sc_hd__a211oi_1 _13865_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net153),
    .B1(_06770_),
    .C1(_06948_),
    .Y(_06949_));
 sky130_fd_sc_hd__nor2_1 _13866_ (.A(_13345_),
    .B(_13481_),
    .Y(_06950_));
 sky130_fd_sc_hd__mux2i_1 _13867_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[44] ),
    .A1(net153),
    .S(_13488_),
    .Y(_06951_));
 sky130_fd_sc_hd__nand2_1 _13868_ (.A(_06818_),
    .B(_06951_),
    .Y(_06952_));
 sky130_fd_sc_hd__o311ai_1 _13869_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[12] ),
    .A2(_06757_),
    .A3(_06950_),
    .B1(_06952_),
    .C1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06953_));
 sky130_fd_sc_hd__a221oi_1 _13870_ (.A1(_09553_),
    .A2(_06828_),
    .B1(_06949_),
    .B2(_06953_),
    .C1(_03724_),
    .Y(_06954_));
 sky130_fd_sc_hd__o21ai_0 _13871_ (.A1(_06947_),
    .A2(_06954_),
    .B1(_06765_),
    .Y(_06955_));
 sky130_fd_sc_hd__nand2_1 _13872_ (.A(_06946_),
    .B(_06955_),
    .Y(_01551_));
 sky130_fd_sc_hd__nor2_1 _13873_ (.A(_10810_),
    .B(_06951_),
    .Y(_06956_));
 sky130_fd_sc_hd__a211oi_1 _13874_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net154),
    .B1(_06770_),
    .C1(_06956_),
    .Y(_06957_));
 sky130_fd_sc_hd__nor2_1 _13875_ (.A(_06869_),
    .B(_13481_),
    .Y(_06958_));
 sky130_fd_sc_hd__mux2i_1 _13876_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[45] ),
    .A1(net154),
    .S(_13488_),
    .Y(_06959_));
 sky130_fd_sc_hd__nand2_1 _13877_ (.A(_06818_),
    .B(_06959_),
    .Y(_06960_));
 sky130_fd_sc_hd__o311ai_1 _13878_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[13] ),
    .A2(_06757_),
    .A3(_06958_),
    .B1(_06960_),
    .C1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06961_));
 sky130_fd_sc_hd__a221oi_1 _13879_ (.A1(net648),
    .A2(_06828_),
    .B1(_06957_),
    .B2(_06961_),
    .C1(_03724_),
    .Y(_06962_));
 sky130_fd_sc_hd__a21oi_1 _13880_ (.A1(_03724_),
    .A2(_03075_),
    .B1(_06962_),
    .Y(_06963_));
 sky130_fd_sc_hd__nand2_1 _13881_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[45] ),
    .B(_06808_),
    .Y(_06964_));
 sky130_fd_sc_hd__o21ai_0 _13882_ (.A1(_06808_),
    .A2(_06963_),
    .B1(_06964_),
    .Y(_01552_));
 sky130_fd_sc_hd__a21oi_1 _13883_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net1583),
    .B1(_06770_),
    .Y(_06965_));
 sky130_fd_sc_hd__nor2_1 _13884_ (.A(_06833_),
    .B(_13481_),
    .Y(_06966_));
 sky130_fd_sc_hd__mux2i_1 _13885_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[46] ),
    .A1(net1583),
    .S(_13488_),
    .Y(_06967_));
 sky130_fd_sc_hd__nand2_1 _13886_ (.A(_06818_),
    .B(_06967_),
    .Y(_06968_));
 sky130_fd_sc_hd__o311ai_1 _13887_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[14] ),
    .A2(_06757_),
    .A3(_06966_),
    .B1(_06968_),
    .C1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06969_));
 sky130_fd_sc_hd__o211ai_1 _13888_ (.A1(_10810_),
    .A2(_06959_),
    .B1(_06965_),
    .C1(_06969_),
    .Y(_06970_));
 sky130_fd_sc_hd__a21oi_1 _13889_ (.A1(_09632_),
    .A2(_06828_),
    .B1(_03724_),
    .Y(_06971_));
 sky130_fd_sc_hd__a21oi_1 _13890_ (.A1(_06970_),
    .A2(_06971_),
    .B1(_03194_),
    .Y(_06972_));
 sky130_fd_sc_hd__nand2_1 _13891_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[46] ),
    .B(_06808_),
    .Y(_06973_));
 sky130_fd_sc_hd__o21ai_0 _13892_ (.A1(_06808_),
    .A2(_06972_),
    .B1(_06973_),
    .Y(_01553_));
 sky130_fd_sc_hd__mux2i_2 _13893_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[47] ),
    .A1(net721),
    .S(_13488_),
    .Y(_06974_));
 sky130_fd_sc_hd__nor2_1 _13894_ (.A(_06844_),
    .B(_13481_),
    .Y(_06975_));
 sky130_fd_sc_hd__nor3_1 _13895_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[15] ),
    .B(_06818_),
    .C(_06975_),
    .Y(_06976_));
 sky130_fd_sc_hd__a21oi_1 _13896_ (.A1(_06757_),
    .A2(_06974_),
    .B1(_06976_),
    .Y(_06977_));
 sky130_fd_sc_hd__a21oi_1 _13897_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net719),
    .B1(_06770_),
    .Y(_06978_));
 sky130_fd_sc_hd__o21ai_0 _13898_ (.A1(_10810_),
    .A2(_06967_),
    .B1(_06978_),
    .Y(_06979_));
 sky130_fd_sc_hd__a21oi_1 _13899_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .A2(_06977_),
    .B1(_06979_),
    .Y(_06980_));
 sky130_fd_sc_hd__o21ai_0 _13900_ (.A1(net837),
    .A2(_06772_),
    .B1(_13335_),
    .Y(_06981_));
 sky130_fd_sc_hd__o22ai_1 _13901_ (.A1(_13335_),
    .A2(_03343_),
    .B1(_06980_),
    .B2(_06981_),
    .Y(_06982_));
 sky130_fd_sc_hd__nand2_1 _13902_ (.A(_06809_),
    .B(_06982_),
    .Y(_06983_));
 sky130_fd_sc_hd__o21ai_0 _13903_ (.A1(_09680_),
    .A2(_06809_),
    .B1(_06983_),
    .Y(_01554_));
 sky130_fd_sc_hd__nand2_1 _13904_ (.A(net308),
    .B(net301),
    .Y(_06984_));
 sky130_fd_sc_hd__o21ai_0 _13905_ (.A1(net175),
    .A2(_06685_),
    .B1(_06984_),
    .Y(_06985_));
 sky130_fd_sc_hd__nand2_1 _13906_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[4] ),
    .B(_10952_),
    .Y(_06986_));
 sky130_fd_sc_hd__o21ai_0 _13907_ (.A1(_10952_),
    .A2(_06985_),
    .B1(_06986_),
    .Y(_01555_));
 sky130_fd_sc_hd__nor2_1 _13908_ (.A(_10810_),
    .B(_06974_),
    .Y(_06987_));
 sky130_fd_sc_hd__a211oi_1 _13909_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net157),
    .B1(_06770_),
    .C1(_06987_),
    .Y(_06988_));
 sky130_fd_sc_hd__a21oi_1 _13910_ (.A1(_13350_),
    .A2(_13490_),
    .B1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[16] ),
    .Y(_06989_));
 sky130_fd_sc_hd__nor2_1 _13911_ (.A(_06818_),
    .B(_06989_),
    .Y(_06990_));
 sky130_fd_sc_hd__mux2i_1 _13912_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[48] ),
    .A1(net157),
    .S(_13488_),
    .Y(_06991_));
 sky130_fd_sc_hd__nor2_1 _13913_ (.A(_06774_),
    .B(_06991_),
    .Y(_06992_));
 sky130_fd_sc_hd__o21ai_0 _13914_ (.A1(_06990_),
    .A2(_06992_),
    .B1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_06993_));
 sky130_fd_sc_hd__a221oi_2 _13915_ (.A1(_09821_),
    .A2(_06828_),
    .B1(_06988_),
    .B2(_06993_),
    .C1(_03724_),
    .Y(_06994_));
 sky130_fd_sc_hd__a21oi_1 _13916_ (.A1(_03724_),
    .A2(_03462_),
    .B1(_06994_),
    .Y(_06995_));
 sky130_fd_sc_hd__nand2_1 _13917_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[48] ),
    .B(_06808_),
    .Y(_06996_));
 sky130_fd_sc_hd__o21ai_0 _13918_ (.A1(_06808_),
    .A2(_06995_),
    .B1(_06996_),
    .Y(_01556_));
 sky130_fd_sc_hd__mux2i_1 _13919_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[49] ),
    .A1(net158),
    .S(_13488_),
    .Y(_06997_));
 sky130_fd_sc_hd__nor2b_1 _13920_ (.A(_10824_),
    .B_N(_13490_),
    .Y(_06998_));
 sky130_fd_sc_hd__o21ai_2 _13921_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[17] ),
    .A2(_06998_),
    .B1(_06774_),
    .Y(_06999_));
 sky130_fd_sc_hd__o21ai_0 _13922_ (.A1(_06774_),
    .A2(_06997_),
    .B1(_06999_),
    .Y(_07000_));
 sky130_fd_sc_hd__a21oi_1 _13923_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net158),
    .B1(_06770_),
    .Y(_07001_));
 sky130_fd_sc_hd__o21ai_0 _13924_ (.A1(_10810_),
    .A2(_06991_),
    .B1(_07001_),
    .Y(_07002_));
 sky130_fd_sc_hd__a21oi_1 _13925_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .A2(_07000_),
    .B1(_07002_),
    .Y(_07003_));
 sky130_fd_sc_hd__o21ai_0 _13926_ (.A1(net777),
    .A2(_06772_),
    .B1(_13335_),
    .Y(_07004_));
 sky130_fd_sc_hd__nor2_1 _13927_ (.A(_07003_),
    .B(_07004_),
    .Y(_07005_));
 sky130_fd_sc_hd__a21oi_1 _13928_ (.A1(_03724_),
    .A2(_03598_),
    .B1(_07005_),
    .Y(_07006_));
 sky130_fd_sc_hd__nand2_1 _13929_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[49] ),
    .B(_06808_),
    .Y(_07007_));
 sky130_fd_sc_hd__o21ai_0 _13930_ (.A1(_06808_),
    .A2(_07006_),
    .B1(_07007_),
    .Y(_01557_));
 sky130_fd_sc_hd__nand2_1 _13931_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[50] ),
    .B(_06808_),
    .Y(_07008_));
 sky130_fd_sc_hd__mux2i_1 _13932_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[50] ),
    .A1(net1241),
    .S(_13488_),
    .Y(_07009_));
 sky130_fd_sc_hd__nor2_1 _13933_ (.A(_06833_),
    .B(_13493_),
    .Y(_07010_));
 sky130_fd_sc_hd__nor3_1 _13934_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[18] ),
    .B(_06818_),
    .C(_07010_),
    .Y(_07011_));
 sky130_fd_sc_hd__a21oi_1 _13935_ (.A1(_06757_),
    .A2(_07009_),
    .B1(_07011_),
    .Y(_07012_));
 sky130_fd_sc_hd__a21oi_1 _13936_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net1241),
    .B1(_06770_),
    .Y(_07013_));
 sky130_fd_sc_hd__o21ai_0 _13937_ (.A1(_10810_),
    .A2(_06997_),
    .B1(_07013_),
    .Y(_07014_));
 sky130_fd_sc_hd__a21oi_1 _13938_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .A2(_07012_),
    .B1(_07014_),
    .Y(_07015_));
 sky130_fd_sc_hd__o21ai_0 _13939_ (.A1(net960),
    .A2(_06772_),
    .B1(_13335_),
    .Y(_07016_));
 sky130_fd_sc_hd__o21ai_0 _13940_ (.A1(_07015_),
    .A2(_07016_),
    .B1(_03725_),
    .Y(_07017_));
 sky130_fd_sc_hd__nand2_1 _13941_ (.A(_06765_),
    .B(_07017_),
    .Y(_07018_));
 sky130_fd_sc_hd__nand2_1 _13942_ (.A(_07008_),
    .B(_07018_),
    .Y(_01558_));
 sky130_fd_sc_hd__nand2_1 _13943_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[51] ),
    .B(_06808_),
    .Y(_07019_));
 sky130_fd_sc_hd__nor2_1 _13944_ (.A(_10810_),
    .B(_07009_),
    .Y(_07020_));
 sky130_fd_sc_hd__a211oi_1 _13945_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net1261),
    .B1(_06770_),
    .C1(_07020_),
    .Y(_07021_));
 sky130_fd_sc_hd__nor2_1 _13946_ (.A(_06844_),
    .B(_13493_),
    .Y(_07022_));
 sky130_fd_sc_hd__mux2i_2 _13947_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[51] ),
    .A1(net1261),
    .S(_13488_),
    .Y(_07023_));
 sky130_fd_sc_hd__nand2_1 _13948_ (.A(_06818_),
    .B(_07023_),
    .Y(_07024_));
 sky130_fd_sc_hd__o311ai_2 _13949_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[19] ),
    .A2(_06757_),
    .A3(_07022_),
    .B1(_07024_),
    .C1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_07025_));
 sky130_fd_sc_hd__a221oi_1 _13950_ (.A1(_09969_),
    .A2(_06828_),
    .B1(_07021_),
    .B2(_07025_),
    .C1(_03724_),
    .Y(_07026_));
 sky130_fd_sc_hd__nor2_1 _13951_ (.A(_13335_),
    .B(_03853_),
    .Y(_07027_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1253 ();
 sky130_fd_sc_hd__o21ai_0 _13953_ (.A1(_07026_),
    .A2(_07027_),
    .B1(_06765_),
    .Y(_07029_));
 sky130_fd_sc_hd__nand2_1 _13954_ (.A(_07019_),
    .B(_07029_),
    .Y(_01559_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1252 ();
 sky130_fd_sc_hd__nor2_1 _13956_ (.A(_10810_),
    .B(_07023_),
    .Y(_07031_));
 sky130_fd_sc_hd__a211oi_1 _13957_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net693),
    .B1(_06770_),
    .C1(_07031_),
    .Y(_07032_));
 sky130_fd_sc_hd__nor2_1 _13958_ (.A(_13345_),
    .B(_13497_),
    .Y(_07033_));
 sky130_fd_sc_hd__mux2i_1 _13959_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[52] ),
    .A1(net692),
    .S(_13488_),
    .Y(_07034_));
 sky130_fd_sc_hd__nand2_1 _13960_ (.A(_06818_),
    .B(_07034_),
    .Y(_07035_));
 sky130_fd_sc_hd__o311ai_1 _13961_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[20] ),
    .A2(_06757_),
    .A3(_07033_),
    .B1(_07035_),
    .C1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_07036_));
 sky130_fd_sc_hd__a221oi_1 _13962_ (.A1(_10061_),
    .A2(_06828_),
    .B1(_07032_),
    .B2(_07036_),
    .C1(_03724_),
    .Y(_07037_));
 sky130_fd_sc_hd__a21oi_1 _13963_ (.A1(_03724_),
    .A2(_03968_),
    .B1(_07037_),
    .Y(_07038_));
 sky130_fd_sc_hd__nand2_1 _13964_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[52] ),
    .B(_06808_),
    .Y(_07039_));
 sky130_fd_sc_hd__o21ai_0 _13965_ (.A1(_06808_),
    .A2(_07038_),
    .B1(_07039_),
    .Y(_01560_));
 sky130_fd_sc_hd__nand2_1 _13966_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[53] ),
    .B(_06808_),
    .Y(_07040_));
 sky130_fd_sc_hd__nand3_1 _13967_ (.A(_03724_),
    .B(_04105_),
    .C(_06765_),
    .Y(_07041_));
 sky130_fd_sc_hd__nor2_1 _13968_ (.A(_06869_),
    .B(_13497_),
    .Y(_07042_));
 sky130_fd_sc_hd__mux2i_1 _13969_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[53] ),
    .A1(net1255),
    .S(_13488_),
    .Y(_07043_));
 sky130_fd_sc_hd__nand2_1 _13970_ (.A(_06818_),
    .B(_07043_),
    .Y(_07044_));
 sky130_fd_sc_hd__o311ai_0 _13971_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[21] ),
    .A2(_06818_),
    .A3(_07042_),
    .B1(_07044_),
    .C1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_07045_));
 sky130_fd_sc_hd__a21oi_1 _13972_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net1256),
    .B1(_06770_),
    .Y(_07046_));
 sky130_fd_sc_hd__o211ai_1 _13973_ (.A1(_10810_),
    .A2(_07034_),
    .B1(_07045_),
    .C1(_07046_),
    .Y(_07047_));
 sky130_fd_sc_hd__nand2_1 _13974_ (.A(_10130_),
    .B(_06828_),
    .Y(_07048_));
 sky130_fd_sc_hd__nand4_1 _13975_ (.A(_13335_),
    .B(_06765_),
    .C(_07047_),
    .D(_07048_),
    .Y(_07049_));
 sky130_fd_sc_hd__nand3_1 _13976_ (.A(_07040_),
    .B(_07041_),
    .C(_07049_),
    .Y(_01561_));
 sky130_fd_sc_hd__nor2_1 _13977_ (.A(_10810_),
    .B(_07043_),
    .Y(_07050_));
 sky130_fd_sc_hd__a211oi_1 _13978_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net992),
    .B1(_06770_),
    .C1(_07050_),
    .Y(_07051_));
 sky130_fd_sc_hd__nor2_1 _13979_ (.A(_06833_),
    .B(_13497_),
    .Y(_07052_));
 sky130_fd_sc_hd__mux2i_1 _13980_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[54] ),
    .A1(net992),
    .S(_13488_),
    .Y(_07053_));
 sky130_fd_sc_hd__nand2_1 _13981_ (.A(_06818_),
    .B(_07053_),
    .Y(_07054_));
 sky130_fd_sc_hd__o311ai_1 _13982_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[22] ),
    .A2(_06818_),
    .A3(_07052_),
    .B1(_07054_),
    .C1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_07055_));
 sky130_fd_sc_hd__a221oi_1 _13983_ (.A1(_10168_),
    .A2(_06828_),
    .B1(_07051_),
    .B2(_07055_),
    .C1(_03724_),
    .Y(_07056_));
 sky130_fd_sc_hd__o21ai_0 _13984_ (.A1(_13335_),
    .A2(_04235_),
    .B1(_06765_),
    .Y(_07057_));
 sky130_fd_sc_hd__o22a_1 _13985_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[54] ),
    .A2(_06765_),
    .B1(_07056_),
    .B2(_07057_),
    .X(_01562_));
 sky130_fd_sc_hd__nand2_1 _13986_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[55] ),
    .B(_06808_),
    .Y(_07058_));
 sky130_fd_sc_hd__nand3_1 _13987_ (.A(_03724_),
    .B(_04378_),
    .C(_06765_),
    .Y(_07059_));
 sky130_fd_sc_hd__nor2_1 _13988_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[55] ),
    .B(_13488_),
    .Y(_07060_));
 sky130_fd_sc_hd__nor2_1 _13989_ (.A(net1244),
    .B(_13468_),
    .Y(_07061_));
 sky130_fd_sc_hd__nor2_1 _13990_ (.A(_07060_),
    .B(_07061_),
    .Y(_07062_));
 sky130_fd_sc_hd__nor2_1 _13991_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[23] ),
    .B(_06757_),
    .Y(_07063_));
 sky130_fd_sc_hd__o21ai_1 _13992_ (.A1(_06844_),
    .A2(_13497_),
    .B1(_07063_),
    .Y(_07064_));
 sky130_fd_sc_hd__o211ai_1 _13993_ (.A1(_13333_),
    .A2(_07062_),
    .B1(_07064_),
    .C1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_07065_));
 sky130_fd_sc_hd__a21oi_1 _13994_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net1244),
    .B1(_06770_),
    .Y(_07066_));
 sky130_fd_sc_hd__o211ai_1 _13995_ (.A1(_10810_),
    .A2(_07053_),
    .B1(_07065_),
    .C1(_07066_),
    .Y(_07067_));
 sky130_fd_sc_hd__o2111ai_1 _13996_ (.A1(_10233_),
    .A2(_06772_),
    .B1(_07067_),
    .C1(_13335_),
    .D1(_06765_),
    .Y(_07068_));
 sky130_fd_sc_hd__nand3_1 _13997_ (.A(_07058_),
    .B(_07059_),
    .C(_07068_),
    .Y(_01563_));
 sky130_fd_sc_hd__a221oi_2 _13998_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net1535),
    .B1(_07062_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(_06770_),
    .Y(_07069_));
 sky130_fd_sc_hd__nor2_1 _13999_ (.A(_13345_),
    .B(_13503_),
    .Y(_07070_));
 sky130_fd_sc_hd__mux2i_1 _14000_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[56] ),
    .A1(net1535),
    .S(_13488_),
    .Y(_07071_));
 sky130_fd_sc_hd__nand2_1 _14001_ (.A(_06818_),
    .B(_07071_),
    .Y(_07072_));
 sky130_fd_sc_hd__o311ai_4 _14002_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[24] ),
    .A2(_06818_),
    .A3(_07070_),
    .B1(_07072_),
    .C1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_07073_));
 sky130_fd_sc_hd__a221oi_4 _14003_ (.A1(_10365_),
    .A2(_06828_),
    .B1(_07069_),
    .B2(_07073_),
    .C1(_03724_),
    .Y(_07074_));
 sky130_fd_sc_hd__a311oi_1 _14004_ (.A1(_03724_),
    .A2(_04530_),
    .A3(_04531_),
    .B1(_06808_),
    .C1(_07074_),
    .Y(_07075_));
 sky130_fd_sc_hd__a21oi_1 _14005_ (.A1(_10343_),
    .A2(_06808_),
    .B1(_07075_),
    .Y(_01564_));
 sky130_fd_sc_hd__o221a_1 _14006_ (.A1(_08502_),
    .A2(_10407_),
    .B1(_07071_),
    .B2(_10810_),
    .C1(_06755_),
    .X(_07076_));
 sky130_fd_sc_hd__nor2_1 _14007_ (.A(_06869_),
    .B(_13503_),
    .Y(_07077_));
 sky130_fd_sc_hd__nor2_1 _14008_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[57] ),
    .B(_13488_),
    .Y(_07078_));
 sky130_fd_sc_hd__a21oi_1 _14009_ (.A1(_10407_),
    .A2(_13488_),
    .B1(_07078_),
    .Y(_07079_));
 sky130_fd_sc_hd__or2_0 _14010_ (.A(_06774_),
    .B(_07079_),
    .X(_07080_));
 sky130_fd_sc_hd__o311ai_2 _14011_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[25] ),
    .A2(_06757_),
    .A3(_07077_),
    .B1(_07080_),
    .C1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_07081_));
 sky130_fd_sc_hd__a221oi_2 _14012_ (.A1(_10299_),
    .A2(_06828_),
    .B1(_07076_),
    .B2(_07081_),
    .C1(_03724_),
    .Y(_07082_));
 sky130_fd_sc_hd__a21oi_1 _14013_ (.A1(_03724_),
    .A2(_04645_),
    .B1(_07082_),
    .Y(_07083_));
 sky130_fd_sc_hd__nand2_1 _14014_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[57] ),
    .B(_06808_),
    .Y(_07084_));
 sky130_fd_sc_hd__o21ai_0 _14015_ (.A1(_06808_),
    .A2(_07083_),
    .B1(_07084_),
    .Y(_01565_));
 sky130_fd_sc_hd__nand2_1 _14016_ (.A(_10865_),
    .B(net301),
    .Y(_07085_));
 sky130_fd_sc_hd__o21ai_0 _14017_ (.A1(net1062),
    .A2(_06685_),
    .B1(_07085_),
    .Y(_07086_));
 sky130_fd_sc_hd__nand2_1 _14018_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[5] ),
    .B(_10952_),
    .Y(_07087_));
 sky130_fd_sc_hd__o21ai_0 _14019_ (.A1(_10952_),
    .A2(_07086_),
    .B1(_07087_),
    .Y(_01566_));
 sky130_fd_sc_hd__nor2_1 _14020_ (.A(_10535_),
    .B(_13468_),
    .Y(_07088_));
 sky130_fd_sc_hd__a21oi_1 _14021_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[58] ),
    .A2(_13468_),
    .B1(_07088_),
    .Y(_07089_));
 sky130_fd_sc_hd__nor2_1 _14022_ (.A(_06833_),
    .B(_13503_),
    .Y(_07090_));
 sky130_fd_sc_hd__o21ai_0 _14023_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[26] ),
    .A2(_07090_),
    .B1(_06774_),
    .Y(_07091_));
 sky130_fd_sc_hd__o21ai_0 _14024_ (.A1(_06774_),
    .A2(_07089_),
    .B1(_07091_),
    .Y(_07092_));
 sky130_fd_sc_hd__a221o_1 _14025_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net167),
    .B1(_07079_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(_06770_),
    .X(_07093_));
 sky130_fd_sc_hd__a21oi_1 _14026_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .A2(_07092_),
    .B1(_07093_),
    .Y(_07094_));
 sky130_fd_sc_hd__nand2_1 _14027_ (.A(_10457_),
    .B(_06828_),
    .Y(_07095_));
 sky130_fd_sc_hd__nand3_1 _14028_ (.A(_13335_),
    .B(_06765_),
    .C(_07095_),
    .Y(_07096_));
 sky130_fd_sc_hd__nand2_1 _14029_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[58] ),
    .B(_06808_),
    .Y(_07097_));
 sky130_fd_sc_hd__nand3_1 _14030_ (.A(_03724_),
    .B(_04747_),
    .C(_06765_),
    .Y(_07098_));
 sky130_fd_sc_hd__o211ai_1 _14031_ (.A1(_07094_),
    .A2(_07096_),
    .B1(_07097_),
    .C1(_07098_),
    .Y(_01567_));
 sky130_fd_sc_hd__a21oi_1 _14032_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net687),
    .B1(_06770_),
    .Y(_07099_));
 sky130_fd_sc_hd__o21a_1 _14033_ (.A1(_10810_),
    .A2(_07089_),
    .B1(_07099_),
    .X(_07100_));
 sky130_fd_sc_hd__nor2_1 _14034_ (.A(_06844_),
    .B(_13503_),
    .Y(_07101_));
 sky130_fd_sc_hd__mux2i_2 _14035_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[59] ),
    .A1(net687),
    .S(_13488_),
    .Y(_07102_));
 sky130_fd_sc_hd__nand2_1 _14036_ (.A(_06818_),
    .B(_07102_),
    .Y(_07103_));
 sky130_fd_sc_hd__o311ai_2 _14037_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[27] ),
    .A2(_06757_),
    .A3(_07101_),
    .B1(_07103_),
    .C1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_07104_));
 sky130_fd_sc_hd__a221oi_2 _14038_ (.A1(_10493_),
    .A2(_06828_),
    .B1(_07100_),
    .B2(_07104_),
    .C1(_03724_),
    .Y(_07105_));
 sky130_fd_sc_hd__a21oi_1 _14039_ (.A1(_03724_),
    .A2(_04852_),
    .B1(_07105_),
    .Y(_07106_));
 sky130_fd_sc_hd__nand2_1 _14040_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[59] ),
    .B(_06808_),
    .Y(_07107_));
 sky130_fd_sc_hd__o21ai_0 _14041_ (.A1(_06808_),
    .A2(_07106_),
    .B1(_07107_),
    .Y(_01568_));
 sky130_fd_sc_hd__nor2_1 _14042_ (.A(_10810_),
    .B(_07102_),
    .Y(_07108_));
 sky130_fd_sc_hd__a211oi_1 _14043_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net492),
    .B1(_06770_),
    .C1(_07108_),
    .Y(_07109_));
 sky130_fd_sc_hd__nor2_1 _14044_ (.A(_13345_),
    .B(_01649_),
    .Y(_07110_));
 sky130_fd_sc_hd__mux2i_1 _14045_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[60] ),
    .A1(net493),
    .S(_13488_),
    .Y(_07111_));
 sky130_fd_sc_hd__nand2_1 _14046_ (.A(_06818_),
    .B(_07111_),
    .Y(_07112_));
 sky130_fd_sc_hd__o311ai_1 _14047_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[28] ),
    .A2(_06818_),
    .A3(_07110_),
    .B1(_07112_),
    .C1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_07113_));
 sky130_fd_sc_hd__a221oi_1 _14048_ (.A1(_10644_),
    .A2(_06828_),
    .B1(_07109_),
    .B2(_07113_),
    .C1(_03724_),
    .Y(_07114_));
 sky130_fd_sc_hd__a311oi_1 _14049_ (.A1(_03724_),
    .A2(_04970_),
    .A3(_04971_),
    .B1(_06808_),
    .C1(_07114_),
    .Y(_07115_));
 sky130_fd_sc_hd__nor2_1 _14050_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[60] ),
    .B(_06765_),
    .Y(_07116_));
 sky130_fd_sc_hd__nor2_1 _14051_ (.A(_07115_),
    .B(_07116_),
    .Y(_01569_));
 sky130_fd_sc_hd__o221a_1 _14052_ (.A1(_08502_),
    .A2(net850),
    .B1(_07111_),
    .B2(_10810_),
    .C1(_06755_),
    .X(_07117_));
 sky130_fd_sc_hd__nor2_1 _14053_ (.A(_06869_),
    .B(_01649_),
    .Y(_07118_));
 sky130_fd_sc_hd__nand2_1 _14054_ (.A(net852),
    .B(_13488_),
    .Y(_07119_));
 sky130_fd_sc_hd__o21ai_1 _14055_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[61] ),
    .A2(_13488_),
    .B1(_07119_),
    .Y(_07120_));
 sky130_fd_sc_hd__nand2_1 _14056_ (.A(_06818_),
    .B(_07120_),
    .Y(_07121_));
 sky130_fd_sc_hd__o311ai_2 _14057_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[29] ),
    .A2(_06818_),
    .A3(_07118_),
    .B1(_07121_),
    .C1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_07122_));
 sky130_fd_sc_hd__a221oi_2 _14058_ (.A1(_10557_),
    .A2(_06828_),
    .B1(_07117_),
    .B2(_07122_),
    .C1(_03724_),
    .Y(_07123_));
 sky130_fd_sc_hd__a21oi_1 _14059_ (.A1(_03724_),
    .A2(_05058_),
    .B1(_07123_),
    .Y(_07124_));
 sky130_fd_sc_hd__nand2_1 _14060_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[61] ),
    .B(_06808_),
    .Y(_07125_));
 sky130_fd_sc_hd__o21ai_0 _14061_ (.A1(_06808_),
    .A2(_07124_),
    .B1(_07125_),
    .Y(_01570_));
 sky130_fd_sc_hd__o221a_1 _14062_ (.A1(_08502_),
    .A2(_10809_),
    .B1(_07120_),
    .B2(_10810_),
    .C1(_06755_),
    .X(_07126_));
 sky130_fd_sc_hd__nor2_1 _14063_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[62] ),
    .B(_13488_),
    .Y(_07127_));
 sky130_fd_sc_hd__a21oi_1 _14064_ (.A1(_10809_),
    .A2(_13488_),
    .B1(_07127_),
    .Y(_07128_));
 sky130_fd_sc_hd__nor2_1 _14065_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[30] ),
    .B(_06818_),
    .Y(_07129_));
 sky130_fd_sc_hd__o21ai_1 _14066_ (.A1(_06833_),
    .A2(_01649_),
    .B1(_07129_),
    .Y(_07130_));
 sky130_fd_sc_hd__o211ai_1 _14067_ (.A1(_06774_),
    .A2(_07128_),
    .B1(_07130_),
    .C1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_07131_));
 sky130_fd_sc_hd__a221o_1 _14068_ (.A1(_10789_),
    .A2(_06828_),
    .B1(_07126_),
    .B2(_07131_),
    .C1(_03724_),
    .X(_07132_));
 sky130_fd_sc_hd__nor2_1 _14069_ (.A(_13335_),
    .B(_05164_),
    .Y(_07133_));
 sky130_fd_sc_hd__o21ai_0 _14070_ (.A1(_01698_),
    .A2(_05162_),
    .B1(_07133_),
    .Y(_07134_));
 sky130_fd_sc_hd__a21oi_1 _14071_ (.A1(_07132_),
    .A2(_07134_),
    .B1(_06808_),
    .Y(_07135_));
 sky130_fd_sc_hd__a21o_1 _14072_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[62] ),
    .A2(_06808_),
    .B1(_07135_),
    .X(_01571_));
 sky130_fd_sc_hd__a21oi_1 _14073_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[63] ),
    .A2(net484),
    .B1(_06774_),
    .Y(_07136_));
 sky130_fd_sc_hd__nor2_1 _14074_ (.A(_06844_),
    .B(_01649_),
    .Y(_07137_));
 sky130_fd_sc_hd__nor3_1 _14075_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[31] ),
    .B(_06818_),
    .C(_07137_),
    .Y(_07138_));
 sky130_fd_sc_hd__nor2_1 _14076_ (.A(_07136_),
    .B(_07138_),
    .Y(_07139_));
 sky130_fd_sc_hd__a221o_1 _14077_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(net481),
    .B1(_07128_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .C1(_06770_),
    .X(_07140_));
 sky130_fd_sc_hd__a21oi_1 _14078_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .A2(_07139_),
    .B1(_07140_),
    .Y(_07141_));
 sky130_fd_sc_hd__nor2_1 _14079_ (.A(_10691_),
    .B(_06772_),
    .Y(_07142_));
 sky130_fd_sc_hd__nor3_1 _14080_ (.A(_03724_),
    .B(_07141_),
    .C(_07142_),
    .Y(_07143_));
 sky130_fd_sc_hd__nor3_1 _14081_ (.A(_13335_),
    .B(_05249_),
    .C(_05250_),
    .Y(_07144_));
 sky130_fd_sc_hd__o21ai_0 _14082_ (.A1(_07143_),
    .A2(_07144_),
    .B1(_06765_),
    .Y(_07145_));
 sky130_fd_sc_hd__o21ai_0 _14083_ (.A1(_10727_),
    .A2(_06765_),
    .B1(_07145_),
    .Y(_01572_));
 sky130_fd_sc_hd__inv_1 _14084_ (.A(_05053_),
    .Y(_07146_));
 sky130_fd_sc_hd__a31oi_1 _14085_ (.A1(_07146_),
    .A2(_05155_),
    .A3(_05160_),
    .B1(_05151_),
    .Y(_07147_));
 sky130_fd_sc_hd__o22ai_1 _14086_ (.A1(_05243_),
    .A2(_05246_),
    .B1(_07147_),
    .B2(_05150_),
    .Y(_07148_));
 sky130_fd_sc_hd__nand2_1 _14087_ (.A(_05243_),
    .B(_05246_),
    .Y(_07149_));
 sky130_fd_sc_hd__nor2_1 _14088_ (.A(_05240_),
    .B(_05241_),
    .Y(_07150_));
 sky130_fd_sc_hd__nand2_1 _14089_ (.A(_05240_),
    .B(_05241_),
    .Y(_07151_));
 sky130_fd_sc_hd__o21ai_0 _14090_ (.A1(_05200_),
    .A2(_07150_),
    .B1(_07151_),
    .Y(_07152_));
 sky130_fd_sc_hd__maj3_2 _14091_ (.A(_05211_),
    .B(_05212_),
    .C(_05239_),
    .X(_07153_));
 sky130_fd_sc_hd__inv_1 _14092_ (.A(_05223_),
    .Y(_07154_));
 sky130_fd_sc_hd__inv_1 _14093_ (.A(_05237_),
    .Y(_07155_));
 sky130_fd_sc_hd__maj3_1 _14094_ (.A(_07154_),
    .B(_05225_),
    .C(_07155_),
    .X(_07156_));
 sky130_fd_sc_hd__a21o_2 _14095_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[63] ),
    .A2(net311),
    .B1(_03772_),
    .X(_07157_));
 sky130_fd_sc_hd__nor2_1 _14096_ (.A(_05092_),
    .B(_05214_),
    .Y(_07158_));
 sky130_fd_sc_hd__nor2_1 _14097_ (.A(_04049_),
    .B(_07157_),
    .Y(_07159_));
 sky130_fd_sc_hd__a211oi_1 _14098_ (.A1(_04049_),
    .A2(_07158_),
    .B1(_07159_),
    .C1(_03933_),
    .Y(_07160_));
 sky130_fd_sc_hd__nor2_1 _14099_ (.A(_04049_),
    .B(_05214_),
    .Y(_07161_));
 sky130_fd_sc_hd__a21oi_1 _14100_ (.A1(_05102_),
    .A2(_05214_),
    .B1(_07161_),
    .Y(_07162_));
 sky130_fd_sc_hd__o21a_1 _14101_ (.A1(_05092_),
    .A2(_07162_),
    .B1(_03933_),
    .X(_07163_));
 sky130_fd_sc_hd__o32ai_1 _14102_ (.A1(_05215_),
    .A2(_05104_),
    .A3(_07157_),
    .B1(_07160_),
    .B2(_07163_),
    .Y(_07164_));
 sky130_fd_sc_hd__nor2_1 _14103_ (.A(_05215_),
    .B(_07157_),
    .Y(_07165_));
 sky130_fd_sc_hd__a21oi_1 _14104_ (.A1(_04049_),
    .A2(_07165_),
    .B1(_07161_),
    .Y(_07166_));
 sky130_fd_sc_hd__nor2_1 _14105_ (.A(_03695_),
    .B(_07166_),
    .Y(_07167_));
 sky130_fd_sc_hd__a21oi_1 _14106_ (.A1(_04677_),
    .A2(_07165_),
    .B1(_07167_),
    .Y(_07168_));
 sky130_fd_sc_hd__nor2_1 _14107_ (.A(_03927_),
    .B(_07168_),
    .Y(_07169_));
 sky130_fd_sc_hd__a21oi_1 _14108_ (.A1(_03927_),
    .A2(_07164_),
    .B1(_07169_),
    .Y(_07170_));
 sky130_fd_sc_hd__xnor2_1 _14109_ (.A(_05225_),
    .B(_07170_),
    .Y(_07171_));
 sky130_fd_sc_hd__a21oi_4 _14110_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ),
    .A2(net311),
    .B1(_03772_),
    .Y(_07172_));
 sky130_fd_sc_hd__o21ai_0 _14111_ (.A1(_05215_),
    .A2(_05214_),
    .B1(_03937_),
    .Y(_07173_));
 sky130_fd_sc_hd__a21oi_1 _14112_ (.A1(_05218_),
    .A2(_07173_),
    .B1(_03941_),
    .Y(_07174_));
 sky130_fd_sc_hd__a21o_1 _14113_ (.A1(_04049_),
    .A2(_07157_),
    .B1(_07174_),
    .X(_07175_));
 sky130_fd_sc_hd__nor3_1 _14114_ (.A(_03933_),
    .B(_03937_),
    .C(_07157_),
    .Y(_07176_));
 sky130_fd_sc_hd__a21oi_1 _14115_ (.A1(_03933_),
    .A2(_07161_),
    .B1(_07176_),
    .Y(_07177_));
 sky130_fd_sc_hd__nor2_1 _14116_ (.A(_03927_),
    .B(_07177_),
    .Y(_07178_));
 sky130_fd_sc_hd__a21oi_1 _14117_ (.A1(_03927_),
    .A2(_07175_),
    .B1(_07178_),
    .Y(_07179_));
 sky130_fd_sc_hd__xnor2_1 _14118_ (.A(_07172_),
    .B(_07179_),
    .Y(_07180_));
 sky130_fd_sc_hd__xnor2_1 _14119_ (.A(_04674_),
    .B(_07180_),
    .Y(_07181_));
 sky130_fd_sc_hd__xnor2_2 _14120_ (.A(_07171_),
    .B(_07181_),
    .Y(_07182_));
 sky130_fd_sc_hd__inv_1 _14121_ (.A(_05207_),
    .Y(_07183_));
 sky130_fd_sc_hd__nand2_1 _14122_ (.A(_07183_),
    .B(_05209_),
    .Y(_07184_));
 sky130_fd_sc_hd__xor2_1 _14123_ (.A(_04272_),
    .B(_04560_),
    .X(_07185_));
 sky130_fd_sc_hd__nor2_1 _14124_ (.A(_03670_),
    .B(_05119_),
    .Y(_07186_));
 sky130_fd_sc_hd__xnor2_1 _14125_ (.A(_07185_),
    .B(_07186_),
    .Y(_07187_));
 sky130_fd_sc_hd__o211ai_1 _14126_ (.A1(_03373_),
    .A2(_05202_),
    .B1(_05026_),
    .C1(_03313_),
    .Y(_07188_));
 sky130_fd_sc_hd__nor2_1 _14127_ (.A(_03370_),
    .B(_03428_),
    .Y(_07189_));
 sky130_fd_sc_hd__a21oi_1 _14128_ (.A1(_03428_),
    .A2(_07188_),
    .B1(_07189_),
    .Y(_07190_));
 sky130_fd_sc_hd__nor2_1 _14129_ (.A(_03670_),
    .B(_05026_),
    .Y(_07191_));
 sky130_fd_sc_hd__xnor2_1 _14130_ (.A(_07191_),
    .B(_05205_),
    .Y(_07192_));
 sky130_fd_sc_hd__nor2_1 _14131_ (.A(_05201_),
    .B(_07192_),
    .Y(_07193_));
 sky130_fd_sc_hd__nand2_1 _14132_ (.A(_05201_),
    .B(_07192_),
    .Y(_07194_));
 sky130_fd_sc_hd__nor2_1 _14133_ (.A(_05133_),
    .B(_07194_),
    .Y(_07195_));
 sky130_fd_sc_hd__a21oi_1 _14134_ (.A1(_05133_),
    .A2(_07193_),
    .B1(_07195_),
    .Y(_07196_));
 sky130_fd_sc_hd__xor2_1 _14135_ (.A(_07190_),
    .B(_07196_),
    .X(_07197_));
 sky130_fd_sc_hd__xnor2_1 _14136_ (.A(_07187_),
    .B(_07197_),
    .Y(_07198_));
 sky130_fd_sc_hd__maj3_1 _14137_ (.A(_05133_),
    .B(_05122_),
    .C(_05208_),
    .X(_07199_));
 sky130_fd_sc_hd__o21ai_1 _14138_ (.A1(_07183_),
    .A2(_07199_),
    .B1(_07187_),
    .Y(_07200_));
 sky130_fd_sc_hd__and3_2 _14139_ (.A(_07184_),
    .B(_07198_),
    .C(_07200_),
    .X(_07201_));
 sky130_fd_sc_hd__a21oi_4 _14140_ (.A1(_07184_),
    .A2(_07200_),
    .B1(_07198_),
    .Y(_07202_));
 sky130_fd_sc_hd__nor2_1 _14141_ (.A(_07201_),
    .B(_07202_),
    .Y(_07203_));
 sky130_fd_sc_hd__xor2_1 _14142_ (.A(_07182_),
    .B(_07203_),
    .X(_07204_));
 sky130_fd_sc_hd__xnor2_1 _14143_ (.A(_07156_),
    .B(_07204_),
    .Y(_07205_));
 sky130_fd_sc_hd__xnor2_1 _14144_ (.A(_07153_),
    .B(_07205_),
    .Y(_07206_));
 sky130_fd_sc_hd__nand2_1 _14145_ (.A(_07152_),
    .B(_07206_),
    .Y(_07207_));
 sky130_fd_sc_hd__or2_0 _14146_ (.A(_07152_),
    .B(_07206_),
    .X(_07208_));
 sky130_fd_sc_hd__a22oi_1 _14147_ (.A1(_07148_),
    .A2(_07149_),
    .B1(_07207_),
    .B2(_07208_),
    .Y(_07209_));
 sky130_fd_sc_hd__and4_1 _14148_ (.A(_07148_),
    .B(_07149_),
    .C(_07207_),
    .D(_07208_),
    .X(_07210_));
 sky130_fd_sc_hd__o21ai_2 _14149_ (.A1(_07209_),
    .A2(_07210_),
    .B1(_02169_),
    .Y(_07211_));
 sky130_fd_sc_hd__o21ai_1 _14150_ (.A1(net445),
    .A2(_06755_),
    .B1(_13335_),
    .Y(_07212_));
 sky130_fd_sc_hd__a311o_1 _14151_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[63] ),
    .A3(net481),
    .B1(_06808_),
    .C1(_07212_),
    .X(_07213_));
 sky130_fd_sc_hd__o21ai_0 _14152_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ),
    .A2(_06765_),
    .B1(_07213_),
    .Y(_07214_));
 sky130_fd_sc_hd__a31oi_1 _14153_ (.A1(_03724_),
    .A2(_06765_),
    .A3(_07211_),
    .B1(_07214_),
    .Y(_01573_));
 sky130_fd_sc_hd__nand2_1 _14154_ (.A(_07157_),
    .B(_07172_),
    .Y(_07215_));
 sky130_fd_sc_hd__nor2_1 _14155_ (.A(_04049_),
    .B(_07172_),
    .Y(_07216_));
 sky130_fd_sc_hd__nor2_1 _14156_ (.A(_03937_),
    .B(_07215_),
    .Y(_07217_));
 sky130_fd_sc_hd__o21ai_0 _14157_ (.A1(_07216_),
    .A2(_07217_),
    .B1(_03941_),
    .Y(_07218_));
 sky130_fd_sc_hd__o21ai_0 _14158_ (.A1(_04352_),
    .A2(_07215_),
    .B1(_07218_),
    .Y(_07219_));
 sky130_fd_sc_hd__nor3_1 _14159_ (.A(_03937_),
    .B(_07157_),
    .C(_07172_),
    .Y(_07220_));
 sky130_fd_sc_hd__a211oi_1 _14160_ (.A1(_03937_),
    .A2(_07172_),
    .B1(_07220_),
    .C1(_03933_),
    .Y(_07221_));
 sky130_fd_sc_hd__nand3_1 _14161_ (.A(_04049_),
    .B(_05092_),
    .C(_07172_),
    .Y(_07222_));
 sky130_fd_sc_hd__o21ai_0 _14162_ (.A1(_04049_),
    .A2(_07172_),
    .B1(_07222_),
    .Y(_07223_));
 sky130_fd_sc_hd__a21oi_1 _14163_ (.A1(_05214_),
    .A2(_07223_),
    .B1(_03941_),
    .Y(_07224_));
 sky130_fd_sc_hd__o22ai_1 _14164_ (.A1(_05227_),
    .A2(_07215_),
    .B1(_07221_),
    .B2(_07224_),
    .Y(_07225_));
 sky130_fd_sc_hd__mux2i_1 _14165_ (.A0(_07219_),
    .A1(_07225_),
    .S(_03927_),
    .Y(_07226_));
 sky130_fd_sc_hd__nand3_1 _14166_ (.A(_03933_),
    .B(_03937_),
    .C(_05214_),
    .Y(_07227_));
 sky130_fd_sc_hd__o221ai_1 _14167_ (.A1(_03937_),
    .A2(_07172_),
    .B1(_07215_),
    .B2(_03941_),
    .C1(_07227_),
    .Y(_07228_));
 sky130_fd_sc_hd__nand3_1 _14168_ (.A(_03941_),
    .B(_04049_),
    .C(_07172_),
    .Y(_07229_));
 sky130_fd_sc_hd__nand2_1 _14169_ (.A(_03933_),
    .B(_07216_),
    .Y(_07230_));
 sky130_fd_sc_hd__a21oi_1 _14170_ (.A1(_07229_),
    .A2(_07230_),
    .B1(_03927_),
    .Y(_07231_));
 sky130_fd_sc_hd__a21oi_1 _14171_ (.A1(_03927_),
    .A2(_07228_),
    .B1(_07231_),
    .Y(_07232_));
 sky130_fd_sc_hd__a21oi_1 _14172_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ),
    .A2(net311),
    .B1(_03772_),
    .Y(_07233_));
 sky130_fd_sc_hd__xor2_1 _14173_ (.A(_07232_),
    .B(_07233_),
    .X(_07234_));
 sky130_fd_sc_hd__xnor2_1 _14174_ (.A(_07226_),
    .B(_07234_),
    .Y(_07235_));
 sky130_fd_sc_hd__inv_1 _14175_ (.A(_07170_),
    .Y(_07236_));
 sky130_fd_sc_hd__nor3_1 _14176_ (.A(_05225_),
    .B(_07236_),
    .C(_07180_),
    .Y(_07237_));
 sky130_fd_sc_hd__and3_1 _14177_ (.A(_05225_),
    .B(_07236_),
    .C(_07180_),
    .X(_07238_));
 sky130_fd_sc_hd__a211oi_1 _14178_ (.A1(_04501_),
    .A2(_07171_),
    .B1(_07237_),
    .C1(_07238_),
    .Y(_07239_));
 sky130_fd_sc_hd__xnor2_1 _14179_ (.A(_07235_),
    .B(_07239_),
    .Y(_07240_));
 sky130_fd_sc_hd__o211a_1 _14180_ (.A1(_07190_),
    .A2(_07193_),
    .B1(_05133_),
    .C1(_07187_),
    .X(_07241_));
 sky130_fd_sc_hd__a21oi_1 _14181_ (.A1(_07153_),
    .A2(_07201_),
    .B1(_07241_),
    .Y(_07242_));
 sky130_fd_sc_hd__xnor2_1 _14182_ (.A(_07240_),
    .B(_07242_),
    .Y(_07243_));
 sky130_fd_sc_hd__nor2_1 _14183_ (.A(_07182_),
    .B(_07201_),
    .Y(_07244_));
 sky130_fd_sc_hd__nor2_1 _14184_ (.A(_07202_),
    .B(_07244_),
    .Y(_07245_));
 sky130_fd_sc_hd__nor2_1 _14185_ (.A(_07153_),
    .B(_07245_),
    .Y(_07246_));
 sky130_fd_sc_hd__nand2_1 _14186_ (.A(_07182_),
    .B(_07201_),
    .Y(_07247_));
 sky130_fd_sc_hd__o31ai_1 _14187_ (.A1(_07156_),
    .A2(_07202_),
    .A3(_07244_),
    .B1(_07247_),
    .Y(_07248_));
 sky130_fd_sc_hd__nand2b_1 _14188_ (.A_N(_07182_),
    .B(_07202_),
    .Y(_07249_));
 sky130_fd_sc_hd__mux2_1 _14189_ (.A0(_07247_),
    .A1(_07249_),
    .S(_07156_),
    .X(_07250_));
 sky130_fd_sc_hd__o21ai_0 _14190_ (.A1(_07153_),
    .A2(_07249_),
    .B1(_07250_),
    .Y(_07251_));
 sky130_fd_sc_hd__a221oi_1 _14191_ (.A1(_07156_),
    .A2(_07246_),
    .B1(_07248_),
    .B2(_07153_),
    .C1(_07251_),
    .Y(_07252_));
 sky130_fd_sc_hd__xnor2_1 _14192_ (.A(_07243_),
    .B(_07252_),
    .Y(_07253_));
 sky130_fd_sc_hd__nor3_1 _14193_ (.A(_05150_),
    .B(_05195_),
    .C(_05196_),
    .Y(_07254_));
 sky130_fd_sc_hd__nor2_1 _14194_ (.A(_05151_),
    .B(_07254_),
    .Y(_07255_));
 sky130_fd_sc_hd__maj3_1 _14195_ (.A(_05243_),
    .B(_05246_),
    .C(_07255_),
    .X(_07256_));
 sky130_fd_sc_hd__nand2_1 _14196_ (.A(_07207_),
    .B(_07256_),
    .Y(_07257_));
 sky130_fd_sc_hd__nand2_1 _14197_ (.A(_07208_),
    .B(_07257_),
    .Y(_07258_));
 sky130_fd_sc_hd__xor2_1 _14198_ (.A(_07253_),
    .B(_07258_),
    .X(_07259_));
 sky130_fd_sc_hd__a21oi_1 _14199_ (.A1(_06774_),
    .A2(_06770_),
    .B1(_06808_),
    .Y(_07260_));
 sky130_fd_sc_hd__mux2i_1 _14200_ (.A0(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ),
    .A1(_07212_),
    .S(_06765_),
    .Y(_07261_));
 sky130_fd_sc_hd__a21oi_1 _14201_ (.A1(_07259_),
    .A2(_07260_),
    .B1(_07261_),
    .Y(_01574_));
 sky130_fd_sc_hd__nor2_1 _14202_ (.A(_09159_),
    .B(net301),
    .Y(_07262_));
 sky130_fd_sc_hd__a21oi_1 _14203_ (.A1(_09148_),
    .A2(net301),
    .B1(_07262_),
    .Y(_07263_));
 sky130_fd_sc_hd__nand2_1 _14204_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[6] ),
    .B(_10952_),
    .Y(_07264_));
 sky130_fd_sc_hd__o21ai_0 _14205_ (.A1(_10952_),
    .A2(_07263_),
    .B1(_07264_),
    .Y(_01575_));
 sky130_fd_sc_hd__nor2_1 _14206_ (.A(net1023),
    .B(net301),
    .Y(_07265_));
 sky130_fd_sc_hd__a21oi_1 _14207_ (.A1(_08494_),
    .A2(net301),
    .B1(_07265_),
    .Y(_07266_));
 sky130_fd_sc_hd__nand2_1 _14208_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[7] ),
    .B(_10952_),
    .Y(_07267_));
 sky130_fd_sc_hd__o21ai_0 _14209_ (.A1(_10952_),
    .A2(_07266_),
    .B1(_07267_),
    .Y(_01576_));
 sky130_fd_sc_hd__nor2_1 _14210_ (.A(_09217_),
    .B(_03369_),
    .Y(_07268_));
 sky130_fd_sc_hd__a21oi_1 _14211_ (.A1(net179),
    .A2(_03369_),
    .B1(_07268_),
    .Y(_07269_));
 sky130_fd_sc_hd__nand2_1 _14212_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[8] ),
    .B(_10952_),
    .Y(_07270_));
 sky130_fd_sc_hd__o21ai_0 _14213_ (.A1(_10952_),
    .A2(_07269_),
    .B1(_07270_),
    .Y(_01577_));
 sky130_fd_sc_hd__mux2i_1 _14214_ (.A0(_09260_),
    .A1(net180),
    .S(_03369_),
    .Y(_07271_));
 sky130_fd_sc_hd__nand2_1 _14215_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[9] ),
    .B(_10952_),
    .Y(_07272_));
 sky130_fd_sc_hd__o21ai_0 _14216_ (.A1(_10952_),
    .A2(_07271_),
    .B1(_07272_),
    .Y(_01578_));
 sky130_fd_sc_hd__nand2_1 _14217_ (.A(\load_store_unit_i.ls_fsm_cs[1] ),
    .B(\load_store_unit_i.lsu_err_q ),
    .Y(_07273_));
 sky130_fd_sc_hd__a21o_1 _14218_ (.A1(\load_store_unit_i.ls_fsm_cs[0] ),
    .A2(_07273_),
    .B1(_11204_),
    .X(_07274_));
 sky130_fd_sc_hd__xor2_1 _14219_ (.A(\load_store_unit_i.ls_fsm_cs[2] ),
    .B(\load_store_unit_i.ls_fsm_cs[1] ),
    .X(_07275_));
 sky130_fd_sc_hd__nand2_2 _14220_ (.A(_10846_),
    .B(_07275_),
    .Y(_07276_));
 sky130_fd_sc_hd__nor2_1 _14221_ (.A(net25),
    .B(_07276_),
    .Y(_07277_));
 sky130_fd_sc_hd__a21oi_2 _14222_ (.A1(_11206_),
    .A2(_07274_),
    .B1(_07277_),
    .Y(_07278_));
 sky130_fd_sc_hd__a21oi_2 _14223_ (.A1(\load_store_unit_i.ls_fsm_cs[2] ),
    .A2(_08302_),
    .B1(net26),
    .Y(_07279_));
 sky130_fd_sc_hd__nor2_8 _14224_ (.A(_07278_),
    .B(_07279_),
    .Y(_07280_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1251 ();
 sky130_fd_sc_hd__mux2_1 _14226_ (.A0(\id_stage_i.controller_i.lsu_addr_last_i[0] ),
    .A1(_10968_),
    .S(_07280_),
    .X(_01580_));
 sky130_fd_sc_hd__mux2_1 _14227_ (.A0(\id_stage_i.controller_i.lsu_addr_last_i[10] ),
    .A1(net1579),
    .S(_07280_),
    .X(_01581_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1249 ();
 sky130_fd_sc_hd__nor2_1 _14230_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[11] ),
    .B(_07280_),
    .Y(_07284_));
 sky130_fd_sc_hd__a21oi_1 _14231_ (.A1(net1590),
    .A2(_07280_),
    .B1(_07284_),
    .Y(_01582_));
 sky130_fd_sc_hd__mux2_1 _14232_ (.A0(\id_stage_i.controller_i.lsu_addr_last_i[12] ),
    .A1(net1559),
    .S(_07280_),
    .X(_01583_));
 sky130_fd_sc_hd__mux2_1 _14233_ (.A0(\id_stage_i.controller_i.lsu_addr_last_i[13] ),
    .A1(net1570),
    .S(_07280_),
    .X(_01584_));
 sky130_fd_sc_hd__mux2_1 _14234_ (.A0(\id_stage_i.controller_i.lsu_addr_last_i[14] ),
    .A1(net1273),
    .S(_07280_),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _14235_ (.A0(\id_stage_i.controller_i.lsu_addr_last_i[15] ),
    .A1(net721),
    .S(_07280_),
    .X(_01586_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1248 ();
 sky130_fd_sc_hd__mux2_1 _14237_ (.A0(\id_stage_i.controller_i.lsu_addr_last_i[16] ),
    .A1(net1581),
    .S(_07280_),
    .X(_01587_));
 sky130_fd_sc_hd__mux2_1 _14238_ (.A0(\id_stage_i.controller_i.lsu_addr_last_i[17] ),
    .A1(net1560),
    .S(_07280_),
    .X(_01588_));
 sky130_fd_sc_hd__mux2_1 _14239_ (.A0(\id_stage_i.controller_i.lsu_addr_last_i[18] ),
    .A1(net1242),
    .S(_07280_),
    .X(_01589_));
 sky130_fd_sc_hd__mux2_1 _14240_ (.A0(\id_stage_i.controller_i.lsu_addr_last_i[19] ),
    .A1(net1260),
    .S(_07280_),
    .X(_01590_));
 sky130_fd_sc_hd__mux2_1 _14241_ (.A0(\id_stage_i.controller_i.lsu_addr_last_i[1] ),
    .A1(_10970_),
    .S(_07280_),
    .X(_01591_));
 sky130_fd_sc_hd__mux2_1 _14242_ (.A0(\id_stage_i.controller_i.lsu_addr_last_i[20] ),
    .A1(net1007),
    .S(_07280_),
    .X(_01592_));
 sky130_fd_sc_hd__mux2_1 _14243_ (.A0(\id_stage_i.controller_i.lsu_addr_last_i[21] ),
    .A1(net1259),
    .S(_07280_),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_1 _14244_ (.A0(\id_stage_i.controller_i.lsu_addr_last_i[22] ),
    .A1(net1547),
    .S(_07280_),
    .X(_01594_));
 sky130_fd_sc_hd__mux2_1 _14245_ (.A0(\id_stage_i.controller_i.lsu_addr_last_i[23] ),
    .A1(net164),
    .S(_07280_),
    .X(_01595_));
 sky130_fd_sc_hd__mux2_1 _14246_ (.A0(\id_stage_i.controller_i.lsu_addr_last_i[24] ),
    .A1(net774),
    .S(_07280_),
    .X(_01596_));
 sky130_fd_sc_hd__nor2_1 _14247_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[25] ),
    .B(_07280_),
    .Y(_07286_));
 sky130_fd_sc_hd__a21oi_1 _14248_ (.A1(net684),
    .A2(_07280_),
    .B1(_07286_),
    .Y(_01597_));
 sky130_fd_sc_hd__mux2_1 _14249_ (.A0(\id_stage_i.controller_i.lsu_addr_last_i[26] ),
    .A1(net167),
    .S(_07280_),
    .X(_01598_));
 sky130_fd_sc_hd__mux2_1 _14250_ (.A0(\id_stage_i.controller_i.lsu_addr_last_i[27] ),
    .A1(net168),
    .S(_07280_),
    .X(_01599_));
 sky130_fd_sc_hd__mux2_1 _14251_ (.A0(\id_stage_i.controller_i.lsu_addr_last_i[28] ),
    .A1(net169),
    .S(_07280_),
    .X(_01600_));
 sky130_fd_sc_hd__nor2_1 _14252_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[29] ),
    .B(_07280_),
    .Y(_07287_));
 sky130_fd_sc_hd__a21oi_1 _14253_ (.A1(_10665_),
    .A2(_07280_),
    .B1(_07287_),
    .Y(_01601_));
 sky130_fd_sc_hd__mux2_1 _14254_ (.A0(\id_stage_i.controller_i.lsu_addr_last_i[2] ),
    .A1(net171),
    .S(_07280_),
    .X(_01602_));
 sky130_fd_sc_hd__nor2_1 _14255_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[30] ),
    .B(_07280_),
    .Y(_07288_));
 sky130_fd_sc_hd__a21oi_1 _14256_ (.A1(_10809_),
    .A2(_07280_),
    .B1(_07288_),
    .Y(_01603_));
 sky130_fd_sc_hd__nor2_1 _14257_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[31] ),
    .B(_07280_),
    .Y(_07289_));
 sky130_fd_sc_hd__a21oi_1 _14258_ (.A1(_13466_),
    .A2(_07280_),
    .B1(_07289_),
    .Y(_01604_));
 sky130_fd_sc_hd__mux2_1 _14259_ (.A0(\id_stage_i.controller_i.lsu_addr_last_i[3] ),
    .A1(net1525),
    .S(_07280_),
    .X(_01605_));
 sky130_fd_sc_hd__mux2_1 _14260_ (.A0(\id_stage_i.controller_i.lsu_addr_last_i[4] ),
    .A1(net175),
    .S(_07280_),
    .X(_01606_));
 sky130_fd_sc_hd__nand2_1 _14261_ (.A(net1062),
    .B(_07280_),
    .Y(_07290_));
 sky130_fd_sc_hd__o21ai_0 _14262_ (.A1(_09108_),
    .A2(_07280_),
    .B1(_07290_),
    .Y(_01607_));
 sky130_fd_sc_hd__nor2_1 _14263_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[6] ),
    .B(_07280_),
    .Y(_07291_));
 sky130_fd_sc_hd__a21oi_1 _14264_ (.A1(net1038),
    .A2(_07280_),
    .B1(_07291_),
    .Y(_01608_));
 sky130_fd_sc_hd__mux2_1 _14265_ (.A0(\id_stage_i.controller_i.lsu_addr_last_i[7] ),
    .A1(net178),
    .S(_07280_),
    .X(_01609_));
 sky130_fd_sc_hd__mux2_1 _14266_ (.A0(\id_stage_i.controller_i.lsu_addr_last_i[8] ),
    .A1(net179),
    .S(_07280_),
    .X(_01610_));
 sky130_fd_sc_hd__mux2_1 _14267_ (.A0(\id_stage_i.controller_i.lsu_addr_last_i[9] ),
    .A1(net1588),
    .S(_07280_),
    .X(_01611_));
 sky130_fd_sc_hd__nand2_1 _14268_ (.A(_08250_),
    .B(_08442_),
    .Y(_07292_));
 sky130_fd_sc_hd__nand2_1 _14269_ (.A(\load_store_unit_i.data_sign_ext_q ),
    .B(_11207_),
    .Y(_07293_));
 sky130_fd_sc_hd__o21ai_0 _14270_ (.A1(_11207_),
    .A2(_07292_),
    .B1(_07293_),
    .Y(_01612_));
 sky130_fd_sc_hd__and2_2 _14271_ (.A(net564),
    .B(_11195_),
    .X(net218));
 sky130_fd_sc_hd__mux2_1 _14272_ (.A0(net218),
    .A1(\load_store_unit_i.data_we_q ),
    .S(_11207_),
    .X(_01613_));
 sky130_fd_sc_hd__a21o_1 _14273_ (.A1(_08302_),
    .A2(_11203_),
    .B1(\load_store_unit_i.ls_fsm_cs[2] ),
    .X(_07294_));
 sky130_fd_sc_hd__a21oi_1 _14274_ (.A1(\load_store_unit_i.ls_fsm_cs[1] ),
    .A2(_10846_),
    .B1(net26),
    .Y(_07295_));
 sky130_fd_sc_hd__or2_2 _14275_ (.A(net677),
    .B(_08214_),
    .X(_07296_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1247 ();
 sky130_fd_sc_hd__a21oi_1 _14277_ (.A1(net491),
    .A2(_10970_),
    .B1(_07296_),
    .Y(_07298_));
 sky130_fd_sc_hd__nor2b_1 _14278_ (.A(_07298_),
    .B_N(_10968_),
    .Y(_07299_));
 sky130_fd_sc_hd__a21oi_2 _14279_ (.A1(_10970_),
    .A2(_07296_),
    .B1(_07299_),
    .Y(_07300_));
 sky130_fd_sc_hd__o21ai_0 _14280_ (.A1(\load_store_unit_i.ls_fsm_cs[2] ),
    .A2(_08302_),
    .B1(_07300_),
    .Y(_07301_));
 sky130_fd_sc_hd__nand2_1 _14281_ (.A(\load_store_unit_i.ls_fsm_cs[1] ),
    .B(_11206_),
    .Y(_07302_));
 sky130_fd_sc_hd__nand2_1 _14282_ (.A(_07301_),
    .B(_07302_),
    .Y(_07303_));
 sky130_fd_sc_hd__o21ai_0 _14283_ (.A1(_07294_),
    .A2(_07295_),
    .B1(\load_store_unit_i.handle_misaligned_q ),
    .Y(_07304_));
 sky130_fd_sc_hd__o31ai_1 _14284_ (.A1(_07294_),
    .A2(_07295_),
    .A3(_07303_),
    .B1(_07304_),
    .Y(_01614_));
 sky130_fd_sc_hd__inv_1 _14285_ (.A(\load_store_unit_i.ls_fsm_cs[0] ),
    .Y(_07305_));
 sky130_fd_sc_hd__a21oi_1 _14286_ (.A1(\load_store_unit_i.ls_fsm_cs[1] ),
    .A2(net59),
    .B1(_11204_),
    .Y(_07306_));
 sky130_fd_sc_hd__a211oi_1 _14287_ (.A1(_07305_),
    .A2(_07306_),
    .B1(net26),
    .C1(\load_store_unit_i.ls_fsm_cs[2] ),
    .Y(_01615_));
 sky130_fd_sc_hd__inv_1 _14288_ (.A(\load_store_unit_i.ls_fsm_cs[1] ),
    .Y(_07307_));
 sky130_fd_sc_hd__nor2b_1 _14289_ (.A(\load_store_unit_i.ls_fsm_cs[0] ),
    .B_N(_07300_),
    .Y(_07308_));
 sky130_fd_sc_hd__inv_2 _14290_ (.A(_07294_),
    .Y(net185));
 sky130_fd_sc_hd__o21ai_0 _14291_ (.A1(net26),
    .A2(_07308_),
    .B1(net185),
    .Y(_07309_));
 sky130_fd_sc_hd__a22oi_1 _14292_ (.A1(net59),
    .A2(_07294_),
    .B1(_07300_),
    .B2(net26),
    .Y(_07310_));
 sky130_fd_sc_hd__a21oi_1 _14293_ (.A1(\load_store_unit_i.ls_fsm_cs[1] ),
    .A2(net26),
    .B1(\load_store_unit_i.ls_fsm_cs[2] ),
    .Y(_07311_));
 sky130_fd_sc_hd__o21ai_0 _14294_ (.A1(\load_store_unit_i.ls_fsm_cs[0] ),
    .A2(_07310_),
    .B1(_07311_),
    .Y(_07312_));
 sky130_fd_sc_hd__a21oi_1 _14295_ (.A1(_07307_),
    .A2(_07309_),
    .B1(_07312_),
    .Y(_01616_));
 sky130_fd_sc_hd__mux2i_1 _14296_ (.A0(\load_store_unit_i.ls_fsm_cs[2] ),
    .A1(_11206_),
    .S(\load_store_unit_i.ls_fsm_cs[1] ),
    .Y(_07313_));
 sky130_fd_sc_hd__nor3_1 _14297_ (.A(\load_store_unit_i.ls_fsm_cs[0] ),
    .B(net59),
    .C(_07313_),
    .Y(_01617_));
 sky130_fd_sc_hd__nor2_1 _14298_ (.A(\load_store_unit_i.ls_fsm_cs[2] ),
    .B(_07306_),
    .Y(_07314_));
 sky130_fd_sc_hd__a31oi_1 _14299_ (.A1(\load_store_unit_i.ls_fsm_cs[2] ),
    .A2(_07307_),
    .A3(net59),
    .B1(_07314_),
    .Y(_07315_));
 sky130_fd_sc_hd__nand2_1 _14300_ (.A(net25),
    .B(_07275_),
    .Y(_07316_));
 sky130_fd_sc_hd__o21ai_0 _14301_ (.A1(\load_store_unit_i.ls_fsm_cs[0] ),
    .A2(_07315_),
    .B1(\load_store_unit_i.lsu_err_q ),
    .Y(_07317_));
 sky130_fd_sc_hd__o31ai_1 _14302_ (.A1(\load_store_unit_i.ls_fsm_cs[0] ),
    .A2(_07315_),
    .A3(_07316_),
    .B1(_07317_),
    .Y(_01618_));
 sky130_fd_sc_hd__mux2_1 _14303_ (.A0(_10968_),
    .A1(\load_store_unit_i.rdata_offset_q[0] ),
    .S(_11207_),
    .X(_01619_));
 sky130_fd_sc_hd__nand2_1 _14304_ (.A(\load_store_unit_i.rdata_offset_q[1] ),
    .B(_11207_),
    .Y(_07318_));
 sky130_fd_sc_hd__o21ai_0 _14305_ (.A1(_13394_),
    .A2(_11207_),
    .B1(_07318_),
    .Y(_01620_));
 sky130_fd_sc_hd__nor2_8 _14306_ (.A(\load_store_unit_i.data_we_q ),
    .B(_07276_),
    .Y(_07319_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1246 ();
 sky130_fd_sc_hd__mux2_1 _14308_ (.A0(\load_store_unit_i.rdata_q[8] ),
    .A1(net57),
    .S(_07319_),
    .X(_01621_));
 sky130_fd_sc_hd__mux2_1 _14309_ (.A0(\load_store_unit_i.rdata_q[18] ),
    .A1(net36),
    .S(_07319_),
    .X(_01622_));
 sky130_fd_sc_hd__mux2_1 _14310_ (.A0(\load_store_unit_i.rdata_q[19] ),
    .A1(net37),
    .S(_07319_),
    .X(_01623_));
 sky130_fd_sc_hd__mux2_1 _14311_ (.A0(\load_store_unit_i.rdata_q[20] ),
    .A1(net39),
    .S(_07319_),
    .X(_01624_));
 sky130_fd_sc_hd__mux2_1 _14312_ (.A0(\load_store_unit_i.rdata_q[21] ),
    .A1(net40),
    .S(_07319_),
    .X(_01625_));
 sky130_fd_sc_hd__mux2_1 _14313_ (.A0(\load_store_unit_i.rdata_q[22] ),
    .A1(net41),
    .S(_07319_),
    .X(_01626_));
 sky130_fd_sc_hd__mux2_1 _14314_ (.A0(\load_store_unit_i.rdata_q[23] ),
    .A1(net42),
    .S(_07319_),
    .X(_01627_));
 sky130_fd_sc_hd__mux2_1 _14315_ (.A0(\load_store_unit_i.rdata_q[24] ),
    .A1(net43),
    .S(_07319_),
    .X(_01628_));
 sky130_fd_sc_hd__mux2_1 _14316_ (.A0(\load_store_unit_i.rdata_q[25] ),
    .A1(net44),
    .S(_07319_),
    .X(_01629_));
 sky130_fd_sc_hd__mux2_1 _14317_ (.A0(\load_store_unit_i.rdata_q[26] ),
    .A1(net45),
    .S(_07319_),
    .X(_01630_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1245 ();
 sky130_fd_sc_hd__mux2_1 _14319_ (.A0(\load_store_unit_i.rdata_q[27] ),
    .A1(net46),
    .S(_07319_),
    .X(_01631_));
 sky130_fd_sc_hd__mux2_1 _14320_ (.A0(\load_store_unit_i.rdata_q[9] ),
    .A1(net58),
    .S(_07319_),
    .X(_01632_));
 sky130_fd_sc_hd__mux2_1 _14321_ (.A0(\load_store_unit_i.rdata_q[28] ),
    .A1(net47),
    .S(_07319_),
    .X(_01633_));
 sky130_fd_sc_hd__mux2_1 _14322_ (.A0(\load_store_unit_i.rdata_q[29] ),
    .A1(net48),
    .S(_07319_),
    .X(_01634_));
 sky130_fd_sc_hd__mux2_1 _14323_ (.A0(\load_store_unit_i.rdata_q[30] ),
    .A1(net50),
    .S(_07319_),
    .X(_01635_));
 sky130_fd_sc_hd__mux2_1 _14324_ (.A0(\load_store_unit_i.rdata_q[31] ),
    .A1(net51),
    .S(_07319_),
    .X(_01636_));
 sky130_fd_sc_hd__mux2_1 _14325_ (.A0(\load_store_unit_i.rdata_q[10] ),
    .A1(net28),
    .S(_07319_),
    .X(_01637_));
 sky130_fd_sc_hd__mux2_1 _14326_ (.A0(\load_store_unit_i.rdata_q[11] ),
    .A1(net29),
    .S(_07319_),
    .X(_01638_));
 sky130_fd_sc_hd__mux2_1 _14327_ (.A0(\load_store_unit_i.rdata_q[12] ),
    .A1(net30),
    .S(_07319_),
    .X(_01639_));
 sky130_fd_sc_hd__mux2_1 _14328_ (.A0(\load_store_unit_i.rdata_q[13] ),
    .A1(net31),
    .S(_07319_),
    .X(_01640_));
 sky130_fd_sc_hd__mux2_1 _14329_ (.A0(\load_store_unit_i.rdata_q[14] ),
    .A1(net32),
    .S(_07319_),
    .X(_01641_));
 sky130_fd_sc_hd__mux2_1 _14330_ (.A0(\load_store_unit_i.rdata_q[15] ),
    .A1(net33),
    .S(_07319_),
    .X(_01642_));
 sky130_fd_sc_hd__mux2_1 _14331_ (.A0(\load_store_unit_i.rdata_q[16] ),
    .A1(net34),
    .S(_07319_),
    .X(_01643_));
 sky130_fd_sc_hd__mux2_1 _14332_ (.A0(\load_store_unit_i.rdata_q[17] ),
    .A1(net35),
    .S(_07319_),
    .X(_01644_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1244 ();
 sky130_fd_sc_hd__nand2_1 _14334_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .Y(_07323_));
 sky130_fd_sc_hd__nand3_1 _14335_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .B(_11126_),
    .C(net94),
    .Y(_07324_));
 sky130_fd_sc_hd__nand2b_1 _14336_ (.A_N(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ),
    .B(\cs_registers_i.pc_if_i[1] ),
    .Y(_07325_));
 sky130_fd_sc_hd__a21oi_1 _14337_ (.A1(_07323_),
    .A2(_07324_),
    .B1(_07325_),
    .Y(_01579_));
 sky130_fd_sc_hd__nor2_1 _14338_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .B(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .Y(_07326_));
 sky130_fd_sc_hd__or3_1 _14339_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .B(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .C(_07326_),
    .X(_07327_));
 sky130_fd_sc_hd__nor2_1 _14340_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .Y(_07328_));
 sky130_fd_sc_hd__nor2_1 _14341_ (.A(_11126_),
    .B(_07328_),
    .Y(_07329_));
 sky130_fd_sc_hd__a2111oi_4 _14342_ (.A1(_10996_),
    .A2(_11004_),
    .B1(_11011_),
    .C1(_11034_),
    .D1(_11042_),
    .Y(_07330_));
 sky130_fd_sc_hd__a221oi_4 _14343_ (.A1(_08106_),
    .A2(_07327_),
    .B1(_07329_),
    .B2(net293),
    .C1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .Y(_07331_));
 sky130_fd_sc_hd__nor2_2 _14344_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(_07331_),
    .Y(_07332_));
 sky130_fd_sc_hd__nor4b_1 _14345_ (.A(\load_store_unit_i.ls_fsm_cs[2] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .C(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .D_N(_08302_),
    .Y(_07333_));
 sky130_fd_sc_hd__o21ai_1 _14346_ (.A1(\cs_registers_i.debug_mode_i ),
    .A2(_06647_),
    .B1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .Y(_07334_));
 sky130_fd_sc_hd__nand4_1 _14347_ (.A(_11162_),
    .B(_07332_),
    .C(_07333_),
    .D(_07334_),
    .Y(core_busy_d));
 sky130_fd_sc_hd__and2_1 _14348_ (.A(clknet_1_0__leaf_clk_i),
    .B(\core_clock_gate_i.en_latch ),
    .X(clk));
 sky130_fd_sc_hd__nand2_1 _14349_ (.A(\load_store_unit_i.handle_misaligned_q ),
    .B(_07296_),
    .Y(_07335_));
 sky130_fd_sc_hd__o21ai_1 _14350_ (.A1(net491),
    .A2(_07296_),
    .B1(\load_store_unit_i.handle_misaligned_q ),
    .Y(_07336_));
 sky130_fd_sc_hd__nor2_1 _14351_ (.A(_10971_),
    .B(_07336_),
    .Y(_07337_));
 sky130_fd_sc_hd__a21o_2 _14352_ (.A1(_10971_),
    .A2(_07335_),
    .B1(_07337_),
    .X(net181));
 sky130_fd_sc_hd__nor2_1 _14353_ (.A(net491),
    .B(_07296_),
    .Y(_07338_));
 sky130_fd_sc_hd__nand2_1 _14354_ (.A(_10968_),
    .B(_07338_),
    .Y(_07339_));
 sky130_fd_sc_hd__o21ai_0 _14355_ (.A1(\load_store_unit_i.handle_misaligned_q ),
    .A2(_07338_),
    .B1(_07339_),
    .Y(_07340_));
 sky130_fd_sc_hd__nand2_1 _14356_ (.A(_13394_),
    .B(_07340_),
    .Y(_07341_));
 sky130_fd_sc_hd__o21ai_4 _14357_ (.A1(_13394_),
    .A2(_07335_),
    .B1(_07341_),
    .Y(net182));
 sky130_fd_sc_hd__a21oi_1 _14358_ (.A1(net491),
    .A2(_10968_),
    .B1(_07296_),
    .Y(_07342_));
 sky130_fd_sc_hd__nand2_1 _14359_ (.A(_10968_),
    .B(_07335_),
    .Y(_07343_));
 sky130_fd_sc_hd__o211ai_2 _14360_ (.A1(_10968_),
    .A2(_07336_),
    .B1(_07343_),
    .C1(_10970_),
    .Y(_07344_));
 sky130_fd_sc_hd__o31ai_4 _14361_ (.A1(\load_store_unit_i.handle_misaligned_q ),
    .A2(_10970_),
    .A3(_07342_),
    .B1(_07344_),
    .Y(net183));
 sky130_fd_sc_hd__o22ai_4 _14362_ (.A1(\load_store_unit_i.handle_misaligned_q ),
    .A2(_07298_),
    .B1(_07339_),
    .B2(_13394_),
    .Y(net184));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1243 ();
 sky130_fd_sc_hd__nand2_1 _14364_ (.A(_08948_),
    .B(net275),
    .Y(_07346_));
 sky130_fd_sc_hd__o21ai_4 _14365_ (.A1(_01711_),
    .A2(net275),
    .B1(_07346_),
    .Y(_07347_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1242 ();
 sky130_fd_sc_hd__nor2_1 _14367_ (.A(_09217_),
    .B(net276),
    .Y(_07349_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1241 ();
 sky130_fd_sc_hd__nor2_1 _14369_ (.A(net1212),
    .B(net287),
    .Y(_07351_));
 sky130_fd_sc_hd__nor2_2 _14370_ (.A(_07349_),
    .B(_07351_),
    .Y(_07352_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1240 ();
 sky130_fd_sc_hd__mux2i_1 _14372_ (.A0(_07347_),
    .A1(_07352_),
    .S(net288),
    .Y(net186));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1239 ();
 sky130_fd_sc_hd__mux2i_1 _14374_ (.A0(net916),
    .A1(_10437_),
    .S(net286),
    .Y(_07355_));
 sky130_fd_sc_hd__nand2_1 _14375_ (.A(net1049),
    .B(net286),
    .Y(_07356_));
 sky130_fd_sc_hd__o21ai_4 _14376_ (.A1(_08795_),
    .A2(net286),
    .B1(_07356_),
    .Y(_07357_));
 sky130_fd_sc_hd__mux2i_1 _14377_ (.A0(_07355_),
    .A1(_07357_),
    .S(net289),
    .Y(net187));
 sky130_fd_sc_hd__nand2_1 _14378_ (.A(net932),
    .B(net275),
    .Y(_07358_));
 sky130_fd_sc_hd__o21ai_0 _14379_ (.A1(_10522_),
    .A2(net275),
    .B1(_07358_),
    .Y(_07359_));
 sky130_fd_sc_hd__nand2_1 _14380_ (.A(net746),
    .B(net286),
    .Y(_07360_));
 sky130_fd_sc_hd__nand2_1 _14381_ (.A(net785),
    .B(net275),
    .Y(_07361_));
 sky130_fd_sc_hd__nand2_1 _14382_ (.A(_07360_),
    .B(_07361_),
    .Y(_07362_));
 sky130_fd_sc_hd__mux2i_1 _14383_ (.A0(_07359_),
    .A1(_07362_),
    .S(net289),
    .Y(net188));
 sky130_fd_sc_hd__nand2_1 _14384_ (.A(_10620_),
    .B(net286),
    .Y(_07363_));
 sky130_fd_sc_hd__o21ai_0 _14385_ (.A1(_09524_),
    .A2(net286),
    .B1(_07363_),
    .Y(_07364_));
 sky130_fd_sc_hd__nand2_1 _14386_ (.A(net476),
    .B(net275),
    .Y(_07365_));
 sky130_fd_sc_hd__o21ai_4 _14387_ (.A1(_10040_),
    .A2(net275),
    .B1(_07365_),
    .Y(_07366_));
 sky130_fd_sc_hd__mux2i_1 _14388_ (.A0(_07364_),
    .A1(_07366_),
    .S(net289),
    .Y(net189));
 sky130_fd_sc_hd__nand2_1 _14389_ (.A(_09486_),
    .B(net276),
    .Y(_07367_));
 sky130_fd_sc_hd__o21ai_4 _14390_ (.A1(_10590_),
    .A2(net276),
    .B1(_07367_),
    .Y(_07368_));
 sky130_fd_sc_hd__nand2_1 _14391_ (.A(_10865_),
    .B(net276),
    .Y(_07369_));
 sky130_fd_sc_hd__o21ai_4 _14392_ (.A1(_10110_),
    .A2(net276),
    .B1(_07369_),
    .Y(_07370_));
 sky130_fd_sc_hd__mux2i_1 _14393_ (.A0(_07368_),
    .A1(_07370_),
    .S(net288),
    .Y(net190));
 sky130_fd_sc_hd__mux2i_1 _14394_ (.A0(net1144),
    .A1(_10792_),
    .S(net286),
    .Y(_07371_));
 sky130_fd_sc_hd__mux2i_1 _14395_ (.A0(net800),
    .A1(_10202_),
    .S(net286),
    .Y(_07372_));
 sky130_fd_sc_hd__mux2i_1 _14396_ (.A0(_07371_),
    .A1(_07372_),
    .S(net289),
    .Y(net191));
 sky130_fd_sc_hd__mux2i_1 _14397_ (.A0(net979),
    .A1(_10721_),
    .S(net286),
    .Y(_07373_));
 sky130_fd_sc_hd__mux2i_1 _14398_ (.A0(_08494_),
    .A1(net1081),
    .S(net286),
    .Y(_07374_));
 sky130_fd_sc_hd__mux2i_1 _14399_ (.A0(_07373_),
    .A1(_07374_),
    .S(net289),
    .Y(net192));
 sky130_fd_sc_hd__nand2_1 _14400_ (.A(_08948_),
    .B(net287),
    .Y(_07375_));
 sky130_fd_sc_hd__o21ai_4 _14401_ (.A1(net1190),
    .A2(net287),
    .B1(_07375_),
    .Y(_07376_));
 sky130_fd_sc_hd__nand2_1 _14402_ (.A(net1212),
    .B(net287),
    .Y(_07377_));
 sky130_fd_sc_hd__nand2_1 _14403_ (.A(_09217_),
    .B(net276),
    .Y(_07378_));
 sky130_fd_sc_hd__nand2_2 _14404_ (.A(_07377_),
    .B(_07378_),
    .Y(_07379_));
 sky130_fd_sc_hd__mux2i_1 _14405_ (.A0(_07376_),
    .A1(_07379_),
    .S(net288),
    .Y(net193));
 sky130_fd_sc_hd__nand2_1 _14406_ (.A(net699),
    .B(net287),
    .Y(_07380_));
 sky130_fd_sc_hd__o21ai_4 _14407_ (.A1(net1272),
    .A2(net287),
    .B1(_07380_),
    .Y(_07381_));
 sky130_fd_sc_hd__nand2_1 _14408_ (.A(_02619_),
    .B(net276),
    .Y(_07382_));
 sky130_fd_sc_hd__o21ai_2 _14409_ (.A1(_10332_),
    .A2(net276),
    .B1(_07382_),
    .Y(_07383_));
 sky130_fd_sc_hd__mux2i_1 _14410_ (.A0(_07381_),
    .A1(_07383_),
    .S(net288),
    .Y(net194));
 sky130_fd_sc_hd__nand2_1 _14411_ (.A(net1049),
    .B(net275),
    .Y(_07384_));
 sky130_fd_sc_hd__o21ai_4 _14412_ (.A1(_08795_),
    .A2(net275),
    .B1(_07384_),
    .Y(_07385_));
 sky130_fd_sc_hd__mux2i_1 _14413_ (.A0(_07385_),
    .A1(_07355_),
    .S(net289),
    .Y(net195));
 sky130_fd_sc_hd__nand2_1 _14414_ (.A(net785),
    .B(net286),
    .Y(_07386_));
 sky130_fd_sc_hd__nand2_1 _14415_ (.A(net746),
    .B(net275),
    .Y(_07387_));
 sky130_fd_sc_hd__nand2_1 _14416_ (.A(_07386_),
    .B(_07387_),
    .Y(_07388_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1238 ();
 sky130_fd_sc_hd__mux2i_1 _14418_ (.A0(_07388_),
    .A1(_07359_),
    .S(net289),
    .Y(net196));
 sky130_fd_sc_hd__nand2_1 _14419_ (.A(net699),
    .B(net276),
    .Y(_07390_));
 sky130_fd_sc_hd__o21ai_4 _14420_ (.A1(net1272),
    .A2(net276),
    .B1(_07390_),
    .Y(_07391_));
 sky130_fd_sc_hd__nand2_1 _14421_ (.A(_02619_),
    .B(net287),
    .Y(_07392_));
 sky130_fd_sc_hd__o21ai_2 _14422_ (.A1(_10332_),
    .A2(net287),
    .B1(_07392_),
    .Y(_07393_));
 sky130_fd_sc_hd__mux2i_1 _14423_ (.A0(_07391_),
    .A1(_07393_),
    .S(net288),
    .Y(net197));
 sky130_fd_sc_hd__nand2_1 _14424_ (.A(net477),
    .B(net286),
    .Y(_07394_));
 sky130_fd_sc_hd__o21ai_4 _14425_ (.A1(_10040_),
    .A2(net286),
    .B1(_07394_),
    .Y(_07395_));
 sky130_fd_sc_hd__mux2i_1 _14426_ (.A0(_07395_),
    .A1(_07364_),
    .S(net289),
    .Y(net198));
 sky130_fd_sc_hd__nand2_1 _14427_ (.A(_10865_),
    .B(net287),
    .Y(_07396_));
 sky130_fd_sc_hd__o21ai_4 _14428_ (.A1(_10110_),
    .A2(net287),
    .B1(_07396_),
    .Y(_07397_));
 sky130_fd_sc_hd__mux2i_1 _14429_ (.A0(_07397_),
    .A1(_07368_),
    .S(net288),
    .Y(net199));
 sky130_fd_sc_hd__mux2i_1 _14430_ (.A0(net800),
    .A1(_10202_),
    .S(net275),
    .Y(_07398_));
 sky130_fd_sc_hd__mux2i_1 _14431_ (.A0(_07398_),
    .A1(_07371_),
    .S(net289),
    .Y(net200));
 sky130_fd_sc_hd__mux2i_1 _14432_ (.A0(_08494_),
    .A1(net1081),
    .S(net275),
    .Y(_07399_));
 sky130_fd_sc_hd__mux2i_1 _14433_ (.A0(_07399_),
    .A1(_07373_),
    .S(net289),
    .Y(net201));
 sky130_fd_sc_hd__mux2i_1 _14434_ (.A0(_07352_),
    .A1(_07376_),
    .S(net288),
    .Y(net202));
 sky130_fd_sc_hd__mux2i_1 _14435_ (.A0(_07393_),
    .A1(_07381_),
    .S(net288),
    .Y(net203));
 sky130_fd_sc_hd__mux2i_1 _14436_ (.A0(net916),
    .A1(_10437_),
    .S(net275),
    .Y(_07400_));
 sky130_fd_sc_hd__mux2i_1 _14437_ (.A0(_07400_),
    .A1(_07385_),
    .S(net289),
    .Y(net204));
 sky130_fd_sc_hd__nand2_1 _14438_ (.A(net932),
    .B(net286),
    .Y(_07401_));
 sky130_fd_sc_hd__o21ai_0 _14439_ (.A1(_10522_),
    .A2(net286),
    .B1(_07401_),
    .Y(_07402_));
 sky130_fd_sc_hd__mux2i_1 _14440_ (.A0(_07402_),
    .A1(_07388_),
    .S(net289),
    .Y(net205));
 sky130_fd_sc_hd__nor2_1 _14441_ (.A(_10620_),
    .B(net286),
    .Y(_07403_));
 sky130_fd_sc_hd__a21oi_1 _14442_ (.A1(_09524_),
    .A2(net286),
    .B1(_07403_),
    .Y(_07404_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1237 ();
 sky130_fd_sc_hd__mux2i_1 _14444_ (.A0(_07404_),
    .A1(_07395_),
    .S(net289),
    .Y(net206));
 sky130_fd_sc_hd__nand2_1 _14445_ (.A(_09486_),
    .B(net287),
    .Y(_07406_));
 sky130_fd_sc_hd__o21ai_4 _14446_ (.A1(_10590_),
    .A2(net287),
    .B1(_07406_),
    .Y(_07407_));
 sky130_fd_sc_hd__mux2i_1 _14447_ (.A0(_07407_),
    .A1(_07397_),
    .S(net288),
    .Y(net207));
 sky130_fd_sc_hd__mux2i_1 _14448_ (.A0(_07357_),
    .A1(_07400_),
    .S(net289),
    .Y(net208));
 sky130_fd_sc_hd__mux2i_1 _14449_ (.A0(net1144),
    .A1(_10792_),
    .S(net275),
    .Y(_07408_));
 sky130_fd_sc_hd__mux2i_1 _14450_ (.A0(_07408_),
    .A1(_07398_),
    .S(net289),
    .Y(net209));
 sky130_fd_sc_hd__mux2i_1 _14451_ (.A0(net979),
    .A1(_10721_),
    .S(net275),
    .Y(_07409_));
 sky130_fd_sc_hd__mux2i_1 _14452_ (.A0(_07409_),
    .A1(_07399_),
    .S(net289),
    .Y(net210));
 sky130_fd_sc_hd__mux2i_1 _14453_ (.A0(_07362_),
    .A1(_07402_),
    .S(net289),
    .Y(net211));
 sky130_fd_sc_hd__mux2i_1 _14454_ (.A0(_07366_),
    .A1(_07404_),
    .S(net289),
    .Y(net212));
 sky130_fd_sc_hd__mux2i_1 _14455_ (.A0(_07370_),
    .A1(_07407_),
    .S(net288),
    .Y(net213));
 sky130_fd_sc_hd__mux2i_1 _14456_ (.A0(_07372_),
    .A1(_07408_),
    .S(net289),
    .Y(net214));
 sky130_fd_sc_hd__mux2i_1 _14457_ (.A0(_07374_),
    .A1(_07409_),
    .S(net289),
    .Y(net215));
 sky130_fd_sc_hd__mux2i_1 _14458_ (.A0(_07379_),
    .A1(_07347_),
    .S(net288),
    .Y(net216));
 sky130_fd_sc_hd__mux2i_1 _14459_ (.A0(_07383_),
    .A1(_07391_),
    .S(net288),
    .Y(net217));
 sky130_fd_sc_hd__inv_1 _14460_ (.A(net94),
    .Y(_07410_));
 sky130_fd_sc_hd__o21ai_0 _14461_ (.A1(_07410_),
    .A2(_11135_),
    .B1(_11126_),
    .Y(_07411_));
 sky130_fd_sc_hd__nand2_1 _14462_ (.A(\cs_registers_i.pc_if_i[1] ),
    .B(_07411_),
    .Y(_07412_));
 sky130_fd_sc_hd__a211oi_1 _14463_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .A2(_11137_),
    .B1(_07325_),
    .C1(_11126_),
    .Y(_07413_));
 sky130_fd_sc_hd__a21oi_1 _14464_ (.A1(_11136_),
    .A2(_07412_),
    .B1(_07413_),
    .Y(\if_stage_i.fetch_err ));
 sky130_fd_sc_hd__inv_1 _14465_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .Y(_07414_));
 sky130_fd_sc_hd__nand2_1 _14466_ (.A(net95),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ),
    .Y(_07415_));
 sky130_fd_sc_hd__o21ai_0 _14467_ (.A1(net128),
    .A2(net1026),
    .B1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .Y(_07416_));
 sky130_fd_sc_hd__nand3_1 _14468_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .B(net95),
    .C(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ),
    .Y(_07417_));
 sky130_fd_sc_hd__a21oi_1 _14469_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .A2(net1026),
    .B1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1] ),
    .Y(_07418_));
 sky130_fd_sc_hd__nand2_1 _14470_ (.A(_07417_),
    .B(_07418_),
    .Y(_07419_));
 sky130_fd_sc_hd__nor2_1 _14471_ (.A(_11130_),
    .B(_07419_),
    .Y(_07420_));
 sky130_fd_sc_hd__a31oi_1 _14472_ (.A1(_07414_),
    .A2(_07415_),
    .A3(_07416_),
    .B1(_07420_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ));
 sky130_fd_sc_hd__and2_0 _14473_ (.A(_11130_),
    .B(_07419_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1236 ();
 sky130_fd_sc_hd__a21oi_2 _14475_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .A2(_10996_),
    .B1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .Y(_07422_));
 sky130_fd_sc_hd__o21ai_4 _14476_ (.A1(_08106_),
    .A2(_07422_),
    .B1(_11009_),
    .Y(_07423_));
 sky130_fd_sc_hd__nor2_1 _14477_ (.A(net1),
    .B(_07423_),
    .Y(_07424_));
 sky130_fd_sc_hd__o21a_4 _14478_ (.A1(_08106_),
    .A2(_07422_),
    .B1(_11009_),
    .X(_07425_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1235 ();
 sky130_fd_sc_hd__nor4_1 _14480_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .B(\id_stage_i.controller_i.store_err_q ),
    .C(\id_stage_i.controller_i.exc_req_q ),
    .D(\id_stage_i.controller_i.load_err_q ),
    .Y(_07427_));
 sky130_fd_sc_hd__o21ai_4 _14481_ (.A1(_10945_),
    .A2(_07427_),
    .B1(_11009_),
    .Y(_07428_));
 sky130_fd_sc_hd__nand2_2 _14482_ (.A(\cs_registers_i.debug_mode_i ),
    .B(_12469_),
    .Y(_07429_));
 sky130_fd_sc_hd__and3_4 _14483_ (.A(_11009_),
    .B(_07428_),
    .C(_07429_),
    .X(_07430_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1234 ();
 sky130_fd_sc_hd__nand2_1 _14485_ (.A(\cs_registers_i.csr_mtvec_o[10] ),
    .B(_07430_),
    .Y(_07432_));
 sky130_fd_sc_hd__nor2_8 _14486_ (.A(_10941_),
    .B(_12451_),
    .Y(_07433_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1233 ();
 sky130_fd_sc_hd__a22oi_1 _14488_ (.A1(\cs_registers_i.csr_mepc_o[10] ),
    .A2(_12455_),
    .B1(_07433_),
    .B2(\cs_registers_i.csr_depc_o[10] ),
    .Y(_07435_));
 sky130_fd_sc_hd__nand2_1 _14489_ (.A(_07432_),
    .B(_07435_),
    .Y(_07436_));
 sky130_fd_sc_hd__a211oi_2 _14490_ (.A1(net319),
    .A2(net1578),
    .B1(_07425_),
    .C1(_07436_),
    .Y(_07437_));
 sky130_fd_sc_hd__nand2_1 _14491_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ),
    .B(net291),
    .Y(_07438_));
 sky130_fd_sc_hd__o31ai_1 _14492_ (.A1(net291),
    .A2(_07424_),
    .A3(_07437_),
    .B1(_07438_),
    .Y(_07439_));
 sky130_fd_sc_hd__a221oi_2 _14493_ (.A1(\cs_registers_i.csr_mepc_o[7] ),
    .A2(_12455_),
    .B1(_07433_),
    .B2(\cs_registers_i.csr_depc_o[7] ),
    .C1(_07425_),
    .Y(_07440_));
 sky130_fd_sc_hd__o211ai_4 _14494_ (.A1(_11037_),
    .A2(net1022),
    .B1(net1554),
    .C1(_07440_),
    .Y(_07441_));
 sky130_fd_sc_hd__o21ai_2 _14495_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7] ),
    .A2(net1026),
    .B1(_07441_),
    .Y(_07442_));
 sky130_fd_sc_hd__a22oi_2 _14496_ (.A1(\cs_registers_i.csr_mepc_o[6] ),
    .A2(_12452_),
    .B1(_12459_),
    .B2(\cs_registers_i.csr_depc_o[6] ),
    .Y(_07443_));
 sky130_fd_sc_hd__o2111ai_4 _14497_ (.A1(_11037_),
    .A2(net1037),
    .B1(net1554),
    .C1(_12753_),
    .D1(_07443_),
    .Y(_07444_));
 sky130_fd_sc_hd__o21ai_2 _14498_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6] ),
    .A2(_11043_),
    .B1(_07444_),
    .Y(_07445_));
 sky130_fd_sc_hd__a22oi_1 _14499_ (.A1(\cs_registers_i.csr_mepc_o[5] ),
    .A2(_12452_),
    .B1(_12459_),
    .B2(\cs_registers_i.csr_depc_o[5] ),
    .Y(_07446_));
 sky130_fd_sc_hd__nand3_1 _14500_ (.A(_11043_),
    .B(_12747_),
    .C(_07446_),
    .Y(_07447_));
 sky130_fd_sc_hd__a21o_1 _14501_ (.A1(net319),
    .A2(net176),
    .B1(_07447_),
    .X(_07448_));
 sky130_fd_sc_hd__o21ai_4 _14502_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5] ),
    .A2(net1554),
    .B1(_07448_),
    .Y(_07449_));
 sky130_fd_sc_hd__a22oi_1 _14503_ (.A1(\cs_registers_i.csr_mepc_o[4] ),
    .A2(_12452_),
    .B1(_12459_),
    .B2(\cs_registers_i.csr_depc_o[4] ),
    .Y(_07450_));
 sky130_fd_sc_hd__nand3_1 _14504_ (.A(_11043_),
    .B(_12742_),
    .C(_07450_),
    .Y(_07451_));
 sky130_fd_sc_hd__a21oi_2 _14505_ (.A1(net319),
    .A2(net175),
    .B1(_07451_),
    .Y(_07452_));
 sky130_fd_sc_hd__o21bai_4 _14506_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4] ),
    .A2(net1554),
    .B1_N(_07452_),
    .Y(_07453_));
 sky130_fd_sc_hd__a22oi_1 _14507_ (.A1(\cs_registers_i.csr_mepc_o[3] ),
    .A2(_12452_),
    .B1(_12459_),
    .B2(\cs_registers_i.csr_depc_o[3] ),
    .Y(_07454_));
 sky130_fd_sc_hd__nand4_1 _14508_ (.A(_11043_),
    .B(_12729_),
    .C(_07429_),
    .D(_07454_),
    .Y(_07455_));
 sky130_fd_sc_hd__a21o_1 _14509_ (.A1(net319),
    .A2(net1525),
    .B1(_07455_),
    .X(_07456_));
 sky130_fd_sc_hd__o21ai_2 _14510_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3] ),
    .A2(_11043_),
    .B1(_07456_),
    .Y(_07457_));
 sky130_fd_sc_hd__nand2_4 _14511_ (.A(_10994_),
    .B(_07331_),
    .Y(_07458_));
 sky130_fd_sc_hd__a22oi_2 _14512_ (.A1(\cs_registers_i.csr_mepc_o[2] ),
    .A2(_12452_),
    .B1(_12459_),
    .B2(\cs_registers_i.csr_depc_o[2] ),
    .Y(_07459_));
 sky130_fd_sc_hd__o2111ai_4 _14513_ (.A1(_11037_),
    .A2(net1464),
    .B1(net1554),
    .C1(_12712_),
    .D1(_07459_),
    .Y(_07460_));
 sky130_fd_sc_hd__o21ai_2 _14514_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2] ),
    .A2(_11043_),
    .B1(_07460_),
    .Y(_07461_));
 sky130_fd_sc_hd__or2_0 _14515_ (.A(_07458_),
    .B(_07461_),
    .X(_07462_));
 sky130_fd_sc_hd__nor2_1 _14516_ (.A(_07457_),
    .B(_07462_),
    .Y(_07463_));
 sky130_fd_sc_hd__nor4b_2 _14517_ (.A(_07445_),
    .B(_07449_),
    .C(_07453_),
    .D_N(_07463_),
    .Y(_07464_));
 sky130_fd_sc_hd__nor2_1 _14518_ (.A(net24),
    .B(_07423_),
    .Y(_07465_));
 sky130_fd_sc_hd__nand2_1 _14519_ (.A(\cs_registers_i.csr_mtvec_o[9] ),
    .B(_07430_),
    .Y(_07466_));
 sky130_fd_sc_hd__a22oi_1 _14520_ (.A1(\cs_registers_i.csr_mepc_o[9] ),
    .A2(_12455_),
    .B1(_07433_),
    .B2(\cs_registers_i.csr_depc_o[9] ),
    .Y(_07467_));
 sky130_fd_sc_hd__nand2_1 _14521_ (.A(_07466_),
    .B(_07467_),
    .Y(_07468_));
 sky130_fd_sc_hd__a211oi_2 _14522_ (.A1(net319),
    .A2(net1587),
    .B1(_07425_),
    .C1(_07468_),
    .Y(_07469_));
 sky130_fd_sc_hd__nand2_1 _14523_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ),
    .B(net292),
    .Y(_07470_));
 sky130_fd_sc_hd__o31ai_2 _14524_ (.A1(net292),
    .A2(_07465_),
    .A3(_07469_),
    .B1(_07470_),
    .Y(_07471_));
 sky130_fd_sc_hd__nor2_1 _14525_ (.A(net23),
    .B(_07423_),
    .Y(_07472_));
 sky130_fd_sc_hd__nand2_1 _14526_ (.A(\cs_registers_i.csr_depc_o[8] ),
    .B(_12459_),
    .Y(_07473_));
 sky130_fd_sc_hd__a22oi_1 _14527_ (.A1(\cs_registers_i.csr_mepc_o[8] ),
    .A2(_12452_),
    .B1(_07430_),
    .B2(\cs_registers_i.csr_mtvec_o[8] ),
    .Y(_07474_));
 sky130_fd_sc_hd__o2111a_2 _14528_ (.A1(_11037_),
    .A2(net1066),
    .B1(_07423_),
    .C1(_07473_),
    .D1(_07474_),
    .X(_07475_));
 sky130_fd_sc_hd__nand2_1 _14529_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ),
    .B(net292),
    .Y(_07476_));
 sky130_fd_sc_hd__o31ai_4 _14530_ (.A1(net292),
    .A2(_07472_),
    .A3(_07475_),
    .B1(_07476_),
    .Y(_07477_));
 sky130_fd_sc_hd__and4b_1 _14531_ (.A_N(_07442_),
    .B(_07464_),
    .C(_07471_),
    .D(_07477_),
    .X(_07478_));
 sky130_fd_sc_hd__and2_1 _14532_ (.A(_07439_),
    .B(_07478_),
    .X(_07479_));
 sky130_fd_sc_hd__nor2_1 _14533_ (.A(_07439_),
    .B(_07478_),
    .Y(_07480_));
 sky130_fd_sc_hd__nor2_1 _14534_ (.A(_07479_),
    .B(_07480_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[10] ));
 sky130_fd_sc_hd__nand2_1 _14535_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11] ),
    .B(net291),
    .Y(_07481_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1232 ();
 sky130_fd_sc_hd__nand2_4 _14537_ (.A(_11009_),
    .B(_07429_),
    .Y(_07483_));
 sky130_fd_sc_hd__o21ai_1 _14538_ (.A1(\cs_registers_i.csr_mtvec_o[11] ),
    .A2(_07483_),
    .B1(_07428_),
    .Y(_07484_));
 sky130_fd_sc_hd__a22oi_2 _14539_ (.A1(\cs_registers_i.csr_mepc_o[11] ),
    .A2(_12452_),
    .B1(_12459_),
    .B2(\cs_registers_i.csr_depc_o[11] ),
    .Y(_07485_));
 sky130_fd_sc_hd__o2111ai_4 _14540_ (.A1(_11037_),
    .A2(net1590),
    .B1(_07423_),
    .C1(_07484_),
    .D1(_07485_),
    .Y(_07486_));
 sky130_fd_sc_hd__o211ai_4 _14541_ (.A1(net2),
    .A2(_07423_),
    .B1(_07486_),
    .C1(net1554),
    .Y(_07487_));
 sky130_fd_sc_hd__nand2_2 _14542_ (.A(_07481_),
    .B(_07487_),
    .Y(_07488_));
 sky130_fd_sc_hd__xor2_1 _14543_ (.A(_07479_),
    .B(_07488_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[11] ));
 sky130_fd_sc_hd__nor2_1 _14544_ (.A(net3),
    .B(_07423_),
    .Y(_07489_));
 sky130_fd_sc_hd__nand2_1 _14545_ (.A(\cs_registers_i.csr_mtvec_o[12] ),
    .B(_07430_),
    .Y(_07490_));
 sky130_fd_sc_hd__a22oi_1 _14546_ (.A1(\cs_registers_i.csr_mepc_o[12] ),
    .A2(_12455_),
    .B1(_07433_),
    .B2(\cs_registers_i.csr_depc_o[12] ),
    .Y(_07491_));
 sky130_fd_sc_hd__nand2_1 _14547_ (.A(_07490_),
    .B(_07491_),
    .Y(_07492_));
 sky130_fd_sc_hd__a211oi_4 _14548_ (.A1(net1557),
    .A2(net319),
    .B1(_07425_),
    .C1(_07492_),
    .Y(_07493_));
 sky130_fd_sc_hd__nand2_1 _14549_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12] ),
    .B(net291),
    .Y(_07494_));
 sky130_fd_sc_hd__o31ai_4 _14550_ (.A1(net291),
    .A2(_07493_),
    .A3(_07489_),
    .B1(_07494_),
    .Y(_07495_));
 sky130_fd_sc_hd__and3_1 _14551_ (.A(_07479_),
    .B(_07488_),
    .C(_07495_),
    .X(_07496_));
 sky130_fd_sc_hd__a21oi_1 _14552_ (.A1(_07479_),
    .A2(_07488_),
    .B1(_07495_),
    .Y(_07497_));
 sky130_fd_sc_hd__nor2_1 _14553_ (.A(_07496_),
    .B(_07497_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[12] ));
 sky130_fd_sc_hd__a22o_1 _14554_ (.A1(\cs_registers_i.csr_depc_o[13] ),
    .A2(_12459_),
    .B1(_07430_),
    .B2(\cs_registers_i.csr_mtvec_o[13] ),
    .X(_07498_));
 sky130_fd_sc_hd__a21oi_1 _14555_ (.A1(\cs_registers_i.csr_mepc_o[13] ),
    .A2(_12452_),
    .B1(_07498_),
    .Y(_07499_));
 sky130_fd_sc_hd__nand2_1 _14556_ (.A(net319),
    .B(net1571),
    .Y(_07500_));
 sky130_fd_sc_hd__nor2_1 _14557_ (.A(net4),
    .B(_07423_),
    .Y(_07501_));
 sky130_fd_sc_hd__a311oi_4 _14558_ (.A1(_07423_),
    .A2(_07500_),
    .A3(_07499_),
    .B1(_07501_),
    .C1(net291),
    .Y(_07502_));
 sky130_fd_sc_hd__a21o_1 _14559_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13] ),
    .A2(net291),
    .B1(_07502_),
    .X(_07503_));
 sky130_fd_sc_hd__xor2_1 _14560_ (.A(_07496_),
    .B(_07503_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[13] ));
 sky130_fd_sc_hd__nand4_1 _14561_ (.A(_07479_),
    .B(_07488_),
    .C(_07495_),
    .D(_07503_),
    .Y(_07504_));
 sky130_fd_sc_hd__a22o_1 _14562_ (.A1(\cs_registers_i.csr_depc_o[14] ),
    .A2(_12459_),
    .B1(_07430_),
    .B2(\cs_registers_i.csr_mtvec_o[14] ),
    .X(_07505_));
 sky130_fd_sc_hd__a221oi_4 _14563_ (.A1(net1273),
    .A2(net319),
    .B1(_12452_),
    .B2(\cs_registers_i.csr_mepc_o[14] ),
    .C1(_07505_),
    .Y(_07506_));
 sky130_fd_sc_hd__nor2_1 _14564_ (.A(net5),
    .B(_07423_),
    .Y(_07507_));
 sky130_fd_sc_hd__a211o_1 _14565_ (.A1(_07506_),
    .A2(_07423_),
    .B1(_07507_),
    .C1(net291),
    .X(_07508_));
 sky130_fd_sc_hd__a21boi_4 _14566_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14] ),
    .A2(net291),
    .B1_N(_07508_),
    .Y(_07509_));
 sky130_fd_sc_hd__xor2_1 _14567_ (.A(_07504_),
    .B(_07509_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[14] ));
 sky130_fd_sc_hd__or2_1 _14568_ (.A(_07504_),
    .B(_07509_),
    .X(_07510_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1231 ();
 sky130_fd_sc_hd__a22o_1 _14570_ (.A1(\cs_registers_i.csr_depc_o[15] ),
    .A2(_12459_),
    .B1(_07430_),
    .B2(\cs_registers_i.csr_mtvec_o[15] ),
    .X(_07512_));
 sky130_fd_sc_hd__a21oi_1 _14571_ (.A1(\cs_registers_i.csr_mepc_o[15] ),
    .A2(_12452_),
    .B1(_07512_),
    .Y(_07513_));
 sky130_fd_sc_hd__nand2_8 _14572_ (.A(_08107_),
    .B(net721),
    .Y(_07514_));
 sky130_fd_sc_hd__nor2_1 _14573_ (.A(net6),
    .B(_07423_),
    .Y(_07515_));
 sky130_fd_sc_hd__a311oi_4 _14574_ (.A1(_07423_),
    .A2(_07513_),
    .A3(_07514_),
    .B1(_07515_),
    .C1(net290),
    .Y(_07516_));
 sky130_fd_sc_hd__a21oi_4 _14575_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ),
    .A2(net291),
    .B1(_07516_),
    .Y(_07517_));
 sky130_fd_sc_hd__xor2_1 _14576_ (.A(_07510_),
    .B(_07517_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[15] ));
 sky130_fd_sc_hd__nor2_1 _14577_ (.A(_07510_),
    .B(_07517_),
    .Y(_07518_));
 sky130_fd_sc_hd__o21ai_0 _14578_ (.A1(\cs_registers_i.csr_mtvec_o[16] ),
    .A2(_07483_),
    .B1(_07428_),
    .Y(_07519_));
 sky130_fd_sc_hd__a22oi_1 _14579_ (.A1(\cs_registers_i.csr_mepc_o[16] ),
    .A2(_12455_),
    .B1(_07433_),
    .B2(\cs_registers_i.csr_depc_o[16] ),
    .Y(_07520_));
 sky130_fd_sc_hd__nand2_1 _14580_ (.A(_07519_),
    .B(_07520_),
    .Y(_07521_));
 sky130_fd_sc_hd__a21oi_1 _14581_ (.A1(net7),
    .A2(_07425_),
    .B1(_07521_),
    .Y(_07522_));
 sky130_fd_sc_hd__nand2_2 _14582_ (.A(_08107_),
    .B(net1581),
    .Y(_07523_));
 sky130_fd_sc_hd__nand3_4 _14583_ (.A(_11043_),
    .B(_07523_),
    .C(_07522_),
    .Y(_07524_));
 sky130_fd_sc_hd__o21ai_2 _14584_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ),
    .A2(net1026),
    .B1(_07524_),
    .Y(_07525_));
 sky130_fd_sc_hd__xnor2_1 _14585_ (.A(_07518_),
    .B(_07525_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[16] ));
 sky130_fd_sc_hd__nand2_2 _14586_ (.A(_08107_),
    .B(net1560),
    .Y(_07526_));
 sky130_fd_sc_hd__a22o_1 _14587_ (.A1(\cs_registers_i.csr_mepc_o[17] ),
    .A2(_12452_),
    .B1(_07430_),
    .B2(\cs_registers_i.csr_mtvec_o[17] ),
    .X(_07527_));
 sky130_fd_sc_hd__a221oi_2 _14588_ (.A1(\cs_registers_i.csr_depc_o[17] ),
    .A2(_12459_),
    .B1(_07425_),
    .B2(net8),
    .C1(_07527_),
    .Y(_07528_));
 sky130_fd_sc_hd__nand3_4 _14589_ (.A(_11043_),
    .B(_07528_),
    .C(_07526_),
    .Y(_07529_));
 sky130_fd_sc_hd__o21ai_4 _14590_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17] ),
    .A2(net1554),
    .B1(_07529_),
    .Y(_07530_));
 sky130_fd_sc_hd__inv_1 _14591_ (.A(_07530_),
    .Y(_07531_));
 sky130_fd_sc_hd__inv_1 _14592_ (.A(_07525_),
    .Y(_07532_));
 sky130_fd_sc_hd__nand2_1 _14593_ (.A(_07518_),
    .B(_07532_),
    .Y(_07533_));
 sky130_fd_sc_hd__xnor2_1 _14594_ (.A(_07531_),
    .B(_07533_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[17] ));
 sky130_fd_sc_hd__nor2_1 _14595_ (.A(net9),
    .B(_07423_),
    .Y(_07534_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1230 ();
 sky130_fd_sc_hd__nand2_1 _14597_ (.A(\cs_registers_i.csr_mtvec_o[18] ),
    .B(_07430_),
    .Y(_07536_));
 sky130_fd_sc_hd__a22oi_1 _14598_ (.A1(\cs_registers_i.csr_mepc_o[18] ),
    .A2(_12455_),
    .B1(_07433_),
    .B2(\cs_registers_i.csr_depc_o[18] ),
    .Y(_07537_));
 sky130_fd_sc_hd__nand2_1 _14599_ (.A(_07536_),
    .B(_07537_),
    .Y(_07538_));
 sky130_fd_sc_hd__a211oi_4 _14600_ (.A1(net319),
    .A2(net1241),
    .B1(_07425_),
    .C1(_07538_),
    .Y(_07539_));
 sky130_fd_sc_hd__nor3_4 _14601_ (.A(_07539_),
    .B(_07534_),
    .C(net290),
    .Y(_07540_));
 sky130_fd_sc_hd__a21o_1 _14602_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18] ),
    .A2(net292),
    .B1(_07540_),
    .X(_07541_));
 sky130_fd_sc_hd__nor4_1 _14603_ (.A(_07510_),
    .B(_07517_),
    .C(_07525_),
    .D(_07530_),
    .Y(_07542_));
 sky130_fd_sc_hd__xor2_1 _14604_ (.A(_07541_),
    .B(_07542_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[18] ));
 sky130_fd_sc_hd__nand2_1 _14605_ (.A(_07541_),
    .B(_07542_),
    .Y(_07543_));
 sky130_fd_sc_hd__nand2_1 _14606_ (.A(net319),
    .B(net1260),
    .Y(_07544_));
 sky130_fd_sc_hd__a22o_1 _14607_ (.A1(\cs_registers_i.csr_depc_o[19] ),
    .A2(_12459_),
    .B1(_07430_),
    .B2(\cs_registers_i.csr_mtvec_o[19] ),
    .X(_07545_));
 sky130_fd_sc_hd__a21oi_1 _14608_ (.A1(\cs_registers_i.csr_mepc_o[19] ),
    .A2(_12452_),
    .B1(_07545_),
    .Y(_07546_));
 sky130_fd_sc_hd__nand2_1 _14609_ (.A(net10),
    .B(_07425_),
    .Y(_07547_));
 sky130_fd_sc_hd__nand4_4 _14610_ (.A(_11043_),
    .B(_07544_),
    .C(_07546_),
    .D(_07547_),
    .Y(_07548_));
 sky130_fd_sc_hd__o21ai_2 _14611_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19] ),
    .A2(net1026),
    .B1(_07548_),
    .Y(_07549_));
 sky130_fd_sc_hd__xor2_1 _14612_ (.A(_07543_),
    .B(_07549_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[19] ));
 sky130_fd_sc_hd__o21ai_0 _14613_ (.A1(\cs_registers_i.csr_mtvec_o[20] ),
    .A2(_07483_),
    .B1(_07428_),
    .Y(_07550_));
 sky130_fd_sc_hd__a22oi_1 _14614_ (.A1(\cs_registers_i.csr_mepc_o[20] ),
    .A2(_12455_),
    .B1(_07433_),
    .B2(\cs_registers_i.csr_depc_o[20] ),
    .Y(_07551_));
 sky130_fd_sc_hd__nand2_1 _14615_ (.A(_07550_),
    .B(_07551_),
    .Y(_07552_));
 sky130_fd_sc_hd__a21oi_1 _14616_ (.A1(net11),
    .A2(_07425_),
    .B1(_07552_),
    .Y(_07553_));
 sky130_fd_sc_hd__nand2_1 _14617_ (.A(net319),
    .B(net1007),
    .Y(_07554_));
 sky130_fd_sc_hd__nand3_4 _14618_ (.A(_11043_),
    .B(_07553_),
    .C(_07554_),
    .Y(_07555_));
 sky130_fd_sc_hd__o21ai_2 _14619_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20] ),
    .A2(net1554),
    .B1(_07555_),
    .Y(_07556_));
 sky130_fd_sc_hd__nor2_1 _14620_ (.A(_07543_),
    .B(_07549_),
    .Y(_07557_));
 sky130_fd_sc_hd__xnor2_1 _14621_ (.A(_07556_),
    .B(_07557_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[20] ));
 sky130_fd_sc_hd__nand2_1 _14622_ (.A(net319),
    .B(net1259),
    .Y(_07558_));
 sky130_fd_sc_hd__a22o_1 _14623_ (.A1(\cs_registers_i.csr_mepc_o[21] ),
    .A2(_12452_),
    .B1(_07430_),
    .B2(\cs_registers_i.csr_mtvec_o[21] ),
    .X(_07559_));
 sky130_fd_sc_hd__a221oi_2 _14624_ (.A1(\cs_registers_i.csr_depc_o[21] ),
    .A2(_12459_),
    .B1(_07425_),
    .B2(net12),
    .C1(_07559_),
    .Y(_07560_));
 sky130_fd_sc_hd__nand3_4 _14625_ (.A(net1554),
    .B(_07558_),
    .C(_07560_),
    .Y(_07561_));
 sky130_fd_sc_hd__o21ai_2 _14626_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ),
    .A2(net1026),
    .B1(_07561_),
    .Y(_07562_));
 sky130_fd_sc_hd__nor3_1 _14627_ (.A(_07543_),
    .B(_07549_),
    .C(_07556_),
    .Y(_07563_));
 sky130_fd_sc_hd__xnor2_1 _14628_ (.A(_07562_),
    .B(_07563_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[21] ));
 sky130_fd_sc_hd__nand2_2 _14629_ (.A(net319),
    .B(net1547),
    .Y(_07564_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1229 ();
 sky130_fd_sc_hd__a22o_1 _14631_ (.A1(\cs_registers_i.csr_mepc_o[22] ),
    .A2(_12452_),
    .B1(_07430_),
    .B2(\cs_registers_i.csr_mtvec_o[22] ),
    .X(_07566_));
 sky130_fd_sc_hd__a221oi_2 _14632_ (.A1(\cs_registers_i.csr_depc_o[22] ),
    .A2(_12459_),
    .B1(_07425_),
    .B2(net13),
    .C1(_07566_),
    .Y(_07567_));
 sky130_fd_sc_hd__nand3_4 _14633_ (.A(net1554),
    .B(_07564_),
    .C(_07567_),
    .Y(_07568_));
 sky130_fd_sc_hd__o21ai_2 _14634_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22] ),
    .A2(net1026),
    .B1(_07568_),
    .Y(_07569_));
 sky130_fd_sc_hd__nand4_1 _14635_ (.A(_07518_),
    .B(_07532_),
    .C(_07531_),
    .D(_07541_),
    .Y(_07570_));
 sky130_fd_sc_hd__nor4_2 _14636_ (.A(_07570_),
    .B(_07549_),
    .C(_07556_),
    .D(_07562_),
    .Y(_07571_));
 sky130_fd_sc_hd__xnor2_1 _14637_ (.A(_07569_),
    .B(_07571_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[22] ));
 sky130_fd_sc_hd__nand2_4 _14638_ (.A(_08107_),
    .B(net164),
    .Y(_07572_));
 sky130_fd_sc_hd__a22o_1 _14639_ (.A1(\cs_registers_i.csr_mepc_o[23] ),
    .A2(_12452_),
    .B1(_07430_),
    .B2(\cs_registers_i.csr_mtvec_o[23] ),
    .X(_07573_));
 sky130_fd_sc_hd__a221oi_4 _14640_ (.A1(\cs_registers_i.csr_depc_o[23] ),
    .A2(_12459_),
    .B1(_07425_),
    .B2(net14),
    .C1(_07573_),
    .Y(_07574_));
 sky130_fd_sc_hd__nand3_4 _14641_ (.A(net1554),
    .B(_07572_),
    .C(_07574_),
    .Y(_07575_));
 sky130_fd_sc_hd__o21ai_2 _14642_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23] ),
    .A2(net1026),
    .B1(_07575_),
    .Y(_07576_));
 sky130_fd_sc_hd__and2b_1 _14643_ (.A_N(_07569_),
    .B(_07571_),
    .X(_07577_));
 sky130_fd_sc_hd__xnor2_1 _14644_ (.A(_07576_),
    .B(_07577_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[23] ));
 sky130_fd_sc_hd__nand2_4 _14645_ (.A(net774),
    .B(net319),
    .Y(_07578_));
 sky130_fd_sc_hd__a22o_1 _14646_ (.A1(\cs_registers_i.csr_mepc_o[24] ),
    .A2(_12452_),
    .B1(_07430_),
    .B2(\cs_registers_i.csr_mtvec_o[24] ),
    .X(_07579_));
 sky130_fd_sc_hd__a221oi_2 _14647_ (.A1(\cs_registers_i.csr_depc_o[24] ),
    .A2(_12459_),
    .B1(_07425_),
    .B2(net15),
    .C1(_07579_),
    .Y(_07580_));
 sky130_fd_sc_hd__nand3_4 _14648_ (.A(_11043_),
    .B(_07578_),
    .C(_07580_),
    .Y(_07581_));
 sky130_fd_sc_hd__o21ai_4 _14649_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24] ),
    .A2(net1026),
    .B1(_07581_),
    .Y(_07582_));
 sky130_fd_sc_hd__nand2b_1 _14650_ (.A_N(_07576_),
    .B(_07577_),
    .Y(_07583_));
 sky130_fd_sc_hd__xor2_1 _14651_ (.A(_07582_),
    .B(_07583_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[24] ));
 sky130_fd_sc_hd__o21ai_0 _14652_ (.A1(\cs_registers_i.csr_mtvec_o[25] ),
    .A2(_07483_),
    .B1(_07428_),
    .Y(_07584_));
 sky130_fd_sc_hd__a22oi_1 _14653_ (.A1(\cs_registers_i.csr_mepc_o[25] ),
    .A2(_12455_),
    .B1(_07433_),
    .B2(\cs_registers_i.csr_depc_o[25] ),
    .Y(_07585_));
 sky130_fd_sc_hd__nand2_1 _14654_ (.A(_07584_),
    .B(_07585_),
    .Y(_07586_));
 sky130_fd_sc_hd__a211oi_1 _14655_ (.A1(net16),
    .A2(_07425_),
    .B1(_07586_),
    .C1(net290),
    .Y(_07587_));
 sky130_fd_sc_hd__o21ai_4 _14656_ (.A1(_11037_),
    .A2(net684),
    .B1(_07587_),
    .Y(_07588_));
 sky130_fd_sc_hd__o21a_1 _14657_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25] ),
    .A2(net1026),
    .B1(_07588_),
    .X(_07589_));
 sky130_fd_sc_hd__nor2_1 _14658_ (.A(_07582_),
    .B(_07583_),
    .Y(_07590_));
 sky130_fd_sc_hd__xor2_1 _14659_ (.A(_07589_),
    .B(_07590_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[25] ));
 sky130_fd_sc_hd__a22o_1 _14660_ (.A1(\cs_registers_i.csr_mepc_o[26] ),
    .A2(_12452_),
    .B1(_07430_),
    .B2(\cs_registers_i.csr_mtvec_o[26] ),
    .X(_07591_));
 sky130_fd_sc_hd__a221oi_2 _14661_ (.A1(\cs_registers_i.csr_depc_o[26] ),
    .A2(_12459_),
    .B1(_07425_),
    .B2(net17),
    .C1(_07591_),
    .Y(_07592_));
 sky130_fd_sc_hd__o211ai_4 _14662_ (.A1(_11037_),
    .A2(_10535_),
    .B1(net1554),
    .C1(_07592_),
    .Y(_07593_));
 sky130_fd_sc_hd__o21ai_4 _14663_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26] ),
    .A2(net1026),
    .B1(_07593_),
    .Y(_07594_));
 sky130_fd_sc_hd__nand2_1 _14664_ (.A(_07589_),
    .B(_07590_),
    .Y(_07595_));
 sky130_fd_sc_hd__xor2_1 _14665_ (.A(_07594_),
    .B(_07595_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[26] ));
 sky130_fd_sc_hd__o21ai_0 _14666_ (.A1(\cs_registers_i.csr_mtvec_o[27] ),
    .A2(_07483_),
    .B1(_07428_),
    .Y(_07596_));
 sky130_fd_sc_hd__a22oi_1 _14667_ (.A1(\cs_registers_i.csr_mepc_o[27] ),
    .A2(_12455_),
    .B1(_07433_),
    .B2(\cs_registers_i.csr_depc_o[27] ),
    .Y(_07597_));
 sky130_fd_sc_hd__nand2_1 _14668_ (.A(_07596_),
    .B(_07597_),
    .Y(_07598_));
 sky130_fd_sc_hd__a21oi_1 _14669_ (.A1(net18),
    .A2(_07425_),
    .B1(_07598_),
    .Y(_07599_));
 sky130_fd_sc_hd__nand2_2 _14670_ (.A(_08107_),
    .B(net168),
    .Y(_07600_));
 sky130_fd_sc_hd__nand3_4 _14671_ (.A(_11043_),
    .B(_07600_),
    .C(_07599_),
    .Y(_07601_));
 sky130_fd_sc_hd__o21ai_4 _14672_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27] ),
    .A2(net1026),
    .B1(_07601_),
    .Y(_07602_));
 sky130_fd_sc_hd__nor2_1 _14673_ (.A(_07594_),
    .B(_07595_),
    .Y(_07603_));
 sky130_fd_sc_hd__xnor2_1 _14674_ (.A(_07602_),
    .B(_07603_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[27] ));
 sky130_fd_sc_hd__o21ai_0 _14675_ (.A1(\cs_registers_i.csr_mtvec_o[28] ),
    .A2(_07483_),
    .B1(_07428_),
    .Y(_07604_));
 sky130_fd_sc_hd__a22oi_1 _14676_ (.A1(\cs_registers_i.csr_mepc_o[28] ),
    .A2(_12455_),
    .B1(_07433_),
    .B2(\cs_registers_i.csr_depc_o[28] ),
    .Y(_07605_));
 sky130_fd_sc_hd__nand2_1 _14677_ (.A(_07604_),
    .B(_07605_),
    .Y(_07606_));
 sky130_fd_sc_hd__a21oi_1 _14678_ (.A1(net19),
    .A2(_07425_),
    .B1(_07606_),
    .Y(_07607_));
 sky130_fd_sc_hd__nand2_2 _14679_ (.A(_08107_),
    .B(net169),
    .Y(_07608_));
 sky130_fd_sc_hd__nand3_4 _14680_ (.A(_11043_),
    .B(_07608_),
    .C(_07607_),
    .Y(_07609_));
 sky130_fd_sc_hd__o21ai_4 _14681_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28] ),
    .A2(net1026),
    .B1(_07609_),
    .Y(_07610_));
 sky130_fd_sc_hd__or3_1 _14682_ (.A(_07594_),
    .B(_07595_),
    .C(_07602_),
    .X(_07611_));
 sky130_fd_sc_hd__xor2_1 _14683_ (.A(_07610_),
    .B(_07611_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[28] ));
 sky130_fd_sc_hd__a22o_1 _14684_ (.A1(\cs_registers_i.csr_mepc_o[29] ),
    .A2(_12452_),
    .B1(_07430_),
    .B2(\cs_registers_i.csr_mtvec_o[29] ),
    .X(_07612_));
 sky130_fd_sc_hd__a221oi_2 _14685_ (.A1(\cs_registers_i.csr_depc_o[29] ),
    .A2(_12459_),
    .B1(_07425_),
    .B2(net20),
    .C1(_07612_),
    .Y(_07613_));
 sky130_fd_sc_hd__o211ai_4 _14686_ (.A1(_11037_),
    .A2(_10665_),
    .B1(_11043_),
    .C1(_07613_),
    .Y(_07614_));
 sky130_fd_sc_hd__o21a_1 _14687_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29] ),
    .A2(net1026),
    .B1(_07614_),
    .X(_07615_));
 sky130_fd_sc_hd__nor2_1 _14688_ (.A(_07610_),
    .B(_07611_),
    .Y(_07616_));
 sky130_fd_sc_hd__xor2_1 _14689_ (.A(_07615_),
    .B(_07616_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[29] ));
 sky130_fd_sc_hd__xor2_1 _14690_ (.A(_07458_),
    .B(_07461_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[2] ));
 sky130_fd_sc_hd__a22o_1 _14691_ (.A1(\cs_registers_i.csr_mepc_o[30] ),
    .A2(_12452_),
    .B1(_07430_),
    .B2(\cs_registers_i.csr_mtvec_o[30] ),
    .X(_07617_));
 sky130_fd_sc_hd__a221oi_2 _14692_ (.A1(\cs_registers_i.csr_depc_o[30] ),
    .A2(_12459_),
    .B1(_07425_),
    .B2(net21),
    .C1(_07617_),
    .Y(_07618_));
 sky130_fd_sc_hd__o211ai_4 _14693_ (.A1(_11037_),
    .A2(_10809_),
    .B1(net1554),
    .C1(_07618_),
    .Y(_07619_));
 sky130_fd_sc_hd__o21ai_4 _14694_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30] ),
    .A2(net1026),
    .B1(_07619_),
    .Y(_07620_));
 sky130_fd_sc_hd__nand2_1 _14695_ (.A(_07615_),
    .B(_07616_),
    .Y(_07621_));
 sky130_fd_sc_hd__xor2_1 _14696_ (.A(_07620_),
    .B(_07621_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[30] ));
 sky130_fd_sc_hd__a22o_1 _14697_ (.A1(\cs_registers_i.csr_mepc_o[31] ),
    .A2(_12452_),
    .B1(_07430_),
    .B2(\cs_registers_i.csr_mtvec_o[31] ),
    .X(_07622_));
 sky130_fd_sc_hd__a221oi_2 _14698_ (.A1(\cs_registers_i.csr_depc_o[31] ),
    .A2(_12459_),
    .B1(_07425_),
    .B2(net22),
    .C1(_07622_),
    .Y(_07623_));
 sky130_fd_sc_hd__o211ai_4 _14699_ (.A1(_11037_),
    .A2(_13466_),
    .B1(net1554),
    .C1(_07623_),
    .Y(_07624_));
 sky130_fd_sc_hd__o21ai_2 _14700_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31] ),
    .A2(net1026),
    .B1(_07624_),
    .Y(_07625_));
 sky130_fd_sc_hd__nor2_1 _14701_ (.A(_07620_),
    .B(_07621_),
    .Y(_07626_));
 sky130_fd_sc_hd__xnor2_1 _14702_ (.A(_07625_),
    .B(_07626_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[31] ));
 sky130_fd_sc_hd__xor2_1 _14703_ (.A(_07457_),
    .B(_07462_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[3] ));
 sky130_fd_sc_hd__xnor2_1 _14704_ (.A(_07453_),
    .B(_07463_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[4] ));
 sky130_fd_sc_hd__nand2b_1 _14705_ (.A_N(_07453_),
    .B(_07463_),
    .Y(_07627_));
 sky130_fd_sc_hd__xor2_1 _14706_ (.A(_07449_),
    .B(_07627_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[5] ));
 sky130_fd_sc_hd__nor2_1 _14707_ (.A(_07449_),
    .B(_07627_),
    .Y(_07628_));
 sky130_fd_sc_hd__xnor2_1 _14708_ (.A(_07445_),
    .B(_07628_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[6] ));
 sky130_fd_sc_hd__xnor2_1 _14709_ (.A(_07442_),
    .B(_07464_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[7] ));
 sky130_fd_sc_hd__nand2b_1 _14710_ (.A_N(_07442_),
    .B(_07464_),
    .Y(_07629_));
 sky130_fd_sc_hd__xnor2_1 _14711_ (.A(_07477_),
    .B(_07629_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[8] ));
 sky130_fd_sc_hd__nand2b_1 _14712_ (.A_N(_07629_),
    .B(_07477_),
    .Y(_07630_));
 sky130_fd_sc_hd__xnor2_1 _14713_ (.A(_07471_),
    .B(_07630_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[9] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1228 ();
 sky130_fd_sc_hd__nand2_8 _14715_ (.A(net293),
    .B(_07458_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ));
 sky130_fd_sc_hd__a21oi_1 _14716_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ),
    .B1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ),
    .Y(_07632_));
 sky130_fd_sc_hd__a211oi_1 _14717_ (.A1(net96),
    .A2(net107),
    .B1(net94),
    .C1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_07633_));
 sky130_fd_sc_hd__a21oi_2 _14718_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .A2(_07632_),
    .B1(_07633_),
    .Y(_07634_));
 sky130_fd_sc_hd__nor2_2 _14719_ (.A(\cs_registers_i.pc_if_i[1] ),
    .B(_07634_),
    .Y(_07635_));
 sky130_fd_sc_hd__nor3_4 _14720_ (.A(_11164_),
    .B(_11201_),
    .C(_07635_),
    .Y(_07636_));
 sky130_fd_sc_hd__nand2b_1 _14721_ (.A_N(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .B(_07636_),
    .Y(_07637_));
 sky130_fd_sc_hd__nand2b_4 _14722_ (.A_N(_07636_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_07638_));
 sky130_fd_sc_hd__nand3_4 _14723_ (.A(_11139_),
    .B(_07637_),
    .C(_07638_),
    .Y(_07639_));
 sky130_fd_sc_hd__nand2_4 _14724_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .B(_07636_),
    .Y(_07640_));
 sky130_fd_sc_hd__nand2_8 _14725_ (.A(_07640_),
    .B(_07639_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ));
 sky130_fd_sc_hd__o21ai_4 _14726_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .A2(_07638_),
    .B1(_07640_),
    .Y(_07641_));
 sky130_fd_sc_hd__a22o_4 _14727_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .A2(net1292),
    .B1(_07641_),
    .B2(_11139_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ));
 sky130_fd_sc_hd__o21ai_0 _14728_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .A2(_07410_),
    .B1(_07323_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_d[0] ));
 sky130_fd_sc_hd__nand2_1 _14729_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2] ),
    .Y(_07642_));
 sky130_fd_sc_hd__o21ai_0 _14730_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .A2(_07410_),
    .B1(_07642_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_d[1] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1227 ();
 sky130_fd_sc_hd__nor2_1 _14732_ (.A(_11037_),
    .B(_13394_),
    .Y(_07644_));
 sky130_fd_sc_hd__a221oi_4 _14733_ (.A1(\cs_registers_i.csr_mepc_o[1] ),
    .A2(_12455_),
    .B1(_07433_),
    .B2(\cs_registers_i.csr_depc_o[1] ),
    .C1(_07644_),
    .Y(_07645_));
 sky130_fd_sc_hd__nor3_1 _14734_ (.A(net1026),
    .B(_11138_),
    .C(_07635_),
    .Y(_07646_));
 sky130_fd_sc_hd__a21oi_1 _14735_ (.A1(net1026),
    .A2(_07645_),
    .B1(_07646_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[1] ));
 sky130_fd_sc_hd__inv_1 _14736_ (.A(\cs_registers_i.pc_if_i[9] ),
    .Y(_07647_));
 sky130_fd_sc_hd__inv_1 _14737_ (.A(\cs_registers_i.pc_if_i[6] ),
    .Y(_07648_));
 sky130_fd_sc_hd__nor2b_2 _14738_ (.A(_07635_),
    .B_N(\cs_registers_i.pc_if_i[2] ),
    .Y(_07649_));
 sky130_fd_sc_hd__nand4_1 _14739_ (.A(\cs_registers_i.pc_if_i[3] ),
    .B(\cs_registers_i.pc_if_i[4] ),
    .C(\cs_registers_i.pc_if_i[5] ),
    .D(_07649_),
    .Y(_07650_));
 sky130_fd_sc_hd__nor2_1 _14740_ (.A(_07648_),
    .B(_07650_),
    .Y(_07651_));
 sky130_fd_sc_hd__nand3_1 _14741_ (.A(\cs_registers_i.pc_if_i[7] ),
    .B(\cs_registers_i.pc_if_i[8] ),
    .C(_07651_),
    .Y(_07652_));
 sky130_fd_sc_hd__nor2_1 _14742_ (.A(_07647_),
    .B(_07652_),
    .Y(_07653_));
 sky130_fd_sc_hd__nand2_1 _14743_ (.A(\cs_registers_i.pc_if_i[10] ),
    .B(_07653_),
    .Y(_07654_));
 sky130_fd_sc_hd__xor2_1 _14744_ (.A(\cs_registers_i.pc_if_i[11] ),
    .B(_07654_),
    .X(_07655_));
 sky130_fd_sc_hd__o21ai_0 _14745_ (.A1(net1026),
    .A2(_07655_),
    .B1(_07487_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[11] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1226 ();
 sky130_fd_sc_hd__and3_1 _14747_ (.A(\cs_registers_i.pc_if_i[10] ),
    .B(\cs_registers_i.pc_if_i[11] ),
    .C(_07653_),
    .X(_07657_));
 sky130_fd_sc_hd__xor2_1 _14748_ (.A(\cs_registers_i.pc_if_i[12] ),
    .B(_07657_),
    .X(_07658_));
 sky130_fd_sc_hd__nand2_1 _14749_ (.A(net291),
    .B(_07658_),
    .Y(_07659_));
 sky130_fd_sc_hd__o31ai_1 _14750_ (.A1(net291),
    .A2(_07489_),
    .A3(_07493_),
    .B1(_07659_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[12] ));
 sky130_fd_sc_hd__nand2_1 _14751_ (.A(\cs_registers_i.pc_if_i[12] ),
    .B(_07657_),
    .Y(_07660_));
 sky130_fd_sc_hd__xnor2_1 _14752_ (.A(\cs_registers_i.pc_if_i[13] ),
    .B(_07660_),
    .Y(_07661_));
 sky130_fd_sc_hd__a21o_1 _14753_ (.A1(net291),
    .A2(_07661_),
    .B1(_07502_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[13] ));
 sky130_fd_sc_hd__inv_1 _14754_ (.A(\cs_registers_i.pc_if_i[14] ),
    .Y(_07662_));
 sky130_fd_sc_hd__nand3_1 _14755_ (.A(\cs_registers_i.pc_if_i[12] ),
    .B(\cs_registers_i.pc_if_i[13] ),
    .C(_07657_),
    .Y(_07663_));
 sky130_fd_sc_hd__xnor2_1 _14756_ (.A(_07662_),
    .B(_07663_),
    .Y(_07664_));
 sky130_fd_sc_hd__o21ai_0 _14757_ (.A1(net1026),
    .A2(_07664_),
    .B1(_07508_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[14] ));
 sky130_fd_sc_hd__nor2_2 _14758_ (.A(_07662_),
    .B(_07663_),
    .Y(_07665_));
 sky130_fd_sc_hd__xor2_1 _14759_ (.A(\cs_registers_i.pc_if_i[15] ),
    .B(_07665_),
    .X(_07666_));
 sky130_fd_sc_hd__a21o_1 _14760_ (.A1(net291),
    .A2(_07666_),
    .B1(_07516_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[15] ));
 sky130_fd_sc_hd__a21oi_1 _14761_ (.A1(\cs_registers_i.pc_if_i[15] ),
    .A2(_07665_),
    .B1(\cs_registers_i.pc_if_i[16] ),
    .Y(_07667_));
 sky130_fd_sc_hd__nand3_2 _14762_ (.A(\cs_registers_i.pc_if_i[15] ),
    .B(\cs_registers_i.pc_if_i[16] ),
    .C(_07665_),
    .Y(_07668_));
 sky130_fd_sc_hd__nor2b_1 _14763_ (.A(_07667_),
    .B_N(_07668_),
    .Y(_07669_));
 sky130_fd_sc_hd__o21a_1 _14764_ (.A1(net1026),
    .A2(_07669_),
    .B1(_07524_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[16] ));
 sky130_fd_sc_hd__inv_1 _14765_ (.A(\cs_registers_i.pc_if_i[17] ),
    .Y(_07670_));
 sky130_fd_sc_hd__xnor2_1 _14766_ (.A(_07670_),
    .B(_07668_),
    .Y(_07671_));
 sky130_fd_sc_hd__a21boi_0 _14767_ (.A1(net290),
    .A2(_07671_),
    .B1_N(_07529_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[17] ));
 sky130_fd_sc_hd__nor2_1 _14768_ (.A(_07670_),
    .B(_07668_),
    .Y(_07672_));
 sky130_fd_sc_hd__xor2_1 _14769_ (.A(\cs_registers_i.pc_if_i[18] ),
    .B(_07672_),
    .X(_07673_));
 sky130_fd_sc_hd__a21o_1 _14770_ (.A1(net290),
    .A2(_07673_),
    .B1(_07540_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[18] ));
 sky130_fd_sc_hd__a21o_1 _14771_ (.A1(\cs_registers_i.pc_if_i[18] ),
    .A2(_07672_),
    .B1(\cs_registers_i.pc_if_i[19] ),
    .X(_07674_));
 sky130_fd_sc_hd__nand3_2 _14772_ (.A(\cs_registers_i.pc_if_i[18] ),
    .B(\cs_registers_i.pc_if_i[19] ),
    .C(_07672_),
    .Y(_07675_));
 sky130_fd_sc_hd__nand2_1 _14773_ (.A(_07674_),
    .B(_07675_),
    .Y(_07676_));
 sky130_fd_sc_hd__a21boi_0 _14774_ (.A1(net290),
    .A2(_07676_),
    .B1_N(_07548_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[19] ));
 sky130_fd_sc_hd__inv_1 _14775_ (.A(\cs_registers_i.pc_if_i[20] ),
    .Y(_07677_));
 sky130_fd_sc_hd__xnor2_1 _14776_ (.A(_07677_),
    .B(_07675_),
    .Y(_07678_));
 sky130_fd_sc_hd__a21boi_0 _14777_ (.A1(net290),
    .A2(_07678_),
    .B1_N(_07555_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[20] ));
 sky130_fd_sc_hd__nor3_1 _14778_ (.A(\cs_registers_i.pc_if_i[1] ),
    .B(\cs_registers_i.pc_if_i[2] ),
    .C(_07634_),
    .Y(_07679_));
 sky130_fd_sc_hd__nor2_1 _14779_ (.A(_07649_),
    .B(_07679_),
    .Y(_07680_));
 sky130_fd_sc_hd__o21a_1 _14780_ (.A1(net1026),
    .A2(_07680_),
    .B1(_07460_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[2] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1225 ();
 sky130_fd_sc_hd__nor2_1 _14782_ (.A(_07677_),
    .B(_07675_),
    .Y(_07682_));
 sky130_fd_sc_hd__xnor2_1 _14783_ (.A(\cs_registers_i.pc_if_i[21] ),
    .B(_07682_),
    .Y(_07683_));
 sky130_fd_sc_hd__a21boi_0 _14784_ (.A1(net290),
    .A2(_07683_),
    .B1_N(_07561_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[21] ));
 sky130_fd_sc_hd__nand2_1 _14785_ (.A(\cs_registers_i.pc_if_i[21] ),
    .B(_07682_),
    .Y(_07684_));
 sky130_fd_sc_hd__xor2_1 _14786_ (.A(\cs_registers_i.pc_if_i[22] ),
    .B(_07684_),
    .X(_07685_));
 sky130_fd_sc_hd__a21boi_0 _14787_ (.A1(net290),
    .A2(_07685_),
    .B1_N(_07568_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[22] ));
 sky130_fd_sc_hd__a31oi_1 _14788_ (.A1(\cs_registers_i.pc_if_i[21] ),
    .A2(\cs_registers_i.pc_if_i[22] ),
    .A3(_07682_),
    .B1(\cs_registers_i.pc_if_i[23] ),
    .Y(_07686_));
 sky130_fd_sc_hd__and4_1 _14789_ (.A(\cs_registers_i.pc_if_i[21] ),
    .B(\cs_registers_i.pc_if_i[22] ),
    .C(\cs_registers_i.pc_if_i[23] ),
    .D(_07682_),
    .X(_07687_));
 sky130_fd_sc_hd__o21ai_0 _14790_ (.A1(_07686_),
    .A2(_07687_),
    .B1(net290),
    .Y(_07688_));
 sky130_fd_sc_hd__and2_0 _14791_ (.A(_07575_),
    .B(_07688_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[23] ));
 sky130_fd_sc_hd__xnor2_1 _14792_ (.A(\cs_registers_i.pc_if_i[24] ),
    .B(_07687_),
    .Y(_07689_));
 sky130_fd_sc_hd__a21boi_0 _14793_ (.A1(net290),
    .A2(_07689_),
    .B1_N(_07581_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[24] ));
 sky130_fd_sc_hd__nand2_1 _14794_ (.A(\cs_registers_i.pc_if_i[24] ),
    .B(_07687_),
    .Y(_07690_));
 sky130_fd_sc_hd__xor2_1 _14795_ (.A(\cs_registers_i.pc_if_i[25] ),
    .B(_07690_),
    .X(_07691_));
 sky130_fd_sc_hd__a21boi_0 _14796_ (.A1(net290),
    .A2(_07691_),
    .B1_N(_07588_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[25] ));
 sky130_fd_sc_hd__a31oi_1 _14797_ (.A1(\cs_registers_i.pc_if_i[24] ),
    .A2(\cs_registers_i.pc_if_i[25] ),
    .A3(_07687_),
    .B1(\cs_registers_i.pc_if_i[26] ),
    .Y(_07692_));
 sky130_fd_sc_hd__and4_1 _14798_ (.A(\cs_registers_i.pc_if_i[24] ),
    .B(\cs_registers_i.pc_if_i[25] ),
    .C(\cs_registers_i.pc_if_i[26] ),
    .D(_07687_),
    .X(_07693_));
 sky130_fd_sc_hd__o21ai_0 _14799_ (.A1(_07692_),
    .A2(_07693_),
    .B1(net290),
    .Y(_07694_));
 sky130_fd_sc_hd__and2_0 _14800_ (.A(_07593_),
    .B(_07694_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[26] ));
 sky130_fd_sc_hd__xnor2_1 _14801_ (.A(\cs_registers_i.pc_if_i[27] ),
    .B(_07693_),
    .Y(_07695_));
 sky130_fd_sc_hd__a21boi_0 _14802_ (.A1(net290),
    .A2(_07695_),
    .B1_N(_07601_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[27] ));
 sky130_fd_sc_hd__a21oi_1 _14803_ (.A1(\cs_registers_i.pc_if_i[27] ),
    .A2(_07693_),
    .B1(\cs_registers_i.pc_if_i[28] ),
    .Y(_07696_));
 sky130_fd_sc_hd__and3_1 _14804_ (.A(\cs_registers_i.pc_if_i[27] ),
    .B(\cs_registers_i.pc_if_i[28] ),
    .C(_07693_),
    .X(_07697_));
 sky130_fd_sc_hd__o21ai_0 _14805_ (.A1(_07696_),
    .A2(_07697_),
    .B1(net290),
    .Y(_07698_));
 sky130_fd_sc_hd__and2_0 _14806_ (.A(_07609_),
    .B(_07698_),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[28] ));
 sky130_fd_sc_hd__xnor2_1 _14807_ (.A(\cs_registers_i.pc_if_i[29] ),
    .B(_07697_),
    .Y(_07699_));
 sky130_fd_sc_hd__a21boi_0 _14808_ (.A1(net290),
    .A2(_07699_),
    .B1_N(_07614_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[29] ));
 sky130_fd_sc_hd__a21o_1 _14809_ (.A1(\cs_registers_i.pc_if_i[29] ),
    .A2(_07697_),
    .B1(\cs_registers_i.pc_if_i[30] ),
    .X(_07700_));
 sky130_fd_sc_hd__nand3_1 _14810_ (.A(\cs_registers_i.pc_if_i[29] ),
    .B(\cs_registers_i.pc_if_i[30] ),
    .C(_07697_),
    .Y(_07701_));
 sky130_fd_sc_hd__nand2_1 _14811_ (.A(_07700_),
    .B(_07701_),
    .Y(_07702_));
 sky130_fd_sc_hd__a21boi_0 _14812_ (.A1(_07330_),
    .A2(_07702_),
    .B1_N(_07619_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[30] ));
 sky130_fd_sc_hd__xnor2_1 _14813_ (.A(\cs_registers_i.pc_if_i[3] ),
    .B(_07649_),
    .Y(_07703_));
 sky130_fd_sc_hd__a21boi_0 _14814_ (.A1(net292),
    .A2(_07703_),
    .B1_N(_07456_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[3] ));
 sky130_fd_sc_hd__xor2_1 _14815_ (.A(\cs_registers_i.pc_if_i[31] ),
    .B(_07701_),
    .X(_07704_));
 sky130_fd_sc_hd__a21boi_0 _14816_ (.A1(_07330_),
    .A2(_07704_),
    .B1_N(_07624_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[31] ));
 sky130_fd_sc_hd__nand3_1 _14817_ (.A(\cs_registers_i.pc_if_i[3] ),
    .B(\cs_registers_i.pc_if_i[4] ),
    .C(_07649_),
    .Y(_07705_));
 sky130_fd_sc_hd__a21o_1 _14818_ (.A1(\cs_registers_i.pc_if_i[3] ),
    .A2(_07649_),
    .B1(\cs_registers_i.pc_if_i[4] ),
    .X(_07706_));
 sky130_fd_sc_hd__nand2_1 _14819_ (.A(_07705_),
    .B(_07706_),
    .Y(_07707_));
 sky130_fd_sc_hd__a21oi_1 _14820_ (.A1(net292),
    .A2(_07707_),
    .B1(_07452_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[4] ));
 sky130_fd_sc_hd__xor2_1 _14821_ (.A(\cs_registers_i.pc_if_i[5] ),
    .B(_07705_),
    .X(_07708_));
 sky130_fd_sc_hd__a21boi_0 _14822_ (.A1(net292),
    .A2(_07708_),
    .B1_N(_07448_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[5] ));
 sky130_fd_sc_hd__xnor2_1 _14823_ (.A(_07648_),
    .B(_07650_),
    .Y(_07709_));
 sky130_fd_sc_hd__a21boi_0 _14824_ (.A1(net292),
    .A2(_07709_),
    .B1_N(_07444_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[6] ));
 sky130_fd_sc_hd__xnor2_1 _14825_ (.A(\cs_registers_i.pc_if_i[7] ),
    .B(_07651_),
    .Y(_07710_));
 sky130_fd_sc_hd__a21boi_0 _14826_ (.A1(net292),
    .A2(_07710_),
    .B1_N(_07441_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[7] ));
 sky130_fd_sc_hd__nand2_1 _14827_ (.A(\cs_registers_i.pc_if_i[7] ),
    .B(_07651_),
    .Y(_07711_));
 sky130_fd_sc_hd__xnor2_1 _14828_ (.A(\cs_registers_i.pc_if_i[8] ),
    .B(_07711_),
    .Y(_07712_));
 sky130_fd_sc_hd__nand2_1 _14829_ (.A(net292),
    .B(_07712_),
    .Y(_07713_));
 sky130_fd_sc_hd__o31ai_1 _14830_ (.A1(net292),
    .A2(_07472_),
    .A3(_07475_),
    .B1(_07713_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[8] ));
 sky130_fd_sc_hd__xnor2_1 _14831_ (.A(\cs_registers_i.pc_if_i[9] ),
    .B(_07652_),
    .Y(_07714_));
 sky130_fd_sc_hd__nand2_1 _14832_ (.A(net292),
    .B(_07714_),
    .Y(_07715_));
 sky130_fd_sc_hd__o31ai_1 _14833_ (.A1(net292),
    .A2(_07465_),
    .A3(_07469_),
    .B1(_07715_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[9] ));
 sky130_fd_sc_hd__xor2_1 _14834_ (.A(\cs_registers_i.pc_if_i[10] ),
    .B(_07653_),
    .X(_07716_));
 sky130_fd_sc_hd__nand2_1 _14835_ (.A(net291),
    .B(_07716_),
    .Y(_07717_));
 sky130_fd_sc_hd__o31ai_1 _14836_ (.A1(net291),
    .A2(_07424_),
    .A3(_07437_),
    .B1(_07717_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[10] ));
 sky130_fd_sc_hd__o21ai_4 _14837_ (.A1(_11164_),
    .A2(_11201_),
    .B1(net293),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ));
 sky130_fd_sc_hd__mux2_1 _14838_ (.A0(net103),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[16] ));
 sky130_fd_sc_hd__mux2_1 _14839_ (.A0(net104),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[17] ));
 sky130_fd_sc_hd__mux2_1 _14840_ (.A0(net105),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[18] ));
 sky130_fd_sc_hd__mux2_1 _14841_ (.A0(net106),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[19] ));
 sky130_fd_sc_hd__mux2_1 _14842_ (.A0(net108),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[20] ));
 sky130_fd_sc_hd__mux2_1 _14843_ (.A0(net109),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[21] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1224 ();
 sky130_fd_sc_hd__mux2_1 _14845_ (.A0(net110),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[22] ));
 sky130_fd_sc_hd__mux2_1 _14846_ (.A0(net111),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[23] ));
 sky130_fd_sc_hd__mux2_1 _14847_ (.A0(net112),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[24] ));
 sky130_fd_sc_hd__mux2_1 _14848_ (.A0(net113),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[25] ));
 sky130_fd_sc_hd__mux2_1 _14849_ (.A0(net114),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[26] ));
 sky130_fd_sc_hd__mux2_1 _14850_ (.A0(net115),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[27] ));
 sky130_fd_sc_hd__mux2_1 _14851_ (.A0(net116),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[28] ));
 sky130_fd_sc_hd__mux2_1 _14852_ (.A0(net117),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[29] ));
 sky130_fd_sc_hd__mux2_1 _14853_ (.A0(net119),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[30] ));
 sky130_fd_sc_hd__mux2_1 _14854_ (.A0(net120),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[31] ));
 sky130_fd_sc_hd__mux2_1 _14855_ (.A0(net96),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[32] ));
 sky130_fd_sc_hd__mux2_1 _14856_ (.A0(net107),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[33] ));
 sky130_fd_sc_hd__mux2_1 _14857_ (.A0(net118),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[34] ));
 sky130_fd_sc_hd__mux2_1 _14858_ (.A0(net121),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[35] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1223 ();
 sky130_fd_sc_hd__mux2_1 _14860_ (.A0(net122),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[36] ));
 sky130_fd_sc_hd__mux2_1 _14861_ (.A0(net123),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[37] ));
 sky130_fd_sc_hd__mux2_1 _14862_ (.A0(net124),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[38] ));
 sky130_fd_sc_hd__mux2_1 _14863_ (.A0(net125),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[39] ));
 sky130_fd_sc_hd__mux2_1 _14864_ (.A0(net126),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[40] ));
 sky130_fd_sc_hd__mux2_1 _14865_ (.A0(net127),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[41] ));
 sky130_fd_sc_hd__mux2_1 _14866_ (.A0(net97),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[42] ));
 sky130_fd_sc_hd__mux2_1 _14867_ (.A0(net98),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[43] ));
 sky130_fd_sc_hd__mux2_1 _14868_ (.A0(net99),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[44] ));
 sky130_fd_sc_hd__mux2_1 _14869_ (.A0(net100),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[45] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1222 ();
 sky130_fd_sc_hd__mux2_1 _14871_ (.A0(net101),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[46] ));
 sky130_fd_sc_hd__mux2_1 _14872_ (.A0(net102),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[47] ));
 sky130_fd_sc_hd__mux2_1 _14873_ (.A0(net103),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[48] ));
 sky130_fd_sc_hd__mux2_1 _14874_ (.A0(net104),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[49] ));
 sky130_fd_sc_hd__mux2_1 _14875_ (.A0(net105),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[50] ));
 sky130_fd_sc_hd__mux2_1 _14876_ (.A0(net106),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[51] ));
 sky130_fd_sc_hd__mux2_1 _14877_ (.A0(net108),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[52] ));
 sky130_fd_sc_hd__mux2_1 _14878_ (.A0(net109),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[53] ));
 sky130_fd_sc_hd__mux2_1 _14879_ (.A0(net110),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[54] ));
 sky130_fd_sc_hd__mux2_1 _14880_ (.A0(net111),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[55] ));
 sky130_fd_sc_hd__mux2_1 _14881_ (.A0(net112),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[56] ));
 sky130_fd_sc_hd__mux2_1 _14882_ (.A0(net113),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[57] ));
 sky130_fd_sc_hd__mux2_1 _14883_ (.A0(net114),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[58] ));
 sky130_fd_sc_hd__mux2_1 _14884_ (.A0(net115),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[59] ));
 sky130_fd_sc_hd__mux2_1 _14885_ (.A0(net116),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[60] ));
 sky130_fd_sc_hd__mux2_1 _14886_ (.A0(net117),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[61] ));
 sky130_fd_sc_hd__mux2_1 _14887_ (.A0(net119),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[62] ));
 sky130_fd_sc_hd__mux2_1 _14888_ (.A0(net120),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[63] ));
 sky130_fd_sc_hd__o31ai_1 _14889_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .A2(_11130_),
    .A3(net1292),
    .B1(_07640_),
    .Y(_07721_));
 sky130_fd_sc_hd__nor2_1 _14890_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .B(_07721_),
    .Y(_07722_));
 sky130_fd_sc_hd__a211oi_1 _14891_ (.A1(_11160_),
    .A2(net1292),
    .B1(_07722_),
    .C1(net1026),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ));
 sky130_fd_sc_hd__o21ai_0 _14892_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .A2(_11130_),
    .B1(_07636_),
    .Y(_07723_));
 sky130_fd_sc_hd__nor3_1 _14893_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .B(_11130_),
    .C(_07638_),
    .Y(_07724_));
 sky130_fd_sc_hd__a221oi_1 _14894_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .A2(net1292),
    .B1(_07723_),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .C1(_07724_),
    .Y(_07725_));
 sky130_fd_sc_hd__nor2_1 _14895_ (.A(net1026),
    .B(_07725_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ));
 sky130_fd_sc_hd__a21oi_1 _14896_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .A2(_11139_),
    .B1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .Y(_07726_));
 sky130_fd_sc_hd__nor3_1 _14897_ (.A(net1026),
    .B(net1292),
    .C(_07726_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1221 ();
 sky130_fd_sc_hd__mux2_1 _14899_ (.A0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10] ),
    .A1(_07439_),
    .S(_10994_),
    .X(net219));
 sky130_fd_sc_hd__mux2_1 _14900_ (.A0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11] ),
    .A1(_07488_),
    .S(_10994_),
    .X(net220));
 sky130_fd_sc_hd__mux2_4 _14901_ (.A0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12] ),
    .A1(_07495_),
    .S(_10994_),
    .X(net221));
 sky130_fd_sc_hd__mux2_1 _14902_ (.A0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13] ),
    .A1(_07503_),
    .S(_10994_),
    .X(net222));
 sky130_fd_sc_hd__nor2_1 _14903_ (.A(_10994_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14] ),
    .Y(_07728_));
 sky130_fd_sc_hd__a21oi_2 _14904_ (.A1(_07509_),
    .A2(_10994_),
    .B1(_07728_),
    .Y(net223));
 sky130_fd_sc_hd__nor2_1 _14905_ (.A(_10994_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15] ),
    .Y(_07729_));
 sky130_fd_sc_hd__a21oi_2 _14906_ (.A1(_10994_),
    .A2(_07517_),
    .B1(_07729_),
    .Y(net224));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1218 ();
 sky130_fd_sc_hd__nand2_1 _14910_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16] ),
    .Y(_07733_));
 sky130_fd_sc_hd__o21ai_1 _14911_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07525_),
    .B1(_07733_),
    .Y(net225));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1217 ();
 sky130_fd_sc_hd__nand2_1 _14913_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17] ),
    .Y(_07735_));
 sky130_fd_sc_hd__o21ai_2 _14914_ (.A1(_07530_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B1(_07735_),
    .Y(net226));
 sky130_fd_sc_hd__mux2_4 _14915_ (.A0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18] ),
    .A1(_07541_),
    .S(_10994_),
    .X(net227));
 sky130_fd_sc_hd__nand2_1 _14916_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19] ),
    .Y(_07736_));
 sky130_fd_sc_hd__o21ai_1 _14917_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07549_),
    .B1(_07736_),
    .Y(net228));
 sky130_fd_sc_hd__nand2_1 _14918_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20] ),
    .Y(_07737_));
 sky130_fd_sc_hd__o21ai_0 _14919_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07556_),
    .B1(_07737_),
    .Y(net229));
 sky130_fd_sc_hd__nand2_1 _14920_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21] ),
    .Y(_07738_));
 sky130_fd_sc_hd__o21ai_1 _14921_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07562_),
    .B1(_07738_),
    .Y(net230));
 sky130_fd_sc_hd__nand2_1 _14922_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22] ),
    .Y(_07739_));
 sky130_fd_sc_hd__o21ai_2 _14923_ (.A1(_07569_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B1(_07739_),
    .Y(net231));
 sky130_fd_sc_hd__nand2_1 _14924_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23] ),
    .Y(_07740_));
 sky130_fd_sc_hd__o21ai_2 _14925_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07576_),
    .B1(_07740_),
    .Y(net232));
 sky130_fd_sc_hd__nand2_1 _14926_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24] ),
    .Y(_07741_));
 sky130_fd_sc_hd__o21ai_2 _14927_ (.A1(_07582_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B1(_07741_),
    .Y(net233));
 sky130_fd_sc_hd__mux2_4 _14928_ (.A0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25] ),
    .A1(_07589_),
    .S(_10994_),
    .X(net234));
 sky130_fd_sc_hd__nand2_1 _14929_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26] ),
    .Y(_07742_));
 sky130_fd_sc_hd__o21ai_2 _14930_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07594_),
    .B1(_07742_),
    .Y(net235));
 sky130_fd_sc_hd__nand2_1 _14931_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27] ),
    .Y(_07743_));
 sky130_fd_sc_hd__o21ai_2 _14932_ (.A1(_07602_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B1(_07743_),
    .Y(net236));
 sky130_fd_sc_hd__nand2_1 _14933_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28] ),
    .Y(_07744_));
 sky130_fd_sc_hd__o21ai_2 _14934_ (.A1(_07610_),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B1(_07744_),
    .Y(net237));
 sky130_fd_sc_hd__mux2_4 _14935_ (.A0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29] ),
    .A1(_07615_),
    .S(_10994_),
    .X(net238));
 sky130_fd_sc_hd__nand2_1 _14936_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2] ),
    .Y(_07745_));
 sky130_fd_sc_hd__o21ai_2 _14937_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07461_),
    .B1(_07745_),
    .Y(net239));
 sky130_fd_sc_hd__nand2_1 _14938_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30] ),
    .Y(_07746_));
 sky130_fd_sc_hd__o21ai_4 _14939_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07620_),
    .B1(_07746_),
    .Y(net240));
 sky130_fd_sc_hd__nand2_1 _14940_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31] ),
    .Y(_07747_));
 sky130_fd_sc_hd__o21ai_2 _14941_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07625_),
    .B1(_07747_),
    .Y(net241));
 sky130_fd_sc_hd__nand2_1 _14942_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3] ),
    .Y(_07748_));
 sky130_fd_sc_hd__o21ai_2 _14943_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07457_),
    .B1(_07748_),
    .Y(net242));
 sky130_fd_sc_hd__nand2_1 _14944_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4] ),
    .Y(_07749_));
 sky130_fd_sc_hd__o21ai_2 _14945_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07453_),
    .B1(_07749_),
    .Y(net243));
 sky130_fd_sc_hd__nand2_1 _14946_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5] ),
    .Y(_07750_));
 sky130_fd_sc_hd__o21ai_2 _14947_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07449_),
    .B1(_07750_),
    .Y(net244));
 sky130_fd_sc_hd__nand2_1 _14948_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6] ),
    .Y(_07751_));
 sky130_fd_sc_hd__o21ai_2 _14949_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07445_),
    .B1(_07751_),
    .Y(net245));
 sky130_fd_sc_hd__nand2_1 _14950_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7] ),
    .Y(_07752_));
 sky130_fd_sc_hd__o21ai_1 _14951_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .A2(_07442_),
    .B1(_07752_),
    .Y(net246));
 sky130_fd_sc_hd__mux2_1 _14952_ (.A0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8] ),
    .A1(_07477_),
    .S(_10994_),
    .X(net247));
 sky130_fd_sc_hd__mux2_1 _14953_ (.A0(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9] ),
    .A1(_07471_),
    .S(_10994_),
    .X(net248));
 sky130_fd_sc_hd__clkinvlp_4 _14954_ (.A(_07332_),
    .Y(net249));
 sky130_fd_sc_hd__nand2b_1 _14955_ (.A_N(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .B(net128),
    .Y(_07753_));
 sky130_fd_sc_hd__a22o_1 _14956_ (.A1(net95),
    .A2(net249),
    .B1(_07753_),
    .B2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ));
 sky130_fd_sc_hd__a31oi_1 _14957_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .A2(net95),
    .A3(net249),
    .B1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .Y(_07754_));
 sky130_fd_sc_hd__a21oi_1 _14958_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .A2(net128),
    .B1(_07754_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ));
 sky130_fd_sc_hd__nor2_8 _14959_ (.A(net95),
    .B(_07458_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ));
 sky130_fd_sc_hd__nor2_1 _14960_ (.A(net95),
    .B(_07332_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ));
 sky130_fd_sc_hd__nand2_8 _14961_ (.A(_10838_),
    .B(\if_stage_i.compressed_decoder_i.instr_i[0] ),
    .Y(_07755_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1214 ();
 sky130_fd_sc_hd__nor2_2 _14965_ (.A(_11082_),
    .B(\if_stage_i.compressed_decoder_i.instr_i[6] ),
    .Y(_07759_));
 sky130_fd_sc_hd__nor4b_4 _14966_ (.A(_11091_),
    .B(_11095_),
    .C(\if_stage_i.compressed_decoder_i.instr_i[4] ),
    .D_N(_07759_),
    .Y(_07760_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1211 ();
 sky130_fd_sc_hd__nand2_4 _14970_ (.A(_11061_),
    .B(_11067_),
    .Y(_07764_));
 sky130_fd_sc_hd__nor2_1 _14971_ (.A(_11053_),
    .B(_07764_),
    .Y(_07765_));
 sky130_fd_sc_hd__a21oi_1 _14972_ (.A1(_11073_),
    .A2(_11078_),
    .B1(_11114_),
    .Y(_07766_));
 sky130_fd_sc_hd__nand2_4 _14973_ (.A(_11053_),
    .B(_11059_),
    .Y(_07767_));
 sky130_fd_sc_hd__nor2_8 _14974_ (.A(_11067_),
    .B(_07767_),
    .Y(_07768_));
 sky130_fd_sc_hd__a32oi_4 _14975_ (.A1(_11114_),
    .A2(_07760_),
    .A3(_07765_),
    .B1(_07766_),
    .B2(_07768_),
    .Y(_07769_));
 sky130_fd_sc_hd__nand2_4 _14976_ (.A(_11053_),
    .B(_11061_),
    .Y(_07770_));
 sky130_fd_sc_hd__nor2_8 _14977_ (.A(_10839_),
    .B(\if_stage_i.compressed_decoder_i.instr_i[0] ),
    .Y(_07771_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1210 ();
 sky130_fd_sc_hd__nand2_1 _14979_ (.A(_07770_),
    .B(_07771_),
    .Y(_07773_));
 sky130_fd_sc_hd__or4_4 _14980_ (.A(_11074_),
    .B(_11078_),
    .C(_11103_),
    .D(\if_stage_i.compressed_decoder_i.instr_i[9] ),
    .X(_07774_));
 sky130_fd_sc_hd__nor2_2 _14981_ (.A(_11107_),
    .B(_07774_),
    .Y(_07775_));
 sky130_fd_sc_hd__nand2_4 _14982_ (.A(_11053_),
    .B(_11067_),
    .Y(_07776_));
 sky130_fd_sc_hd__a31oi_2 _14983_ (.A1(_11114_),
    .A2(_07775_),
    .A3(_07759_),
    .B1(_07776_),
    .Y(_07777_));
 sky130_fd_sc_hd__nor2_4 _14984_ (.A(_11055_),
    .B(_11068_),
    .Y(_07778_));
 sky130_fd_sc_hd__nand2_4 _14985_ (.A(_11059_),
    .B(_07778_),
    .Y(_07779_));
 sky130_fd_sc_hd__nor2_4 _14986_ (.A(_10838_),
    .B(\if_stage_i.compressed_decoder_i.instr_i[0] ),
    .Y(_07780_));
 sky130_fd_sc_hd__or2_0 _14987_ (.A(_11107_),
    .B(_07774_),
    .X(_07781_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1209 ();
 sky130_fd_sc_hd__a31oi_1 _14989_ (.A1(_11114_),
    .A2(_07775_),
    .A3(_07760_),
    .B1(_11067_),
    .Y(_07783_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1208 ();
 sky130_fd_sc_hd__o221ai_1 _14991_ (.A1(_11068_),
    .A2(_07781_),
    .B1(_07783_),
    .B2(_11061_),
    .C1(_11053_),
    .Y(_07785_));
 sky130_fd_sc_hd__o211ai_1 _14992_ (.A1(_11115_),
    .A2(_07779_),
    .B1(_07780_),
    .C1(_07785_),
    .Y(_07786_));
 sky130_fd_sc_hd__o221ai_4 _14993_ (.A1(_07755_),
    .A2(_07769_),
    .B1(_07773_),
    .B2(_07777_),
    .C1(_07786_),
    .Y(\if_stage_i.compressed_decoder_i.illegal_instr_o ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1206 ();
 sky130_fd_sc_hd__nand2_1 _14996_ (.A(_11059_),
    .B(_11068_),
    .Y(_07789_));
 sky130_fd_sc_hd__o21ai_0 _14997_ (.A1(_10839_),
    .A2(_07789_),
    .B1(_11053_),
    .Y(_07790_));
 sky130_fd_sc_hd__nand2_1 _14998_ (.A(_10844_),
    .B(_07790_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[0] ));
 sky130_fd_sc_hd__o21ai_0 _14999_ (.A1(_11061_),
    .A2(_07755_),
    .B1(_11074_),
    .Y(_07791_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1205 ();
 sky130_fd_sc_hd__nand2_1 _15001_ (.A(_10844_),
    .B(_11067_),
    .Y(_07793_));
 sky130_fd_sc_hd__o21ai_0 _15002_ (.A1(_10844_),
    .A2(_07789_),
    .B1(_07793_),
    .Y(_07794_));
 sky130_fd_sc_hd__a21oi_1 _15003_ (.A1(_10838_),
    .A2(_07794_),
    .B1(_11074_),
    .Y(_07795_));
 sky130_fd_sc_hd__nand2_2 _15004_ (.A(_10839_),
    .B(_10844_),
    .Y(_07796_));
 sky130_fd_sc_hd__nand2_1 _15005_ (.A(_07760_),
    .B(_07768_),
    .Y(_07797_));
 sky130_fd_sc_hd__nor2_1 _15006_ (.A(_07796_),
    .B(_07797_),
    .Y(_07798_));
 sky130_fd_sc_hd__a211oi_1 _15007_ (.A1(_11055_),
    .A2(_07791_),
    .B1(_07795_),
    .C1(_07798_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[10] ));
 sky130_fd_sc_hd__nor2_4 _15008_ (.A(_10839_),
    .B(_10844_),
    .Y(_07799_));
 sky130_fd_sc_hd__nor2_2 _15009_ (.A(_11055_),
    .B(_11061_),
    .Y(_07800_));
 sky130_fd_sc_hd__nand2_2 _15010_ (.A(_11068_),
    .B(_07800_),
    .Y(_07801_));
 sky130_fd_sc_hd__and2_2 _15011_ (.A(_11074_),
    .B(_11078_),
    .X(_07802_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1204 ();
 sky130_fd_sc_hd__nand2_2 _15013_ (.A(_11115_),
    .B(_07802_),
    .Y(_07804_));
 sky130_fd_sc_hd__nor2_1 _15014_ (.A(_07801_),
    .B(_07804_),
    .Y(_07805_));
 sky130_fd_sc_hd__nand2_1 _15015_ (.A(_07799_),
    .B(_07805_),
    .Y(_07806_));
 sky130_fd_sc_hd__nor2_1 _15016_ (.A(\if_stage_i.compressed_decoder_i.instr_i[0] ),
    .B(_07797_),
    .Y(_07807_));
 sky130_fd_sc_hd__nor2_1 _15017_ (.A(_10838_),
    .B(_07807_),
    .Y(_07808_));
 sky130_fd_sc_hd__nor2_1 _15018_ (.A(_10844_),
    .B(_11061_),
    .Y(_07809_));
 sky130_fd_sc_hd__nor2_1 _15019_ (.A(\if_stage_i.compressed_decoder_i.instr_i[0] ),
    .B(_07776_),
    .Y(_07810_));
 sky130_fd_sc_hd__a211oi_1 _15020_ (.A1(_07776_),
    .A2(_07809_),
    .B1(_07810_),
    .C1(_10839_),
    .Y(_07811_));
 sky130_fd_sc_hd__o21ai_0 _15021_ (.A1(_07808_),
    .A2(_07811_),
    .B1(_11078_),
    .Y(_07812_));
 sky130_fd_sc_hd__nand2_1 _15022_ (.A(_07806_),
    .B(_07812_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[11] ));
 sky130_fd_sc_hd__nor2_4 _15023_ (.A(_11061_),
    .B(_07776_),
    .Y(_07813_));
 sky130_fd_sc_hd__nor2_1 _15024_ (.A(_10844_),
    .B(_11114_),
    .Y(_07814_));
 sky130_fd_sc_hd__a21oi_1 _15025_ (.A1(_10844_),
    .A2(_07813_),
    .B1(_07814_),
    .Y(_07815_));
 sky130_fd_sc_hd__nand2_1 _15026_ (.A(_11082_),
    .B(\if_stage_i.compressed_decoder_i.instr_i[6] ),
    .Y(_07816_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1203 ();
 sky130_fd_sc_hd__a31oi_1 _15028_ (.A1(_11114_),
    .A2(_07802_),
    .A3(_07816_),
    .B1(_11067_),
    .Y(_07818_));
 sky130_fd_sc_hd__nor2_4 _15029_ (.A(_11053_),
    .B(_11061_),
    .Y(_07819_));
 sky130_fd_sc_hd__nand2_4 _15030_ (.A(_07779_),
    .B(_07799_),
    .Y(_07820_));
 sky130_fd_sc_hd__a21oi_1 _15031_ (.A1(_11114_),
    .A2(_07819_),
    .B1(_07820_),
    .Y(_07821_));
 sky130_fd_sc_hd__nand2b_1 _15032_ (.A_N(_07774_),
    .B(_11107_),
    .Y(_07822_));
 sky130_fd_sc_hd__a21oi_1 _15033_ (.A1(_11091_),
    .A2(_07822_),
    .B1(_11068_),
    .Y(_07823_));
 sky130_fd_sc_hd__o21ai_0 _15034_ (.A1(_11053_),
    .A2(_07823_),
    .B1(_11061_),
    .Y(_07824_));
 sky130_fd_sc_hd__o211ai_1 _15035_ (.A1(_11055_),
    .A2(_07818_),
    .B1(_07821_),
    .C1(_07824_),
    .Y(_07825_));
 sky130_fd_sc_hd__o221ai_2 _15036_ (.A1(_11114_),
    .A2(\if_stage_i.compressed_decoder_i.instr_o[0] ),
    .B1(_07815_),
    .B2(_10838_),
    .C1(_07825_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[12] ));
 sky130_fd_sc_hd__and3_1 _15037_ (.A(_11068_),
    .B(_11078_),
    .C(_07800_),
    .X(_07826_));
 sky130_fd_sc_hd__o21ai_0 _15038_ (.A1(_11086_),
    .A2(_11115_),
    .B1(_11074_),
    .Y(_07827_));
 sky130_fd_sc_hd__nand3_4 _15039_ (.A(_11055_),
    .B(_11061_),
    .C(_11067_),
    .Y(_07828_));
 sky130_fd_sc_hd__nor2b_4 _15040_ (.A(_07774_),
    .B_N(_11107_),
    .Y(_07829_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1202 ();
 sky130_fd_sc_hd__nor2_2 _15042_ (.A(_07828_),
    .B(_07829_),
    .Y(_07831_));
 sky130_fd_sc_hd__a222oi_1 _15043_ (.A1(_11115_),
    .A2(_07819_),
    .B1(_07826_),
    .B2(_07827_),
    .C1(_07831_),
    .C2(_11095_),
    .Y(_07832_));
 sky130_fd_sc_hd__a21oi_1 _15044_ (.A1(_10839_),
    .A2(_11055_),
    .B1(_10844_),
    .Y(_07833_));
 sky130_fd_sc_hd__o22ai_2 _15045_ (.A1(_07820_),
    .A2(_07832_),
    .B1(_07833_),
    .B2(_07800_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[13] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1201 ();
 sky130_fd_sc_hd__nor2_2 _15047_ (.A(\if_stage_i.compressed_decoder_i.instr_i[0] ),
    .B(_11055_),
    .Y(_07835_));
 sky130_fd_sc_hd__o21ai_0 _15048_ (.A1(_11115_),
    .A2(_07759_),
    .B1(_07802_),
    .Y(_07836_));
 sky130_fd_sc_hd__a222oi_1 _15049_ (.A1(_11115_),
    .A2(_07819_),
    .B1(_07836_),
    .B2(_07768_),
    .C1(_07831_),
    .C2(\if_stage_i.compressed_decoder_i.instr_i[4] ),
    .Y(_07837_));
 sky130_fd_sc_hd__o32ai_1 _15050_ (.A1(_11059_),
    .A2(_07799_),
    .A3(_07835_),
    .B1(_07820_),
    .B2(_07837_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[14] ));
 sky130_fd_sc_hd__nand2b_1 _15051_ (.A_N(_07760_),
    .B(_11114_),
    .Y(_07838_));
 sky130_fd_sc_hd__a21oi_1 _15052_ (.A1(_11103_),
    .A2(_07838_),
    .B1(_11067_),
    .Y(_07839_));
 sky130_fd_sc_hd__o22ai_1 _15053_ (.A1(_11053_),
    .A2(_11067_),
    .B1(_07767_),
    .B2(_07839_),
    .Y(_07840_));
 sky130_fd_sc_hd__nand2_1 _15054_ (.A(_07780_),
    .B(_07840_),
    .Y(_07841_));
 sky130_fd_sc_hd__inv_1 _15055_ (.A(_07841_),
    .Y(_07842_));
 sky130_fd_sc_hd__nor3_1 _15056_ (.A(_11115_),
    .B(_07801_),
    .C(_07816_),
    .Y(_07843_));
 sky130_fd_sc_hd__nand2_4 _15057_ (.A(_11055_),
    .B(_11059_),
    .Y(_07844_));
 sky130_fd_sc_hd__nand2_1 _15058_ (.A(_07768_),
    .B(_07802_),
    .Y(_07845_));
 sky130_fd_sc_hd__a21oi_1 _15059_ (.A1(_07844_),
    .A2(_07845_),
    .B1(_11114_),
    .Y(_07846_));
 sky130_fd_sc_hd__a221oi_1 _15060_ (.A1(_11082_),
    .A2(_07831_),
    .B1(_07843_),
    .B2(_11103_),
    .C1(_07846_),
    .Y(_07847_));
 sky130_fd_sc_hd__nand2_1 _15061_ (.A(_11074_),
    .B(_11078_),
    .Y(_07848_));
 sky130_fd_sc_hd__a21oi_1 _15062_ (.A1(_11114_),
    .A2(_07816_),
    .B1(_07848_),
    .Y(_07849_));
 sky130_fd_sc_hd__a21oi_1 _15063_ (.A1(_11068_),
    .A2(_07849_),
    .B1(_11055_),
    .Y(_07850_));
 sky130_fd_sc_hd__o21ai_1 _15064_ (.A1(_11061_),
    .A2(_07850_),
    .B1(_07764_),
    .Y(_07851_));
 sky130_fd_sc_hd__a21oi_1 _15065_ (.A1(_07847_),
    .A2(_07851_),
    .B1(_07755_),
    .Y(_07852_));
 sky130_fd_sc_hd__a21oi_1 _15066_ (.A1(_07841_),
    .A2(_07847_),
    .B1(_07813_),
    .Y(_07853_));
 sky130_fd_sc_hd__o22ai_1 _15067_ (.A1(_07842_),
    .A2(_07852_),
    .B1(_07853_),
    .B2(_11103_),
    .Y(_07854_));
 sky130_fd_sc_hd__nor2_2 _15068_ (.A(_11055_),
    .B(_11059_),
    .Y(_07855_));
 sky130_fd_sc_hd__nor2_1 _15069_ (.A(_11067_),
    .B(_07855_),
    .Y(_07856_));
 sky130_fd_sc_hd__a21oi_1 _15070_ (.A1(_11103_),
    .A2(_07855_),
    .B1(_07856_),
    .Y(_07857_));
 sky130_fd_sc_hd__nand2_4 _15071_ (.A(_10838_),
    .B(_10844_),
    .Y(_07858_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1200 ();
 sky130_fd_sc_hd__o21ai_0 _15073_ (.A1(_10844_),
    .A2(_11067_),
    .B1(_07854_),
    .Y(_07860_));
 sky130_fd_sc_hd__nand2_1 _15074_ (.A(_10839_),
    .B(_07860_),
    .Y(_07861_));
 sky130_fd_sc_hd__o221ai_1 _15075_ (.A1(_10844_),
    .A2(_07854_),
    .B1(_07857_),
    .B2(_07858_),
    .C1(_07861_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[15] ));
 sky130_fd_sc_hd__mux2_1 _15076_ (.A0(_10842_),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[0] ),
    .S(net451),
    .X(_07862_));
 sky130_fd_sc_hd__a21oi_2 _15077_ (.A1(_11059_),
    .A2(_11068_),
    .B1(_11055_),
    .Y(_07863_));
 sky130_fd_sc_hd__o22ai_1 _15078_ (.A1(_11107_),
    .A2(_07770_),
    .B1(_07862_),
    .B2(_07863_),
    .Y(_07864_));
 sky130_fd_sc_hd__nand2_2 _15079_ (.A(_10844_),
    .B(_11053_),
    .Y(_07865_));
 sky130_fd_sc_hd__or3_1 _15080_ (.A(_11067_),
    .B(_11115_),
    .C(_07760_),
    .X(_07866_));
 sky130_fd_sc_hd__a21oi_1 _15081_ (.A1(_11107_),
    .A2(_07866_),
    .B1(_11061_),
    .Y(_07867_));
 sky130_fd_sc_hd__nand2_1 _15082_ (.A(_07865_),
    .B(_07862_),
    .Y(_07868_));
 sky130_fd_sc_hd__o21ai_0 _15083_ (.A1(_07865_),
    .A2(_07867_),
    .B1(_07868_),
    .Y(_07869_));
 sky130_fd_sc_hd__a31oi_1 _15084_ (.A1(_07768_),
    .A2(_07802_),
    .A3(_07862_),
    .B1(_07819_),
    .Y(_07870_));
 sky130_fd_sc_hd__nor2_1 _15085_ (.A(_07774_),
    .B(_07828_),
    .Y(_07871_));
 sky130_fd_sc_hd__o21ai_0 _15086_ (.A1(_07843_),
    .A2(_07871_),
    .B1(_11107_),
    .Y(_07872_));
 sky130_fd_sc_hd__o221ai_1 _15087_ (.A1(_11086_),
    .A2(_07828_),
    .B1(_07870_),
    .B2(_11114_),
    .C1(_07872_),
    .Y(_07873_));
 sky130_fd_sc_hd__nor2_2 _15088_ (.A(_07813_),
    .B(_07755_),
    .Y(_07874_));
 sky130_fd_sc_hd__inv_1 _15089_ (.A(_07851_),
    .Y(_07875_));
 sky130_fd_sc_hd__a21oi_1 _15090_ (.A1(_11107_),
    .A2(_07875_),
    .B1(_10844_),
    .Y(_07876_));
 sky130_fd_sc_hd__nor2_1 _15091_ (.A(_10839_),
    .B(_07876_),
    .Y(_07877_));
 sky130_fd_sc_hd__a221oi_1 _15092_ (.A1(_10839_),
    .A2(_07869_),
    .B1(_07873_),
    .B2(_07874_),
    .C1(_07877_),
    .Y(_07878_));
 sky130_fd_sc_hd__a21oi_1 _15093_ (.A1(_07771_),
    .A2(_07864_),
    .B1(_07878_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[16] ));
 sky130_fd_sc_hd__o21ai_4 _15094_ (.A1(_07828_),
    .A2(_07829_),
    .B1(_07844_),
    .Y(_07879_));
 sky130_fd_sc_hd__mux2i_4 _15095_ (.A0(_10836_),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[1] ),
    .S(\cs_registers_i.pc_if_i[1] ),
    .Y(_07880_));
 sky130_fd_sc_hd__nand4_1 _15096_ (.A(_11082_),
    .B(\if_stage_i.compressed_decoder_i.instr_i[6] ),
    .C(\if_stage_i.compressed_decoder_i.instr_i[9] ),
    .D(_11114_),
    .Y(_07881_));
 sky130_fd_sc_hd__o21ai_0 _15097_ (.A1(_07804_),
    .A2(_07880_),
    .B1(_07881_),
    .Y(_07882_));
 sky130_fd_sc_hd__a222oi_1 _15098_ (.A1(\if_stage_i.compressed_decoder_i.instr_i[9] ),
    .A2(_07875_),
    .B1(_07879_),
    .B2(_11115_),
    .C1(_07882_),
    .C2(_07768_),
    .Y(_07883_));
 sky130_fd_sc_hd__o2111ai_1 _15099_ (.A1(_11067_),
    .A2(_07838_),
    .B1(\if_stage_i.compressed_decoder_i.instr_i[9] ),
    .C1(_11053_),
    .D1(_11059_),
    .Y(_07884_));
 sky130_fd_sc_hd__o21ai_0 _15100_ (.A1(_11053_),
    .A2(_07880_),
    .B1(_07884_),
    .Y(_07885_));
 sky130_fd_sc_hd__nand2_4 _15101_ (.A(_11053_),
    .B(_07789_),
    .Y(_07886_));
 sky130_fd_sc_hd__nor2_2 _15102_ (.A(_10838_),
    .B(_10844_),
    .Y(_07887_));
 sky130_fd_sc_hd__a21oi_2 _15103_ (.A1(_07771_),
    .A2(_07886_),
    .B1(_07887_),
    .Y(_07888_));
 sky130_fd_sc_hd__nand2_1 _15104_ (.A(\if_stage_i.compressed_decoder_i.instr_i[9] ),
    .B(_07771_),
    .Y(_07889_));
 sky130_fd_sc_hd__o22ai_1 _15105_ (.A1(_07880_),
    .A2(_07888_),
    .B1(_07889_),
    .B2(_07770_),
    .Y(_07890_));
 sky130_fd_sc_hd__a21oi_1 _15106_ (.A1(_07780_),
    .A2(_07885_),
    .B1(_07890_),
    .Y(_07891_));
 sky130_fd_sc_hd__o21ai_0 _15107_ (.A1(_07755_),
    .A2(_07883_),
    .B1(_07891_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[17] ));
 sky130_fd_sc_hd__a21oi_2 _15108_ (.A1(_11115_),
    .A2(_07879_),
    .B1(_07813_),
    .Y(_07892_));
 sky130_fd_sc_hd__nand2_2 _15109_ (.A(_11061_),
    .B(_11068_),
    .Y(_07893_));
 sky130_fd_sc_hd__nor2_1 _15110_ (.A(net449),
    .B(_11089_),
    .Y(_07894_));
 sky130_fd_sc_hd__a21oi_4 _15111_ (.A1(net449),
    .A2(_11118_),
    .B1(_07894_),
    .Y(_07895_));
 sky130_fd_sc_hd__o21ai_0 _15112_ (.A1(_07804_),
    .A2(_07895_),
    .B1(_07768_),
    .Y(_07896_));
 sky130_fd_sc_hd__a31oi_1 _15113_ (.A1(_07892_),
    .A2(_07893_),
    .A3(_07896_),
    .B1(_07755_),
    .Y(_07897_));
 sky130_fd_sc_hd__a32oi_1 _15114_ (.A1(_11074_),
    .A2(_07800_),
    .A3(_07866_),
    .B1(_07895_),
    .B2(_11055_),
    .Y(_07898_));
 sky130_fd_sc_hd__nor2_1 _15115_ (.A(_07796_),
    .B(_07898_),
    .Y(_07899_));
 sky130_fd_sc_hd__o22ai_2 _15116_ (.A1(_11074_),
    .A2(_07779_),
    .B1(_07897_),
    .B2(_07899_),
    .Y(_07900_));
 sky130_fd_sc_hd__a21oi_1 _15117_ (.A1(_07776_),
    .A2(_07895_),
    .B1(_07855_),
    .Y(_07901_));
 sky130_fd_sc_hd__nand2_1 _15118_ (.A(\if_stage_i.compressed_decoder_i.instr_i[0] ),
    .B(_07895_),
    .Y(_07902_));
 sky130_fd_sc_hd__nand2_1 _15119_ (.A(_07900_),
    .B(_07902_),
    .Y(_07903_));
 sky130_fd_sc_hd__nand2_1 _15120_ (.A(_10839_),
    .B(_07903_),
    .Y(_07904_));
 sky130_fd_sc_hd__o221ai_1 _15121_ (.A1(_10844_),
    .A2(_07900_),
    .B1(_07901_),
    .B2(_07858_),
    .C1(_07904_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[18] ));
 sky130_fd_sc_hd__mux2i_4 _15122_ (.A0(_11093_),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[3] ),
    .S(net450),
    .Y(_07905_));
 sky130_fd_sc_hd__a21oi_1 _15123_ (.A1(_11078_),
    .A2(_07838_),
    .B1(_11067_),
    .Y(_07906_));
 sky130_fd_sc_hd__o22ai_1 _15124_ (.A1(_11053_),
    .A2(_07905_),
    .B1(_07906_),
    .B2(_07767_),
    .Y(_07907_));
 sky130_fd_sc_hd__o22ai_1 _15125_ (.A1(_10839_),
    .A2(_07892_),
    .B1(_07905_),
    .B2(_07806_),
    .Y(_07908_));
 sky130_fd_sc_hd__a21oi_1 _15126_ (.A1(_07780_),
    .A2(_07907_),
    .B1(_07908_),
    .Y(_07909_));
 sky130_fd_sc_hd__o21ai_0 _15127_ (.A1(_11078_),
    .A2(_07779_),
    .B1(_07858_),
    .Y(_07910_));
 sky130_fd_sc_hd__o22ai_1 _15128_ (.A1(_07888_),
    .A2(_07905_),
    .B1(_07909_),
    .B2(_07910_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[19] ));
 sky130_fd_sc_hd__a22oi_1 _15129_ (.A1(_07799_),
    .A2(_07805_),
    .B1(_07886_),
    .B2(_07771_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[1] ));
 sky130_fd_sc_hd__nor2_1 _15130_ (.A(_11091_),
    .B(_07779_),
    .Y(_07911_));
 sky130_fd_sc_hd__nand2_1 _15131_ (.A(_11068_),
    .B(_11091_),
    .Y(_07912_));
 sky130_fd_sc_hd__nor2_1 _15132_ (.A(net449),
    .B(_11097_),
    .Y(_07913_));
 sky130_fd_sc_hd__a21oi_2 _15133_ (.A1(net449),
    .A2(_11120_),
    .B1(_07913_),
    .Y(_07914_));
 sky130_fd_sc_hd__a31oi_1 _15134_ (.A1(_11115_),
    .A2(_07775_),
    .A3(_07760_),
    .B1(_11091_),
    .Y(_07915_));
 sky130_fd_sc_hd__nor2_1 _15135_ (.A(_07767_),
    .B(_07915_),
    .Y(_07916_));
 sky130_fd_sc_hd__a21oi_1 _15136_ (.A1(_11055_),
    .A2(_07914_),
    .B1(_07916_),
    .Y(_07917_));
 sky130_fd_sc_hd__o21ai_0 _15137_ (.A1(_07770_),
    .A2(_07912_),
    .B1(_07917_),
    .Y(_07918_));
 sky130_fd_sc_hd__nor2_1 _15138_ (.A(_11114_),
    .B(_07848_),
    .Y(_07919_));
 sky130_fd_sc_hd__nand2_1 _15139_ (.A(_11067_),
    .B(_07855_),
    .Y(_07920_));
 sky130_fd_sc_hd__o21ai_1 _15140_ (.A1(_07801_),
    .A2(_07919_),
    .B1(_07920_),
    .Y(_07921_));
 sky130_fd_sc_hd__a22oi_1 _15141_ (.A1(_11091_),
    .A2(_07921_),
    .B1(_07914_),
    .B2(_07805_),
    .Y(_07922_));
 sky130_fd_sc_hd__a21oi_1 _15142_ (.A1(_07892_),
    .A2(_07922_),
    .B1(_07755_),
    .Y(_07923_));
 sky130_fd_sc_hd__a21oi_1 _15143_ (.A1(_07780_),
    .A2(_07918_),
    .B1(_07923_),
    .Y(_07924_));
 sky130_fd_sc_hd__nand2_1 _15144_ (.A(_07886_),
    .B(_07914_),
    .Y(_07925_));
 sky130_fd_sc_hd__o21ai_0 _15145_ (.A1(_07770_),
    .A2(_07912_),
    .B1(_07925_),
    .Y(_07926_));
 sky130_fd_sc_hd__a22oi_1 _15146_ (.A1(_07887_),
    .A2(_07914_),
    .B1(_07926_),
    .B2(_07771_),
    .Y(_07927_));
 sky130_fd_sc_hd__o21ai_0 _15147_ (.A1(_07911_),
    .A2(_07924_),
    .B1(_07927_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[20] ));
 sky130_fd_sc_hd__mux2i_2 _15148_ (.A0(_11080_),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[5] ),
    .S(net450),
    .Y(_07928_));
 sky130_fd_sc_hd__nand2_2 _15149_ (.A(_10839_),
    .B(_07865_),
    .Y(_07929_));
 sky130_fd_sc_hd__a311o_1 _15150_ (.A1(_11053_),
    .A2(_11068_),
    .A3(_07849_),
    .B1(_11061_),
    .C1(_10844_),
    .X(_07930_));
 sky130_fd_sc_hd__nand3_1 _15151_ (.A(_10839_),
    .B(_07764_),
    .C(_07835_),
    .Y(_07931_));
 sky130_fd_sc_hd__o21ai_0 _15152_ (.A1(_10839_),
    .A2(_07930_),
    .B1(_07931_),
    .Y(_07932_));
 sky130_fd_sc_hd__nor2_1 _15153_ (.A(_07845_),
    .B(_07928_),
    .Y(_07933_));
 sky130_fd_sc_hd__o21ai_0 _15154_ (.A1(_07831_),
    .A2(_07933_),
    .B1(_11115_),
    .Y(_07934_));
 sky130_fd_sc_hd__nor2_1 _15155_ (.A(_11068_),
    .B(_07770_),
    .Y(_07935_));
 sky130_fd_sc_hd__o21ai_0 _15156_ (.A1(_07843_),
    .A2(_07935_),
    .B1(_11095_),
    .Y(_07936_));
 sky130_fd_sc_hd__a21oi_1 _15157_ (.A1(_07934_),
    .A2(_07936_),
    .B1(_07820_),
    .Y(_07937_));
 sky130_fd_sc_hd__a21oi_1 _15158_ (.A1(_11095_),
    .A2(_07932_),
    .B1(_07937_),
    .Y(_07938_));
 sky130_fd_sc_hd__nor2_1 _15159_ (.A(_11061_),
    .B(_07928_),
    .Y(_07939_));
 sky130_fd_sc_hd__a31oi_1 _15160_ (.A1(_11053_),
    .A2(_11061_),
    .A3(_11095_),
    .B1(_07939_),
    .Y(_07940_));
 sky130_fd_sc_hd__o22ai_1 _15161_ (.A1(_11053_),
    .A2(_07928_),
    .B1(_07940_),
    .B2(_11067_),
    .Y(_07941_));
 sky130_fd_sc_hd__nand2_1 _15162_ (.A(_07771_),
    .B(_07941_),
    .Y(_07942_));
 sky130_fd_sc_hd__o211ai_1 _15163_ (.A1(_07928_),
    .A2(_07929_),
    .B1(_07938_),
    .C1(_07942_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[21] ));
 sky130_fd_sc_hd__nand2_1 _15164_ (.A(_11053_),
    .B(_11068_),
    .Y(_07943_));
 sky130_fd_sc_hd__nor2_1 _15165_ (.A(_10838_),
    .B(_07865_),
    .Y(_07944_));
 sky130_fd_sc_hd__a31oi_2 _15166_ (.A1(_10838_),
    .A2(_07809_),
    .A3(_07943_),
    .B1(_07944_),
    .Y(_07945_));
 sky130_fd_sc_hd__nand2_1 _15167_ (.A(_07874_),
    .B(_07921_),
    .Y(_07946_));
 sky130_fd_sc_hd__nand2_1 _15168_ (.A(_07945_),
    .B(_07946_),
    .Y(_07947_));
 sky130_fd_sc_hd__nor2_2 _15169_ (.A(_11059_),
    .B(_11067_),
    .Y(_07948_));
 sky130_fd_sc_hd__a22oi_1 _15170_ (.A1(_11067_),
    .A2(_11086_),
    .B1(_11099_),
    .B2(_07948_),
    .Y(_07949_));
 sky130_fd_sc_hd__o21ai_1 _15171_ (.A1(_11055_),
    .A2(_07949_),
    .B1(_07771_),
    .Y(_07950_));
 sky130_fd_sc_hd__nand2_1 _15172_ (.A(_11115_),
    .B(_07831_),
    .Y(_07951_));
 sky130_fd_sc_hd__o22ai_1 _15173_ (.A1(_07886_),
    .A2(_07950_),
    .B1(_07951_),
    .B2(_07820_),
    .Y(_07952_));
 sky130_fd_sc_hd__mux2i_1 _15174_ (.A0(_11084_),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[6] ),
    .S(net449),
    .Y(_07953_));
 sky130_fd_sc_hd__a31oi_1 _15175_ (.A1(_07806_),
    .A2(_07929_),
    .A3(_07950_),
    .B1(_07953_),
    .Y(_07954_));
 sky130_fd_sc_hd__a211o_1 _15176_ (.A1(\if_stage_i.compressed_decoder_i.instr_i[4] ),
    .A2(_07947_),
    .B1(_07952_),
    .C1(_07954_),
    .X(\if_stage_i.compressed_decoder_i.instr_o[22] ));
 sky130_fd_sc_hd__inv_1 _15177_ (.A(_11082_),
    .Y(_07955_));
 sky130_fd_sc_hd__nand2_1 _15178_ (.A(net449),
    .B(_11121_),
    .Y(_07956_));
 sky130_fd_sc_hd__o21ai_2 _15179_ (.A1(net449),
    .A2(_11101_),
    .B1(_07956_),
    .Y(_07957_));
 sky130_fd_sc_hd__a22oi_1 _15180_ (.A1(_07955_),
    .A2(_07778_),
    .B1(_07957_),
    .B2(_11068_),
    .Y(_07958_));
 sky130_fd_sc_hd__o221ai_1 _15181_ (.A1(_11074_),
    .A2(_07920_),
    .B1(_07958_),
    .B2(_11061_),
    .C1(_07771_),
    .Y(_07959_));
 sky130_fd_sc_hd__o21ai_0 _15182_ (.A1(_11055_),
    .A2(_07959_),
    .B1(_07957_),
    .Y(_07960_));
 sky130_fd_sc_hd__nand2_1 _15183_ (.A(_07929_),
    .B(_07959_),
    .Y(_07961_));
 sky130_fd_sc_hd__a21oi_1 _15184_ (.A1(_07919_),
    .A2(_07957_),
    .B1(_07801_),
    .Y(_07962_));
 sky130_fd_sc_hd__nand2_1 _15185_ (.A(_07802_),
    .B(_07962_),
    .Y(_07963_));
 sky130_fd_sc_hd__o21ai_0 _15186_ (.A1(_07935_),
    .A2(_07962_),
    .B1(_11082_),
    .Y(_07964_));
 sky130_fd_sc_hd__a31oi_1 _15187_ (.A1(_07951_),
    .A2(_07963_),
    .A3(_07964_),
    .B1(_07820_),
    .Y(_07965_));
 sky130_fd_sc_hd__a21oi_1 _15188_ (.A1(_07960_),
    .A2(_07961_),
    .B1(_07965_),
    .Y(_07966_));
 sky130_fd_sc_hd__o21ai_0 _15189_ (.A1(_07955_),
    .A2(_07945_),
    .B1(_07966_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[23] ));
 sky130_fd_sc_hd__mux2_2 _15190_ (.A0(_11105_),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[8] ),
    .S(net450),
    .X(_07967_));
 sky130_fd_sc_hd__nor2_2 _15191_ (.A(_11114_),
    .B(_07829_),
    .Y(_07968_));
 sky130_fd_sc_hd__a21oi_1 _15192_ (.A1(\if_stage_i.compressed_decoder_i.instr_i[6] ),
    .A2(_07829_),
    .B1(_07968_),
    .Y(_07969_));
 sky130_fd_sc_hd__nand3_1 _15193_ (.A(_11115_),
    .B(_07802_),
    .C(_07967_),
    .Y(_07970_));
 sky130_fd_sc_hd__o211ai_1 _15194_ (.A1(_11086_),
    .A2(_07802_),
    .B1(_07970_),
    .C1(_11068_),
    .Y(_07971_));
 sky130_fd_sc_hd__o21ai_0 _15195_ (.A1(_11068_),
    .A2(_11086_),
    .B1(_11061_),
    .Y(_07972_));
 sky130_fd_sc_hd__a32oi_1 _15196_ (.A1(_11053_),
    .A2(_07971_),
    .A3(_07972_),
    .B1(_11078_),
    .B2(_07819_),
    .Y(_07973_));
 sky130_fd_sc_hd__o21ai_1 _15197_ (.A1(_07828_),
    .A2(_07969_),
    .B1(_07973_),
    .Y(_07974_));
 sky130_fd_sc_hd__o211ai_1 _15198_ (.A1(_11061_),
    .A2(_11068_),
    .B1(_07799_),
    .C1(_07974_),
    .Y(_07975_));
 sky130_fd_sc_hd__o21ai_0 _15199_ (.A1(_11053_),
    .A2(_07967_),
    .B1(_07780_),
    .Y(_07976_));
 sky130_fd_sc_hd__nand2_1 _15200_ (.A(_07799_),
    .B(_07974_),
    .Y(_07977_));
 sky130_fd_sc_hd__a32oi_1 _15201_ (.A1(_11053_),
    .A2(_11086_),
    .A3(_07975_),
    .B1(_07976_),
    .B2(_07977_),
    .Y(_07978_));
 sky130_fd_sc_hd__a21oi_1 _15202_ (.A1(_07887_),
    .A2(_07967_),
    .B1(_07978_),
    .Y(_07979_));
 sky130_fd_sc_hd__a221oi_1 _15203_ (.A1(_11078_),
    .A2(_07778_),
    .B1(_07886_),
    .B2(_07967_),
    .C1(_07858_),
    .Y(_07980_));
 sky130_fd_sc_hd__a21oi_1 _15204_ (.A1(_07858_),
    .A2(_07979_),
    .B1(_07980_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[24] ));
 sky130_fd_sc_hd__nand2_1 _15205_ (.A(net450),
    .B(_11122_),
    .Y(_07981_));
 sky130_fd_sc_hd__o21ai_2 _15206_ (.A1(net451),
    .A2(_11109_),
    .B1(_07981_),
    .Y(_07982_));
 sky130_fd_sc_hd__nor2_1 _15207_ (.A(_10838_),
    .B(_07835_),
    .Y(_07983_));
 sky130_fd_sc_hd__a21oi_4 _15208_ (.A1(_07771_),
    .A2(_07886_),
    .B1(_07983_),
    .Y(_07984_));
 sky130_fd_sc_hd__nor2_1 _15209_ (.A(_07796_),
    .B(_07770_),
    .Y(_07985_));
 sky130_fd_sc_hd__a21oi_1 _15210_ (.A1(_07771_),
    .A2(_07863_),
    .B1(_07985_),
    .Y(_07986_));
 sky130_fd_sc_hd__nand3_1 _15211_ (.A(_11055_),
    .B(_11067_),
    .C(_07968_),
    .Y(_07987_));
 sky130_fd_sc_hd__a21oi_1 _15212_ (.A1(_07912_),
    .A2(_07987_),
    .B1(_11059_),
    .Y(_07988_));
 sky130_fd_sc_hd__nand2_1 _15213_ (.A(_11074_),
    .B(_07982_),
    .Y(_07989_));
 sky130_fd_sc_hd__a21oi_1 _15214_ (.A1(_07826_),
    .A2(_07989_),
    .B1(_07778_),
    .Y(_07990_));
 sky130_fd_sc_hd__nand2_1 _15215_ (.A(_11055_),
    .B(_11091_),
    .Y(_07991_));
 sky130_fd_sc_hd__nor2_1 _15216_ (.A(_11059_),
    .B(_07829_),
    .Y(_07992_));
 sky130_fd_sc_hd__o22ai_1 _15217_ (.A1(_11114_),
    .A2(_07990_),
    .B1(_07991_),
    .B2(_07992_),
    .Y(_07993_));
 sky130_fd_sc_hd__o21ai_0 _15218_ (.A1(_07988_),
    .A2(_07993_),
    .B1(_07799_),
    .Y(_07994_));
 sky130_fd_sc_hd__o221ai_2 _15219_ (.A1(_07982_),
    .A2(_07984_),
    .B1(_07986_),
    .B2(_11114_),
    .C1(_07994_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[25] ));
 sky130_fd_sc_hd__mux2_2 _15220_ (.A0(_11071_),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[10] ),
    .S(net450),
    .X(_07995_));
 sky130_fd_sc_hd__nand2_1 _15221_ (.A(_11115_),
    .B(_07826_),
    .Y(_07996_));
 sky130_fd_sc_hd__nor2_1 _15222_ (.A(_11073_),
    .B(_07995_),
    .Y(_07997_));
 sky130_fd_sc_hd__a21oi_1 _15223_ (.A1(_11082_),
    .A2(_07829_),
    .B1(_07968_),
    .Y(_07998_));
 sky130_fd_sc_hd__a21oi_1 _15224_ (.A1(_11061_),
    .A2(_11114_),
    .B1(_07776_),
    .Y(_07999_));
 sky130_fd_sc_hd__a221oi_1 _15225_ (.A1(_11103_),
    .A2(_07819_),
    .B1(_07948_),
    .B2(_11082_),
    .C1(_07999_),
    .Y(_08000_));
 sky130_fd_sc_hd__o221ai_1 _15226_ (.A1(_07996_),
    .A2(_07997_),
    .B1(_07998_),
    .B2(_07828_),
    .C1(_08000_),
    .Y(_08001_));
 sky130_fd_sc_hd__a21oi_2 _15227_ (.A1(_11114_),
    .A2(_07813_),
    .B1(_07755_),
    .Y(_08002_));
 sky130_fd_sc_hd__nand2_1 _15228_ (.A(_11068_),
    .B(_11103_),
    .Y(_08003_));
 sky130_fd_sc_hd__nand2_1 _15229_ (.A(_11067_),
    .B(_11091_),
    .Y(_08004_));
 sky130_fd_sc_hd__nand2_1 _15230_ (.A(_08003_),
    .B(_08004_),
    .Y(_08005_));
 sky130_fd_sc_hd__a222oi_1 _15231_ (.A1(_07983_),
    .A2(_07995_),
    .B1(_08001_),
    .B2(_08002_),
    .C1(_08005_),
    .C2(_07985_),
    .Y(_08006_));
 sky130_fd_sc_hd__nand2_1 _15232_ (.A(_11067_),
    .B(_11103_),
    .Y(_08007_));
 sky130_fd_sc_hd__nand2_1 _15233_ (.A(_11061_),
    .B(_11082_),
    .Y(_08008_));
 sky130_fd_sc_hd__o21ai_0 _15234_ (.A1(_11061_),
    .A2(_08007_),
    .B1(_08008_),
    .Y(_08009_));
 sky130_fd_sc_hd__a221oi_1 _15235_ (.A1(_07886_),
    .A2(_07995_),
    .B1(_08009_),
    .B2(_11053_),
    .C1(_07858_),
    .Y(_08010_));
 sky130_fd_sc_hd__a21oi_1 _15236_ (.A1(_07858_),
    .A2(_08006_),
    .B1(_08010_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[26] ));
 sky130_fd_sc_hd__a21oi_1 _15237_ (.A1(_07844_),
    .A2(_07893_),
    .B1(_11086_),
    .Y(_08011_));
 sky130_fd_sc_hd__nand2_1 _15238_ (.A(net450),
    .B(_11123_),
    .Y(_08012_));
 sky130_fd_sc_hd__o21ai_2 _15239_ (.A1(net450),
    .A2(_11076_),
    .B1(_08012_),
    .Y(_08013_));
 sky130_fd_sc_hd__a21oi_1 _15240_ (.A1(_11074_),
    .A2(_08013_),
    .B1(_07996_),
    .Y(_08014_));
 sky130_fd_sc_hd__a21oi_1 _15241_ (.A1(_11095_),
    .A2(_07829_),
    .B1(_07968_),
    .Y(_08015_));
 sky130_fd_sc_hd__nor2_1 _15242_ (.A(_07828_),
    .B(_08015_),
    .Y(_08016_));
 sky130_fd_sc_hd__o41ai_1 _15243_ (.A1(_07999_),
    .A2(_08011_),
    .A3(_08014_),
    .A4(_08016_),
    .B1(_08002_),
    .Y(_08017_));
 sky130_fd_sc_hd__nand2_1 _15244_ (.A(_11068_),
    .B(_11107_),
    .Y(_08018_));
 sky130_fd_sc_hd__nand2_1 _15245_ (.A(_11067_),
    .B(_11095_),
    .Y(_08019_));
 sky130_fd_sc_hd__nand2_1 _15246_ (.A(_08018_),
    .B(_08019_),
    .Y(_08020_));
 sky130_fd_sc_hd__o21ai_0 _15247_ (.A1(_07929_),
    .A2(_08013_),
    .B1(_07858_),
    .Y(_08021_));
 sky130_fd_sc_hd__a21oi_1 _15248_ (.A1(_07985_),
    .A2(_08020_),
    .B1(_08021_),
    .Y(_08022_));
 sky130_fd_sc_hd__nor2_1 _15249_ (.A(_07863_),
    .B(_08013_),
    .Y(_08023_));
 sky130_fd_sc_hd__a211oi_1 _15250_ (.A1(_11107_),
    .A2(_07813_),
    .B1(_07858_),
    .C1(_08023_),
    .Y(_08024_));
 sky130_fd_sc_hd__a21oi_2 _15251_ (.A1(_08017_),
    .A2(_08022_),
    .B1(_08024_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[27] ));
 sky130_fd_sc_hd__nand2_1 _15252_ (.A(net451),
    .B(_11124_),
    .Y(_08025_));
 sky130_fd_sc_hd__o21ai_2 _15253_ (.A1(net451),
    .A2(_11112_),
    .B1(_08025_),
    .Y(_08026_));
 sky130_fd_sc_hd__o21ai_0 _15254_ (.A1(_11061_),
    .A2(\if_stage_i.compressed_decoder_i.instr_i[9] ),
    .B1(_07764_),
    .Y(_08027_));
 sky130_fd_sc_hd__a221oi_1 _15255_ (.A1(_11061_),
    .A2(_11114_),
    .B1(_08027_),
    .B2(_11055_),
    .C1(_07768_),
    .Y(_08028_));
 sky130_fd_sc_hd__a21oi_1 _15256_ (.A1(_11074_),
    .A2(_08026_),
    .B1(_07996_),
    .Y(_08029_));
 sky130_fd_sc_hd__a21oi_1 _15257_ (.A1(\if_stage_i.compressed_decoder_i.instr_i[4] ),
    .A2(_07829_),
    .B1(_07968_),
    .Y(_08030_));
 sky130_fd_sc_hd__nor2_1 _15258_ (.A(_07828_),
    .B(_08030_),
    .Y(_08031_));
 sky130_fd_sc_hd__o31ai_1 _15259_ (.A1(_08028_),
    .A2(_08029_),
    .A3(_08031_),
    .B1(_08002_),
    .Y(_08032_));
 sky130_fd_sc_hd__o221ai_1 _15260_ (.A1(_07779_),
    .A2(_07889_),
    .B1(_07984_),
    .B2(_08026_),
    .C1(_08032_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[28] ));
 sky130_fd_sc_hd__mux2i_4 _15261_ (.A0(_11051_),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[13] ),
    .S(net451),
    .Y(_08033_));
 sky130_fd_sc_hd__a21oi_1 _15262_ (.A1(_11059_),
    .A2(_07776_),
    .B1(_11114_),
    .Y(_08034_));
 sky130_fd_sc_hd__a21oi_1 _15263_ (.A1(_11074_),
    .A2(_08033_),
    .B1(_07996_),
    .Y(_08035_));
 sky130_fd_sc_hd__a211oi_1 _15264_ (.A1(_11074_),
    .A2(_07819_),
    .B1(_08034_),
    .C1(_08035_),
    .Y(_08036_));
 sky130_fd_sc_hd__nand3_1 _15265_ (.A(_11074_),
    .B(_07813_),
    .C(_07771_),
    .Y(_08037_));
 sky130_fd_sc_hd__o221ai_2 _15266_ (.A1(_07984_),
    .A2(_08033_),
    .B1(_08036_),
    .B2(_07755_),
    .C1(_08037_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[29] ));
 sky130_fd_sc_hd__nand2_1 _15267_ (.A(_07806_),
    .B(_07888_),
    .Y(_08038_));
 sky130_fd_sc_hd__nand2_1 _15268_ (.A(_11115_),
    .B(_07775_),
    .Y(_08039_));
 sky130_fd_sc_hd__nand3_1 _15269_ (.A(_07760_),
    .B(_07768_),
    .C(_08039_),
    .Y(_08040_));
 sky130_fd_sc_hd__nand2_1 _15270_ (.A(_07780_),
    .B(_07779_),
    .Y(_08041_));
 sky130_fd_sc_hd__a21oi_2 _15271_ (.A1(_07991_),
    .A2(_08040_),
    .B1(_08041_),
    .Y(_08042_));
 sky130_fd_sc_hd__a221o_1 _15272_ (.A1(_07874_),
    .A2(_07879_),
    .B1(_08038_),
    .B2(_11091_),
    .C1(_08042_),
    .X(\if_stage_i.compressed_decoder_i.instr_o[2] ));
 sky130_fd_sc_hd__o21ai_1 _15273_ (.A1(_07858_),
    .A2(_07863_),
    .B1(_07929_),
    .Y(_08043_));
 sky130_fd_sc_hd__nor2_1 _15274_ (.A(net451),
    .B(_11057_),
    .Y(_08044_));
 sky130_fd_sc_hd__a21oi_2 _15275_ (.A1(net451),
    .A2(_11125_),
    .B1(_08044_),
    .Y(_08045_));
 sky130_fd_sc_hd__nand2_1 _15276_ (.A(_11074_),
    .B(_11115_),
    .Y(_08046_));
 sky130_fd_sc_hd__o22ai_1 _15277_ (.A1(_11115_),
    .A2(_07759_),
    .B1(_08045_),
    .B2(_08046_),
    .Y(_08047_));
 sky130_fd_sc_hd__a21oi_1 _15278_ (.A1(_11078_),
    .A2(_11115_),
    .B1(_11074_),
    .Y(_08048_));
 sky130_fd_sc_hd__a21oi_1 _15279_ (.A1(_11078_),
    .A2(_08047_),
    .B1(_08048_),
    .Y(_08049_));
 sky130_fd_sc_hd__o221ai_1 _15280_ (.A1(_11053_),
    .A2(_11107_),
    .B1(_07943_),
    .B2(_08049_),
    .C1(_11059_),
    .Y(_08050_));
 sky130_fd_sc_hd__o21ai_0 _15281_ (.A1(_11059_),
    .A2(_11114_),
    .B1(_08050_),
    .Y(_08051_));
 sky130_fd_sc_hd__a22o_1 _15282_ (.A1(_08043_),
    .A2(_08045_),
    .B1(_08051_),
    .B2(_08002_),
    .X(\if_stage_i.compressed_decoder_i.instr_o[30] ));
 sky130_fd_sc_hd__mux2i_4 _15283_ (.A0(_11065_),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[15] ),
    .S(net451),
    .Y(_08052_));
 sky130_fd_sc_hd__nand2_1 _15284_ (.A(_11074_),
    .B(_08052_),
    .Y(_08053_));
 sky130_fd_sc_hd__a21oi_1 _15285_ (.A1(_11078_),
    .A2(_08053_),
    .B1(_07801_),
    .Y(_08054_));
 sky130_fd_sc_hd__o32ai_2 _15286_ (.A1(_11114_),
    .A2(_07755_),
    .A3(_08054_),
    .B1(_08052_),
    .B2(_07984_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[31] ));
 sky130_fd_sc_hd__nor3_1 _15287_ (.A(_07801_),
    .B(_07804_),
    .C(_07820_),
    .Y(_08055_));
 sky130_fd_sc_hd__o21ai_0 _15288_ (.A1(_08043_),
    .A2(_08055_),
    .B1(_11095_),
    .Y(_08056_));
 sky130_fd_sc_hd__o21ai_2 _15289_ (.A1(_07755_),
    .A2(_07844_),
    .B1(_08056_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[3] ));
 sky130_fd_sc_hd__a21oi_1 _15290_ (.A1(_11099_),
    .A2(_07776_),
    .B1(_07855_),
    .Y(_08057_));
 sky130_fd_sc_hd__o21ai_0 _15291_ (.A1(\if_stage_i.compressed_decoder_i.instr_i[4] ),
    .A2(_07804_),
    .B1(_11059_),
    .Y(_08058_));
 sky130_fd_sc_hd__a211oi_1 _15292_ (.A1(_11068_),
    .A2(_08058_),
    .B1(_07819_),
    .C1(_07755_),
    .Y(_08059_));
 sky130_fd_sc_hd__a21oi_1 _15293_ (.A1(_10844_),
    .A2(_08057_),
    .B1(_08059_),
    .Y(_08060_));
 sky130_fd_sc_hd__a21oi_1 _15294_ (.A1(_07760_),
    .A2(_08039_),
    .B1(_07801_),
    .Y(_08061_));
 sky130_fd_sc_hd__nor2_1 _15295_ (.A(_08041_),
    .B(_08061_),
    .Y(_08062_));
 sky130_fd_sc_hd__nand2_1 _15296_ (.A(_11053_),
    .B(_08062_),
    .Y(_08063_));
 sky130_fd_sc_hd__o21ai_0 _15297_ (.A1(\if_stage_i.compressed_decoder_i.instr_i[0] ),
    .A2(_08062_),
    .B1(_11099_),
    .Y(_08064_));
 sky130_fd_sc_hd__a21oi_1 _15298_ (.A1(_08063_),
    .A2(_08064_),
    .B1(_08059_),
    .Y(_08065_));
 sky130_fd_sc_hd__a21oi_1 _15299_ (.A1(_10838_),
    .A2(_08060_),
    .B1(_08065_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[4] ));
 sky130_fd_sc_hd__o21ai_0 _15300_ (.A1(_11082_),
    .A2(_11114_),
    .B1(_07802_),
    .Y(_08066_));
 sky130_fd_sc_hd__a21oi_1 _15301_ (.A1(_11059_),
    .A2(_08066_),
    .B1(_11067_),
    .Y(_08067_));
 sky130_fd_sc_hd__o21ai_0 _15302_ (.A1(_07879_),
    .A2(_08067_),
    .B1(_07874_),
    .Y(_08068_));
 sky130_fd_sc_hd__o21ai_0 _15303_ (.A1(_11061_),
    .A2(_11082_),
    .B1(_10844_),
    .Y(_08069_));
 sky130_fd_sc_hd__a221o_1 _15304_ (.A1(_07955_),
    .A2(_07865_),
    .B1(_08069_),
    .B2(_10838_),
    .C1(_07810_),
    .X(_08070_));
 sky130_fd_sc_hd__nand2_1 _15305_ (.A(_08068_),
    .B(_08070_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[5] ));
 sky130_fd_sc_hd__a21oi_1 _15306_ (.A1(\if_stage_i.compressed_decoder_i.instr_i[6] ),
    .A2(_07919_),
    .B1(_11061_),
    .Y(_08071_));
 sky130_fd_sc_hd__o21ai_0 _15307_ (.A1(_11067_),
    .A2(_08071_),
    .B1(_07844_),
    .Y(_08072_));
 sky130_fd_sc_hd__nand2_1 _15308_ (.A(_07799_),
    .B(_08072_),
    .Y(_08073_));
 sky130_fd_sc_hd__o221ai_2 _15309_ (.A1(_11086_),
    .A2(_07984_),
    .B1(_08041_),
    .B2(_07797_),
    .C1(_08073_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[6] ));
 sky130_fd_sc_hd__a22oi_1 _15310_ (.A1(_11091_),
    .A2(_07778_),
    .B1(_07886_),
    .B2(_11103_),
    .Y(_08074_));
 sky130_fd_sc_hd__o211ai_1 _15311_ (.A1(_07760_),
    .A2(_07789_),
    .B1(_07764_),
    .C1(_07835_),
    .Y(_08075_));
 sky130_fd_sc_hd__a31oi_1 _15312_ (.A1(_11115_),
    .A2(_07781_),
    .A3(_07760_),
    .B1(_11067_),
    .Y(_08076_));
 sky130_fd_sc_hd__a21oi_1 _15313_ (.A1(_11053_),
    .A2(_11103_),
    .B1(_11067_),
    .Y(_08077_));
 sky130_fd_sc_hd__o221ai_1 _15314_ (.A1(_11114_),
    .A2(_07893_),
    .B1(_08077_),
    .B2(_11061_),
    .C1(_08007_),
    .Y(_08078_));
 sky130_fd_sc_hd__nand2_1 _15315_ (.A(_07799_),
    .B(_08078_),
    .Y(_08079_));
 sky130_fd_sc_hd__o31ai_2 _15316_ (.A1(_07796_),
    .A2(_07767_),
    .A3(_08076_),
    .B1(_08079_),
    .Y(_08080_));
 sky130_fd_sc_hd__a21oi_1 _15317_ (.A1(_10839_),
    .A2(_08075_),
    .B1(_08080_),
    .Y(_08081_));
 sky130_fd_sc_hd__a21oi_1 _15318_ (.A1(_07779_),
    .A2(_08080_),
    .B1(_11103_),
    .Y(_08082_));
 sky130_fd_sc_hd__o22ai_1 _15319_ (.A1(_07858_),
    .A2(_08074_),
    .B1(_08081_),
    .B2(_08082_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[7] ));
 sky130_fd_sc_hd__a22oi_1 _15320_ (.A1(_11061_),
    .A2(_11095_),
    .B1(_11107_),
    .B2(_07800_),
    .Y(_08083_));
 sky130_fd_sc_hd__nand3_1 _15321_ (.A(_11095_),
    .B(_07778_),
    .C(_07771_),
    .Y(_08084_));
 sky130_fd_sc_hd__a21oi_1 _15322_ (.A1(_10839_),
    .A2(_07760_),
    .B1(_11061_),
    .Y(_08085_));
 sky130_fd_sc_hd__a21oi_1 _15323_ (.A1(_11067_),
    .A2(_07844_),
    .B1(_10844_),
    .Y(_08086_));
 sky130_fd_sc_hd__o21ai_0 _15324_ (.A1(_07810_),
    .A2(_08086_),
    .B1(_10838_),
    .Y(_08087_));
 sky130_fd_sc_hd__o311ai_1 _15325_ (.A1(_11067_),
    .A2(_07865_),
    .A3(_08085_),
    .B1(_08087_),
    .C1(_11107_),
    .Y(_08088_));
 sky130_fd_sc_hd__o311ai_2 _15326_ (.A1(_11067_),
    .A2(_07755_),
    .A3(_08083_),
    .B1(_08084_),
    .C1(_08088_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[8] ));
 sky130_fd_sc_hd__o22ai_1 _15327_ (.A1(_11068_),
    .A2(_11099_),
    .B1(_07893_),
    .B2(_11086_),
    .Y(_08089_));
 sky130_fd_sc_hd__a31oi_1 _15328_ (.A1(_11053_),
    .A2(_07771_),
    .A3(_08089_),
    .B1(\if_stage_i.compressed_decoder_i.instr_i[9] ),
    .Y(_08090_));
 sky130_fd_sc_hd__a22oi_1 _15329_ (.A1(\if_stage_i.compressed_decoder_i.instr_i[9] ),
    .A2(_07800_),
    .B1(_07948_),
    .B2(\if_stage_i.compressed_decoder_i.instr_i[4] ),
    .Y(_08091_));
 sky130_fd_sc_hd__nor2_1 _15330_ (.A(_10844_),
    .B(_08091_),
    .Y(_08092_));
 sky130_fd_sc_hd__o22ai_1 _15331_ (.A1(\if_stage_i.compressed_decoder_i.instr_i[4] ),
    .A2(_07793_),
    .B1(_07893_),
    .B2(\if_stage_i.compressed_decoder_i.instr_i[6] ),
    .Y(_08093_));
 sky130_fd_sc_hd__a221oi_1 _15332_ (.A1(\if_stage_i.compressed_decoder_i.instr_i[0] ),
    .A2(_07764_),
    .B1(_08093_),
    .B2(_11053_),
    .C1(_08090_),
    .Y(_08094_));
 sky130_fd_sc_hd__o21ai_0 _15333_ (.A1(_08092_),
    .A2(_08094_),
    .B1(_10838_),
    .Y(_08095_));
 sky130_fd_sc_hd__o31ai_1 _15334_ (.A1(_10838_),
    .A2(_07807_),
    .A3(_08090_),
    .B1(_08095_),
    .Y(\if_stage_i.compressed_decoder_i.instr_o[9] ));
 sky130_fd_sc_hd__inv_1 _15335_ (.A(_07887_),
    .Y(\if_stage_i.compressed_decoder_i.is_compressed_o ));
 sky130_fd_sc_hd__nand3b_1 _15336_ (.A_N(_11162_),
    .B(\id_stage_i.controller_i.instr_valid_i ),
    .C(_11010_),
    .Y(_08096_));
 sky130_fd_sc_hd__nor2_1 _15337_ (.A(_11004_),
    .B(_08096_),
    .Y(_08097_));
 sky130_fd_sc_hd__nand2_1 _15338_ (.A(_11201_),
    .B(_08097_),
    .Y(_08098_));
 sky130_fd_sc_hd__o31ai_1 _15339_ (.A1(net1026),
    .A2(_11164_),
    .A3(_11201_),
    .B1(_08098_),
    .Y(\if_stage_i.instr_valid_id_d ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1199 ();
 sky130_fd_sc_hd__clkinv_16 _15341_ (.A(net444),
    .Y(_08100_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1196 ();
 sky130_fd_sc_hd__clkinvlp_4 _15345_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .Y(_08104_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1195 ();
 sky130_fd_sc_hd__nand2b_4 _15347_ (.A_N(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .B(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .Y(_08106_));
 sky130_fd_sc_hd__nor3_4 _15348_ (.A(_08104_),
    .B(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .C(_08106_),
    .Y(_08107_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1194 ();
 sky130_fd_sc_hd__nand3b_4 _15350_ (.A_N(\id_stage_i.controller_i.instr_fetch_err_i ),
    .B(_08107_),
    .C(\id_stage_i.controller_i.instr_valid_i ),
    .Y(_08109_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1193 ();
 sky130_fd_sc_hd__nor3_4 _15352_ (.A(\id_stage_i.controller_i.instr_i[30] ),
    .B(\id_stage_i.controller_i.instr_i[26] ),
    .C(net1033),
    .Y(_08111_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1188 ();
 sky130_fd_sc_hd__nor3_2 _15358_ (.A(net801),
    .B(net821),
    .C(net754),
    .Y(_08117_));
 sky130_fd_sc_hd__nand2_1 _15359_ (.A(_08111_),
    .B(_08117_),
    .Y(_08118_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1186 ();
 sky130_fd_sc_hd__nand2_1 _15362_ (.A(net575),
    .B(net801),
    .Y(_08121_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1185 ();
 sky130_fd_sc_hd__nand2_1 _15364_ (.A(\id_stage_i.controller_i.instr_i[30] ),
    .B(net754),
    .Y(_08123_));
 sky130_fd_sc_hd__or4_1 _15365_ (.A(net663),
    .B(net821),
    .C(_08121_),
    .D(_08123_),
    .X(_08124_));
 sky130_fd_sc_hd__nand2_1 _15366_ (.A(_08118_),
    .B(_08124_),
    .Y(_08125_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1173 ();
 sky130_fd_sc_hd__nor2b_1 _15379_ (.A(net545),
    .B_N(net811),
    .Y(_08138_));
 sky130_fd_sc_hd__nand2_1 _15380_ (.A(net670),
    .B(_08138_),
    .Y(_08139_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1171 ();
 sky130_fd_sc_hd__nand2b_4 _15383_ (.A_N(net382),
    .B(net372),
    .Y(_08142_));
 sky130_fd_sc_hd__nor3_4 _15384_ (.A(net552),
    .B(_08139_),
    .C(_08142_),
    .Y(_08143_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1163 ();
 sky130_fd_sc_hd__and2_4 _15393_ (.A(net810),
    .B(net343),
    .X(_08152_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1159 ();
 sky130_fd_sc_hd__nand2_1 _15398_ (.A(net1543),
    .B(_08138_),
    .Y(_08157_));
 sky130_fd_sc_hd__nor4_2 _15399_ (.A(net669),
    .B(net372),
    .C(_08118_),
    .D(_08157_),
    .Y(_08158_));
 sky130_fd_sc_hd__nor4_4 _15400_ (.A(net821),
    .B(net811),
    .C(net669),
    .D(net801),
    .Y(_08159_));
 sky130_fd_sc_hd__nand2_1 _15401_ (.A(net1302),
    .B(_08111_),
    .Y(_08160_));
 sky130_fd_sc_hd__clkinv_16 _15402_ (.A(net334),
    .Y(_08161_));
 sky130_fd_sc_hd__inv_4 _15403_ (.A(net336),
    .Y(_08162_));
 sky130_fd_sc_hd__nand2_8 _15404_ (.A(_08161_),
    .B(_08162_),
    .Y(_08163_));
 sky130_fd_sc_hd__nor4_4 _15405_ (.A(net372),
    .B(net552),
    .C(_08160_),
    .D(_08163_),
    .Y(_08164_));
 sky130_fd_sc_hd__a211oi_2 _15406_ (.A1(_08125_),
    .A2(_08143_),
    .B1(_08158_),
    .C1(_08164_),
    .Y(_08165_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1146 ();
 sky130_fd_sc_hd__nor2_8 _15420_ (.A(net385),
    .B(net390),
    .Y(_08179_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1139 ();
 sky130_fd_sc_hd__nor2_8 _15428_ (.A(net393),
    .B(net405),
    .Y(_08187_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1137 ();
 sky130_fd_sc_hd__nand3b_4 _15431_ (.A_N(net436),
    .B(_08179_),
    .C(net649),
    .Y(_08190_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1134 ();
 sky130_fd_sc_hd__or3_4 _15435_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .B(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .C(net448),
    .X(_08194_));
 sky130_fd_sc_hd__or4_2 _15436_ (.A(\id_stage_i.controller_i.instr_i[14] ),
    .B(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .C(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .D(_08194_),
    .X(_08195_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1130 ();
 sky130_fd_sc_hd__nor2_1 _15441_ (.A(net491),
    .B(net680),
    .Y(_08200_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1129 ();
 sky130_fd_sc_hd__nor4bb_4 _15443_ (.A(\id_stage_i.controller_i.instr_i[3] ),
    .B(\id_stage_i.controller_i.instr_i[2] ),
    .C_N(\id_stage_i.controller_i.instr_i[1] ),
    .D_N(\id_stage_i.controller_i.instr_i[0] ),
    .Y(_08202_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1127 ();
 sky130_fd_sc_hd__and2_2 _15446_ (.A(net1094),
    .B(\id_stage_i.controller_i.instr_i[5] ),
    .X(_08205_));
 sky130_fd_sc_hd__and3_4 _15447_ (.A(net1125),
    .B(net594),
    .C(_08205_),
    .X(_08206_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1126 ();
 sky130_fd_sc_hd__o311ai_4 _15449_ (.A1(_08165_),
    .A2(_08190_),
    .A3(_08195_),
    .B1(_08200_),
    .C1(_08206_),
    .Y(_08208_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1124 ();
 sky130_fd_sc_hd__nand2_1 _15452_ (.A(net491),
    .B(net681),
    .Y(_08211_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1123 ();
 sky130_fd_sc_hd__nor2_1 _15454_ (.A(net1099),
    .B(net1125),
    .Y(_08213_));
 sky130_fd_sc_hd__nand2_2 _15455_ (.A(net595),
    .B(_08213_),
    .Y(_08214_));
 sky130_fd_sc_hd__a21oi_1 _15456_ (.A1(_08100_),
    .A2(_08211_),
    .B1(_08214_),
    .Y(_08215_));
 sky130_fd_sc_hd__nor2b_4 _15457_ (.A(net1095),
    .B_N(net1124),
    .Y(_08216_));
 sky130_fd_sc_hd__nand2_4 _15458_ (.A(net599),
    .B(_08216_),
    .Y(_08217_));
 sky130_fd_sc_hd__nor2_1 _15459_ (.A(net813),
    .B(net673),
    .Y(_08218_));
 sky130_fd_sc_hd__nor2_1 _15460_ (.A(net803),
    .B(net825),
    .Y(_08219_));
 sky130_fd_sc_hd__nand2_1 _15461_ (.A(_08218_),
    .B(_08219_),
    .Y(_08220_));
 sky130_fd_sc_hd__nor2_1 _15462_ (.A(net576),
    .B(net664),
    .Y(_08221_));
 sky130_fd_sc_hd__nand2b_1 _15463_ (.A_N(net1089),
    .B(net917),
    .Y(_08222_));
 sky130_fd_sc_hd__nand2_1 _15464_ (.A(_08221_),
    .B(_08222_),
    .Y(_08223_));
 sky130_fd_sc_hd__nor2b_4 _15465_ (.A(net680),
    .B_N(net967),
    .Y(_08224_));
 sky130_fd_sc_hd__o21ai_0 _15466_ (.A1(_08220_),
    .A2(_08223_),
    .B1(_08224_),
    .Y(_08225_));
 sky130_fd_sc_hd__nor3_1 _15467_ (.A(net564),
    .B(_08217_),
    .C(_08225_),
    .Y(_08226_));
 sky130_fd_sc_hd__nand2_4 _15468_ (.A(\id_stage_i.controller_i.instr_i[1] ),
    .B(\id_stage_i.controller_i.instr_i[0] ),
    .Y(_08227_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1122 ();
 sky130_fd_sc_hd__and4b_2 _15470_ (.A_N(net1127),
    .B(\id_stage_i.controller_i.instr_i[2] ),
    .C(\id_stage_i.controller_i.instr_i[0] ),
    .D(\id_stage_i.controller_i.instr_i[1] ),
    .X(_08229_));
 sky130_fd_sc_hd__nor2_2 _15471_ (.A(net1096),
    .B(net995),
    .Y(_08230_));
 sky130_fd_sc_hd__or2_1 _15472_ (.A(net677),
    .B(net1086),
    .X(_08231_));
 sky130_fd_sc_hd__nand4_1 _15473_ (.A(net844),
    .B(_08229_),
    .C(_08230_),
    .D(_08231_),
    .Y(_08232_));
 sky130_fd_sc_hd__nor2b_2 _15474_ (.A(_08227_),
    .B_N(_08232_),
    .Y(_08233_));
 sky130_fd_sc_hd__inv_1 _15475_ (.A(\id_stage_i.controller_i.instr_i[3] ),
    .Y(_08234_));
 sky130_fd_sc_hd__or3_4 _15476_ (.A(net966),
    .B(net677),
    .C(net1086),
    .X(_08235_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1121 ();
 sky130_fd_sc_hd__and3b_2 _15478_ (.A_N(\id_stage_i.controller_i.instr_i[4] ),
    .B(net1000),
    .C(\id_stage_i.controller_i.instr_i[6] ),
    .X(_08237_));
 sky130_fd_sc_hd__a41oi_1 _15479_ (.A1(\id_stage_i.controller_i.instr_i[2] ),
    .A2(_08234_),
    .A3(_08235_),
    .A4(_08237_),
    .B1(\id_stage_i.decoder_i.illegal_c_insn_i ),
    .Y(_08238_));
 sky130_fd_sc_hd__clkinv_2 _15480_ (.A(\id_stage_i.controller_i.instr_i[2] ),
    .Y(_08239_));
 sky130_fd_sc_hd__nand2b_1 _15481_ (.A_N(net995),
    .B(net1094),
    .Y(_08240_));
 sky130_fd_sc_hd__a21oi_1 _15482_ (.A1(_08239_),
    .A2(_08240_),
    .B1(_08216_),
    .Y(_08241_));
 sky130_fd_sc_hd__nor3b_1 _15483_ (.A(net1094),
    .B(\id_stage_i.controller_i.instr_i[5] ),
    .C_N(\id_stage_i.controller_i.instr_i[3] ),
    .Y(_08242_));
 sky130_fd_sc_hd__nor2b_1 _15484_ (.A(net1124),
    .B_N(\id_stage_i.controller_i.instr_i[2] ),
    .Y(_08243_));
 sky130_fd_sc_hd__o21ai_2 _15485_ (.A1(_08205_),
    .A2(_08242_),
    .B1(_08243_),
    .Y(_08244_));
 sky130_fd_sc_hd__o21ai_0 _15486_ (.A1(net841),
    .A2(_08241_),
    .B1(_08244_),
    .Y(_08245_));
 sky130_fd_sc_hd__nor2_1 _15487_ (.A(net968),
    .B(net444),
    .Y(_08246_));
 sky130_fd_sc_hd__nand3b_1 _15488_ (.A_N(net444),
    .B(net564),
    .C(net1098),
    .Y(_08247_));
 sky130_fd_sc_hd__o31ai_1 _15489_ (.A1(net1097),
    .A2(net564),
    .A3(_08246_),
    .B1(_08247_),
    .Y(_08248_));
 sky130_fd_sc_hd__nand4bb_2 _15490_ (.A_N(\id_stage_i.controller_i.instr_i[2] ),
    .B_N(\id_stage_i.controller_i.instr_i[3] ),
    .C(\id_stage_i.controller_i.instr_i[1] ),
    .D(\id_stage_i.controller_i.instr_i[0] ),
    .Y(_08249_));
 sky130_fd_sc_hd__nor2_1 _15491_ (.A(net1127),
    .B(_08249_),
    .Y(_08250_));
 sky130_fd_sc_hd__nand3_1 _15492_ (.A(net679),
    .B(_08248_),
    .C(_08250_),
    .Y(_08251_));
 sky130_fd_sc_hd__nand4_1 _15493_ (.A(_08233_),
    .B(_08238_),
    .C(_08245_),
    .D(_08251_),
    .Y(_08252_));
 sky130_fd_sc_hd__a211oi_2 _15494_ (.A1(net564),
    .A2(_08215_),
    .B1(_08226_),
    .C1(_08252_),
    .Y(_08253_));
 sky130_fd_sc_hd__inv_2 _15495_ (.A(net973),
    .Y(_08254_));
 sky130_fd_sc_hd__nand2_1 _15496_ (.A(net1089),
    .B(net922),
    .Y(_08255_));
 sky130_fd_sc_hd__or3_1 _15497_ (.A(net445),
    .B(net1089),
    .C(net917),
    .X(_08256_));
 sky130_fd_sc_hd__a32oi_4 _15498_ (.A1(_08254_),
    .A2(_08255_),
    .A3(_08256_),
    .B1(_08224_),
    .B2(_08222_),
    .Y(_08257_));
 sky130_fd_sc_hd__nor4_4 _15499_ (.A(net802),
    .B(net672),
    .C(net812),
    .D(net664),
    .Y(_08258_));
 sky130_fd_sc_hd__a21oi_2 _15500_ (.A1(net445),
    .A2(net917),
    .B1(net823),
    .Y(_08259_));
 sky130_fd_sc_hd__nand3b_1 _15501_ (.A_N(net576),
    .B(_08258_),
    .C(_08259_),
    .Y(_08260_));
 sky130_fd_sc_hd__nor3_4 _15502_ (.A(net444),
    .B(net679),
    .C(net969),
    .Y(_08261_));
 sky130_fd_sc_hd__nor2_4 _15503_ (.A(net824),
    .B(net918),
    .Y(_08262_));
 sky130_fd_sc_hd__o211ai_2 _15504_ (.A1(net577),
    .A2(_08261_),
    .B1(net528),
    .C1(_08262_),
    .Y(_08263_));
 sky130_fd_sc_hd__o21ai_0 _15505_ (.A1(_08257_),
    .A2(_08260_),
    .B1(_08263_),
    .Y(_08264_));
 sky130_fd_sc_hd__nand3_4 _15506_ (.A(net996),
    .B(net597),
    .C(_08216_),
    .Y(_08265_));
 sky130_fd_sc_hd__nand4_2 _15507_ (.A(net970),
    .B(net680),
    .C(_08159_),
    .D(_08111_),
    .Y(_08266_));
 sky130_fd_sc_hd__or3b_1 _15508_ (.A(_08264_),
    .B(_08265_),
    .C_N(_08266_),
    .X(_08267_));
 sky130_fd_sc_hd__nand3_4 _15509_ (.A(_08208_),
    .B(_08253_),
    .C(_08267_),
    .Y(_08268_));
 sky130_fd_sc_hd__nor2_8 _15510_ (.A(_08268_),
    .B(_08109_),
    .Y(_08269_));
 sky130_fd_sc_hd__nor3b_2 _15511_ (.A(net802),
    .B(net664),
    .C_N(net578),
    .Y(_08270_));
 sky130_fd_sc_hd__nand3_4 _15512_ (.A(_08218_),
    .B(_08262_),
    .C(_08270_),
    .Y(_08271_));
 sky130_fd_sc_hd__nor2_8 _15513_ (.A(_08265_),
    .B(_08271_),
    .Y(_08272_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1117 ();
 sky130_fd_sc_hd__nand3_2 _15518_ (.A(_08100_),
    .B(net1524),
    .C(_08272_),
    .Y(_08277_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1115 ();
 sky130_fd_sc_hd__inv_8 _15521_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .Y(_08280_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1114 ();
 sky130_fd_sc_hd__nand2b_2 _15523_ (.A_N(net1097),
    .B(net1127),
    .Y(_08282_));
 sky130_fd_sc_hd__nand2_1 _15524_ (.A(net564),
    .B(net597),
    .Y(_08283_));
 sky130_fd_sc_hd__nor4_2 _15525_ (.A(net488),
    .B(_08282_),
    .C(_08283_),
    .D(_08271_),
    .Y(_08284_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1112 ();
 sky130_fd_sc_hd__nor2_1 _15528_ (.A(_08280_),
    .B(net316),
    .Y(_08287_));
 sky130_fd_sc_hd__nor2_1 _15529_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .B(_08287_),
    .Y(_08288_));
 sky130_fd_sc_hd__nand2_1 _15530_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .B(_08277_),
    .Y(_08289_));
 sky130_fd_sc_hd__o21ai_0 _15531_ (.A1(_08277_),
    .A2(_08288_),
    .B1(_08289_),
    .Y(_00000_));
 sky130_fd_sc_hd__or2_4 _15532_ (.A(_08265_),
    .B(_08271_),
    .X(_08290_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1111 ();
 sky130_fd_sc_hd__nor3_4 _15534_ (.A(_08280_),
    .B(net489),
    .C(_08290_),
    .Y(_08292_));
 sky130_fd_sc_hd__mux2_1 _15535_ (.A0(_08292_),
    .A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .S(_08277_),
    .X(_00001_));
 sky130_fd_sc_hd__or2_1 _15536_ (.A(net824),
    .B(net918),
    .X(_08293_));
 sky130_fd_sc_hd__nand2_8 _15537_ (.A(net579),
    .B(net529),
    .Y(_08294_));
 sky130_fd_sc_hd__or3_4 _15538_ (.A(_08293_),
    .B(_08294_),
    .C(_08265_),
    .X(_08295_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1109 ();
 sky130_fd_sc_hd__a22oi_2 _15541_ (.A1(net1124),
    .A2(_08230_),
    .B1(_08240_),
    .B2(_08239_),
    .Y(_08298_));
 sky130_fd_sc_hd__o21ai_4 _15542_ (.A1(_08298_),
    .A2(\id_stage_i.controller_i.instr_i[3] ),
    .B1(_08244_),
    .Y(_08299_));
 sky130_fd_sc_hd__a21oi_4 _15543_ (.A1(net1087),
    .A2(_08206_),
    .B1(_08227_),
    .Y(_08300_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1108 ();
 sky130_fd_sc_hd__nor2_4 _15545_ (.A(\load_store_unit_i.ls_fsm_cs[0] ),
    .B(\load_store_unit_i.ls_fsm_cs[1] ),
    .Y(_08302_));
 sky130_fd_sc_hd__nand2b_1 _15546_ (.A_N(\load_store_unit_i.handle_misaligned_q ),
    .B(\load_store_unit_i.ls_fsm_cs[0] ),
    .Y(_08303_));
 sky130_fd_sc_hd__nor2b_1 _15547_ (.A(\load_store_unit_i.ls_fsm_cs[2] ),
    .B_N(\load_store_unit_i.ls_fsm_cs[1] ),
    .Y(_08304_));
 sky130_fd_sc_hd__a22oi_4 _15548_ (.A1(\load_store_unit_i.ls_fsm_cs[2] ),
    .A2(_08302_),
    .B1(_08303_),
    .B2(_08304_),
    .Y(_08305_));
 sky130_fd_sc_hd__and2_2 _15549_ (.A(_08232_),
    .B(_08305_),
    .X(_08306_));
 sky130_fd_sc_hd__nand3_4 _15550_ (.A(_08299_),
    .B(_08306_),
    .C(_08300_),
    .Y(_08307_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1107 ();
 sky130_fd_sc_hd__clkinv_4 _15552_ (.A(net390),
    .Y(_08309_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1103 ();
 sky130_fd_sc_hd__mux4_1 _15557_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[135] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[167] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[199] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[231] ),
    .S0(net853),
    .S1(net403),
    .X(_08314_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1101 ();
 sky130_fd_sc_hd__nand2b_1 _15560_ (.A_N(_08314_),
    .B(net398),
    .Y(_08317_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1099 ();
 sky130_fd_sc_hd__mux2_1 _15563_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[71] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[103] ),
    .S(net439),
    .X(_08320_));
 sky130_fd_sc_hd__nor2b_4 _15564_ (.A(net413),
    .B_N(net438),
    .Y(_08321_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1098 ();
 sky130_fd_sc_hd__a221o_1 _15566_ (.A1(net1072),
    .A2(_08320_),
    .B1(net540),
    .B2(\gen_regfile_ff.register_file_i.rf_reg[39] ),
    .C1(net399),
    .X(_08323_));
 sky130_fd_sc_hd__and2_4 _15567_ (.A(net394),
    .B(net1225),
    .X(_08324_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1095 ();
 sky130_fd_sc_hd__mux4_2 _15571_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[391] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[423] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[455] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[487] ),
    .S0(net419),
    .S1(net412),
    .X(_08328_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1094 ();
 sky130_fd_sc_hd__mux4_1 _15573_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[263] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[295] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[327] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[359] ),
    .S0(net419),
    .S1(net1235),
    .X(_08330_));
 sky130_fd_sc_hd__nor2b_4 _15574_ (.A(net394),
    .B_N(net1152),
    .Y(_08331_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1093 ();
 sky130_fd_sc_hd__a22o_1 _15576_ (.A1(_08324_),
    .A2(_08328_),
    .B1(_08330_),
    .B2(net330),
    .X(_08333_));
 sky130_fd_sc_hd__a31o_1 _15577_ (.A1(_08309_),
    .A2(_08317_),
    .A3(_08323_),
    .B1(_08333_),
    .X(_08334_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1089 ();
 sky130_fd_sc_hd__mux4_1 _15582_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[519] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[551] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[583] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[615] ),
    .S0(net427),
    .S1(net1112),
    .X(_08339_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1087 ();
 sky130_fd_sc_hd__nor2_8 _15585_ (.A(net1225),
    .B(net394),
    .Y(_08342_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1086 ();
 sky130_fd_sc_hd__nor2b_4 _15587_ (.A(net1225),
    .B_N(net394),
    .Y(_08344_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1082 ();
 sky130_fd_sc_hd__mux4_1 _15592_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[647] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[679] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[711] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[743] ),
    .S0(net427),
    .S1(net1112),
    .X(_08349_));
 sky130_fd_sc_hd__a22oi_2 _15593_ (.A1(_08339_),
    .A2(_08342_),
    .B1(net608),
    .B2(_08349_),
    .Y(_08350_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1080 ();
 sky130_fd_sc_hd__mux4_2 _15596_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[775] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[807] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[839] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[871] ),
    .S0(net416),
    .S1(net1070),
    .X(_08353_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1078 ();
 sky130_fd_sc_hd__mux4_2 _15599_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[903] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[935] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[967] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[999] ),
    .S0(net419),
    .S1(net412),
    .X(_08356_));
 sky130_fd_sc_hd__a22oi_4 _15600_ (.A1(_08353_),
    .A2(net330),
    .B1(_08324_),
    .B2(_08356_),
    .Y(_08357_));
 sky130_fd_sc_hd__nand3_1 _15601_ (.A(net386),
    .B(_08350_),
    .C(_08357_),
    .Y(_08358_));
 sky130_fd_sc_hd__o21ai_4 _15602_ (.A1(_08334_),
    .A2(net386),
    .B1(_08358_),
    .Y(_08359_));
 sky130_fd_sc_hd__nor2_1 _15603_ (.A(_08359_),
    .B(_08307_),
    .Y(_08360_));
 sky130_fd_sc_hd__a21oi_1 _15604_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[7] ),
    .A2(_08307_),
    .B1(_08360_),
    .Y(_08361_));
 sky130_fd_sc_hd__nand2b_4 _15605_ (.A_N(\id_stage_i.id_fsm_q ),
    .B(\id_stage_i.controller_i.instr_valid_i ),
    .Y(_08362_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1077 ();
 sky130_fd_sc_hd__a32oi_4 _15607_ (.A1(net1580),
    .A2(net1128),
    .A3(_08230_),
    .B1(_08237_),
    .B2(_08362_),
    .Y(_08364_));
 sky130_fd_sc_hd__a21oi_2 _15608_ (.A1(_08230_),
    .A2(_08235_),
    .B1(_08205_),
    .Y(_08365_));
 sky130_fd_sc_hd__nand2_1 _15609_ (.A(net842),
    .B(_08229_),
    .Y(_08366_));
 sky130_fd_sc_hd__o32a_1 _15610_ (.A1(net842),
    .A2(_08227_),
    .A3(_08364_),
    .B1(_08365_),
    .B2(_08366_),
    .X(_08367_));
 sky130_fd_sc_hd__a22o_4 _15611_ (.A1(\load_store_unit_i.ls_fsm_cs[2] ),
    .A2(_08302_),
    .B1(_08303_),
    .B2(_08304_),
    .X(_08368_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1076 ();
 sky130_fd_sc_hd__a31oi_4 _15613_ (.A1(_08299_),
    .A2(_08367_),
    .A3(_08300_),
    .B1(_08368_),
    .Y(_08370_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1075 ();
 sky130_fd_sc_hd__and3_4 _15615_ (.A(_08299_),
    .B(_08300_),
    .C(_08306_),
    .X(_08372_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1074 ();
 sky130_fd_sc_hd__nand3_1 _15617_ (.A(\cs_registers_i.pc_id_i[7] ),
    .B(_08372_),
    .C(net941),
    .Y(_08374_));
 sky130_fd_sc_hd__o21ai_4 _15618_ (.A1(_08361_),
    .A2(net941),
    .B1(_08374_),
    .Y(_08375_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1073 ();
 sky130_fd_sc_hd__or2_4 _15620_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .X(_08377_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1072 ();
 sky130_fd_sc_hd__and3_1 _15622_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[39] ),
    .B(_08272_),
    .C(_08377_),
    .X(_08379_));
 sky130_fd_sc_hd__a21o_2 _15623_ (.A1(_08295_),
    .A2(_08375_),
    .B1(_08379_),
    .X(_08380_));
 sky130_fd_sc_hd__nor2b_4 _15624_ (.A(\id_stage_i.id_fsm_q ),
    .B_N(\id_stage_i.controller_i.instr_valid_i ),
    .Y(_08381_));
 sky130_fd_sc_hd__and3_2 _15625_ (.A(net598),
    .B(_08237_),
    .C(_08381_),
    .X(_08382_));
 sky130_fd_sc_hd__o21ai_0 _15626_ (.A1(_08205_),
    .A2(_08242_),
    .B1(\id_stage_i.controller_i.instr_i[2] ),
    .Y(_08383_));
 sky130_fd_sc_hd__nand3_1 _15627_ (.A(_08239_),
    .B(_08234_),
    .C(net1000),
    .Y(_08384_));
 sky130_fd_sc_hd__a21oi_2 _15628_ (.A1(_08383_),
    .A2(_08384_),
    .B1(net1124),
    .Y(_08385_));
 sky130_fd_sc_hd__nor3_2 _15629_ (.A(net840),
    .B(net1094),
    .C(_08243_),
    .Y(_08386_));
 sky130_fd_sc_hd__nor2b_2 _15630_ (.A(net1089),
    .B_N(net445),
    .Y(_08387_));
 sky130_fd_sc_hd__nand2_1 _15631_ (.A(net968),
    .B(net1088),
    .Y(_08388_));
 sky130_fd_sc_hd__nor3_1 _15632_ (.A(net680),
    .B(net1299),
    .C(_08388_),
    .Y(_08389_));
 sky130_fd_sc_hd__nor3_1 _15633_ (.A(net996),
    .B(_08249_),
    .C(_08282_),
    .Y(_08390_));
 sky130_fd_sc_hd__o21ai_2 _15634_ (.A1(_08387_),
    .A2(_08389_),
    .B1(_08390_),
    .Y(_08391_));
 sky130_fd_sc_hd__o211ai_4 _15635_ (.A1(_08385_),
    .A2(_08386_),
    .B1(_08391_),
    .C1(_08233_),
    .Y(_08392_));
 sky130_fd_sc_hd__nand2b_1 _15636_ (.A_N(net577),
    .B(_08258_),
    .Y(_08393_));
 sky130_fd_sc_hd__nor2b_1 _15637_ (.A(net968),
    .B_N(net445),
    .Y(_08394_));
 sky130_fd_sc_hd__nand4b_1 _15638_ (.A_N(_08393_),
    .B(_08100_),
    .C(_08262_),
    .D(_08394_),
    .Y(_08395_));
 sky130_fd_sc_hd__o221ai_4 _15639_ (.A1(_08257_),
    .A2(_08260_),
    .B1(_08266_),
    .B2(_08100_),
    .C1(_08263_),
    .Y(_08396_));
 sky130_fd_sc_hd__nor3b_1 _15640_ (.A(net445),
    .B(net1092),
    .C_N(net968),
    .Y(_08397_));
 sky130_fd_sc_hd__nor2b_1 _15641_ (.A(net972),
    .B_N(net1089),
    .Y(_08398_));
 sky130_fd_sc_hd__o21ai_2 _15642_ (.A1(_08397_),
    .A2(_08398_),
    .B1(_08262_),
    .Y(_08399_));
 sky130_fd_sc_hd__or2_0 _15643_ (.A(_08393_),
    .B(_08399_),
    .X(_08400_));
 sky130_fd_sc_hd__a31oi_2 _15644_ (.A1(_08395_),
    .A2(_08396_),
    .A3(_08400_),
    .B1(_08265_),
    .Y(_08401_));
 sky130_fd_sc_hd__nor2_1 _15645_ (.A(net680),
    .B(net1301),
    .Y(_08402_));
 sky130_fd_sc_hd__nor2_1 _15646_ (.A(_08388_),
    .B(_08402_),
    .Y(_08403_));
 sky130_fd_sc_hd__nor4_4 _15647_ (.A(net564),
    .B(_08246_),
    .C(_08217_),
    .D(_08403_),
    .Y(_08404_));
 sky130_fd_sc_hd__nor4_4 _15648_ (.A(_08401_),
    .B(_08392_),
    .C(_08382_),
    .D(_08404_),
    .Y(_08405_));
 sky130_fd_sc_hd__a21oi_2 _15649_ (.A1(_08395_),
    .A2(_08396_),
    .B1(_08265_),
    .Y(_08406_));
 sky130_fd_sc_hd__nand3_1 _15650_ (.A(net1089),
    .B(net1301),
    .C(_08111_),
    .Y(_08407_));
 sky130_fd_sc_hd__a211oi_2 _15651_ (.A1(net998),
    .A2(_08407_),
    .B1(_08211_),
    .C1(_08217_),
    .Y(_08408_));
 sky130_fd_sc_hd__and2_2 _15652_ (.A(net597),
    .B(_08237_),
    .X(_08409_));
 sky130_fd_sc_hd__nand2_4 _15653_ (.A(_08381_),
    .B(_08409_),
    .Y(_08410_));
 sky130_fd_sc_hd__xnor2_1 _15654_ (.A(net971),
    .B(net1089),
    .Y(_08411_));
 sky130_fd_sc_hd__nor2_1 _15655_ (.A(net445),
    .B(_08411_),
    .Y(_08412_));
 sky130_fd_sc_hd__nor2_1 _15656_ (.A(_08410_),
    .B(_08412_),
    .Y(_08413_));
 sky130_fd_sc_hd__nor4_4 _15657_ (.A(_08413_),
    .B(_08392_),
    .C(_08408_),
    .D(_08406_),
    .Y(_08414_));
 sky130_fd_sc_hd__nor2_1 _15658_ (.A(net831),
    .B(_08393_),
    .Y(_08415_));
 sky130_fd_sc_hd__nand2b_4 _15659_ (.A_N(\id_stage_i.controller_i.instr_i[13] ),
    .B(net967),
    .Y(_08416_));
 sky130_fd_sc_hd__mux2_1 _15660_ (.A0(_08222_),
    .A1(net922),
    .S(net445),
    .X(_08417_));
 sky130_fd_sc_hd__o32ai_1 _15661_ (.A1(_08100_),
    .A2(net923),
    .A3(_08416_),
    .B1(_08417_),
    .B2(net491),
    .Y(_08418_));
 sky130_fd_sc_hd__inv_1 _15662_ (.A(net917),
    .Y(_08419_));
 sky130_fd_sc_hd__a41oi_1 _15663_ (.A1(net1090),
    .A2(_08419_),
    .A3(net1298),
    .A4(_08224_),
    .B1(_08394_),
    .Y(_08420_));
 sky130_fd_sc_hd__nor2_1 _15664_ (.A(net564),
    .B(_08420_),
    .Y(_08421_));
 sky130_fd_sc_hd__a31oi_2 _15665_ (.A1(net564),
    .A2(_08415_),
    .A3(_08418_),
    .B1(_08421_),
    .Y(_08422_));
 sky130_fd_sc_hd__a211oi_4 _15666_ (.A1(net491),
    .A2(_08100_),
    .B1(_08410_),
    .C1(net445),
    .Y(_08423_));
 sky130_fd_sc_hd__o21bai_4 _15667_ (.A1(_08422_),
    .A2(_08217_),
    .B1_N(_08423_),
    .Y(_08424_));
 sky130_fd_sc_hd__nor2_1 _15668_ (.A(net997),
    .B(_08235_),
    .Y(_08425_));
 sky130_fd_sc_hd__a2111oi_2 _15669_ (.A1(net564),
    .A2(_08223_),
    .B1(_08217_),
    .C1(_08425_),
    .D1(_08220_),
    .Y(_08426_));
 sky130_fd_sc_hd__o21a_1 _15670_ (.A1(_08390_),
    .A2(_08382_),
    .B1(_08100_),
    .X(_08427_));
 sky130_fd_sc_hd__o21ai_4 _15671_ (.A1(_08426_),
    .A2(_08427_),
    .B1(_08224_),
    .Y(_08428_));
 sky130_fd_sc_hd__or3_4 _15672_ (.A(_08406_),
    .B(_08382_),
    .C(_08392_),
    .X(_08429_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1071 ();
 sky130_fd_sc_hd__a41oi_4 _15674_ (.A1(_08405_),
    .A2(_08414_),
    .A3(_08424_),
    .A4(_08428_),
    .B1(_08429_),
    .Y(_08431_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1070 ();
 sky130_fd_sc_hd__o21ai_1 _15676_ (.A1(net1126),
    .A2(_08362_),
    .B1(net1100),
    .Y(_08433_));
 sky130_fd_sc_hd__nand2_1 _15677_ (.A(_08100_),
    .B(_08213_),
    .Y(_08434_));
 sky130_fd_sc_hd__nand4_4 _15678_ (.A(net999),
    .B(net596),
    .C(_08433_),
    .D(_08434_),
    .Y(_08435_));
 sky130_fd_sc_hd__or2_4 _15679_ (.A(_08368_),
    .B(_08435_),
    .X(_08436_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1069 ();
 sky130_fd_sc_hd__nor4_2 _15681_ (.A(_08239_),
    .B(net845),
    .C(_08227_),
    .D(_08282_),
    .Y(_08438_));
 sky130_fd_sc_hd__a211o_4 _15682_ (.A1(_08362_),
    .A2(_08409_),
    .B1(_08438_),
    .C1(_08368_),
    .X(_08439_));
 sky130_fd_sc_hd__nand2_2 _15683_ (.A(_08205_),
    .B(_08229_),
    .Y(_08440_));
 sky130_fd_sc_hd__nor2_1 _15684_ (.A(net847),
    .B(_08362_),
    .Y(_08441_));
 sky130_fd_sc_hd__nor3_2 _15685_ (.A(net1099),
    .B(net995),
    .C(net444),
    .Y(_08442_));
 sky130_fd_sc_hd__nand4_4 _15686_ (.A(net844),
    .B(_08229_),
    .C(_08224_),
    .D(_08442_),
    .Y(_08443_));
 sky130_fd_sc_hd__o211ai_4 _15687_ (.A1(_08440_),
    .A2(_08441_),
    .B1(_08305_),
    .C1(_08443_),
    .Y(_08444_));
 sky130_fd_sc_hd__or4_2 _15688_ (.A(_08239_),
    .B(net844),
    .C(_08227_),
    .D(_08282_),
    .X(_08445_));
 sky130_fd_sc_hd__nand3_2 _15689_ (.A(_08205_),
    .B(_08229_),
    .C(_08362_),
    .Y(_08446_));
 sky130_fd_sc_hd__nand4_2 _15690_ (.A(net996),
    .B(_08100_),
    .C(net594),
    .D(_08213_),
    .Y(_08447_));
 sky130_fd_sc_hd__nand4_2 _15691_ (.A(_08445_),
    .B(_08443_),
    .C(_08446_),
    .D(_08447_),
    .Y(_08448_));
 sky130_fd_sc_hd__o22ai_4 _15692_ (.A1(_08439_),
    .A2(_08444_),
    .B1(_08448_),
    .B2(_08368_),
    .Y(_08449_));
 sky130_fd_sc_hd__and2_4 _15693_ (.A(_08436_),
    .B(_08449_),
    .X(_08450_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1067 ();
 sky130_fd_sc_hd__nor2b_4 _15696_ (.A(net338),
    .B_N(net377),
    .Y(_08453_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1065 ();
 sky130_fd_sc_hd__mux2i_1 _15699_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[551] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[615] ),
    .S(net355),
    .Y(_08456_));
 sky130_fd_sc_hd__nor2b_4 _15700_ (.A(net376),
    .B_N(net339),
    .Y(_08457_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1063 ();
 sky130_fd_sc_hd__mux2i_1 _15703_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[647] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[711] ),
    .S(net355),
    .Y(_08460_));
 sky130_fd_sc_hd__a22oi_1 _15704_ (.A1(net891),
    .A2(_08456_),
    .B1(net590),
    .B2(_08460_),
    .Y(_08461_));
 sky130_fd_sc_hd__nor2_8 _15705_ (.A(net337),
    .B(_08161_),
    .Y(_08462_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1062 ();
 sky130_fd_sc_hd__nor2_8 _15707_ (.A(net377),
    .B(net338),
    .Y(_08464_));
 sky130_fd_sc_hd__mux2i_1 _15708_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[519] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[583] ),
    .S(net355),
    .Y(_08465_));
 sky130_fd_sc_hd__mux2i_1 _15709_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[679] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[743] ),
    .S(net355),
    .Y(_08466_));
 sky130_fd_sc_hd__a22oi_1 _15710_ (.A1(net1047),
    .A2(_08465_),
    .B1(_08466_),
    .B2(net1024),
    .Y(_08467_));
 sky130_fd_sc_hd__nand3_2 _15711_ (.A(_08461_),
    .B(_08462_),
    .C(_08467_),
    .Y(_08468_));
 sky130_fd_sc_hd__nand4b_4 _15712_ (.A_N(net332),
    .B(net335),
    .C(net376),
    .D(net339),
    .Y(_08469_));
 sky130_fd_sc_hd__mux2i_1 _15713_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[423] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[487] ),
    .S(net369),
    .Y(_08470_));
 sky130_fd_sc_hd__nand4b_4 _15714_ (.A_N(net339),
    .B(net335),
    .C(net376),
    .D(net332),
    .Y(_08471_));
 sky130_fd_sc_hd__mux2i_1 _15715_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[807] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[871] ),
    .S(net370),
    .Y(_08472_));
 sky130_fd_sc_hd__o22ai_2 _15716_ (.A1(net868),
    .A2(_08470_),
    .B1(net523),
    .B2(_08472_),
    .Y(_08473_));
 sky130_fd_sc_hd__nand4bb_4 _15717_ (.A_N(net376),
    .B_N(net332),
    .C(net339),
    .D(net335),
    .Y(_08474_));
 sky130_fd_sc_hd__mux2i_1 _15718_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[391] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[455] ),
    .S(net369),
    .Y(_08475_));
 sky130_fd_sc_hd__nand4bb_4 _15719_ (.A_N(net376),
    .B_N(net338),
    .C(net335),
    .D(net333),
    .Y(_08476_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1061 ();
 sky130_fd_sc_hd__mux2i_1 _15721_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[775] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[839] ),
    .S(net369),
    .Y(_08478_));
 sky130_fd_sc_hd__o22ai_2 _15722_ (.A1(net895),
    .A2(_08475_),
    .B1(net502),
    .B2(_08478_),
    .Y(_08479_));
 sky130_fd_sc_hd__nor2_4 _15723_ (.A(_08473_),
    .B(_08479_),
    .Y(_08480_));
 sky130_fd_sc_hd__clkinv_16 _15724_ (.A(net338),
    .Y(_08481_));
 sky130_fd_sc_hd__mux4_1 _15725_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[135] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[167] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[199] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[231] ),
    .S0(net381),
    .S1(net366),
    .X(_08482_));
 sky130_fd_sc_hd__nor2_1 _15726_ (.A(_08481_),
    .B(_08482_),
    .Y(_08483_));
 sky130_fd_sc_hd__nor2b_4 _15727_ (.A(net381),
    .B_N(net366),
    .Y(_08484_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1060 ();
 sky130_fd_sc_hd__mux2_1 _15729_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[39] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[103] ),
    .S(net356),
    .X(_08486_));
 sky130_fd_sc_hd__a221oi_1 _15730_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[71] ),
    .A2(net324),
    .B1(_08486_),
    .B2(net378),
    .C1(net342),
    .Y(_08487_));
 sky130_fd_sc_hd__mux4_4 _15731_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[903] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[935] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[967] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[999] ),
    .S0(net379),
    .S1(net371),
    .X(_08488_));
 sky130_fd_sc_hd__and2_0 _15732_ (.A(net334),
    .B(net339),
    .X(_08489_));
 sky130_fd_sc_hd__mux4_1 _15733_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[263] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[295] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[327] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[359] ),
    .S0(net379),
    .S1(net371),
    .X(_08490_));
 sky130_fd_sc_hd__nor2_4 _15734_ (.A(net333),
    .B(net339),
    .Y(_08491_));
 sky130_fd_sc_hd__a22oi_2 _15735_ (.A1(_08488_),
    .A2(_08489_),
    .B1(_08490_),
    .B2(_08491_),
    .Y(_08492_));
 sky130_fd_sc_hd__o32a_2 _15736_ (.A1(_08163_),
    .A2(_08483_),
    .A3(_08487_),
    .B1(_08492_),
    .B2(_08162_),
    .X(_08493_));
 sky130_fd_sc_hd__nand3_4 _15737_ (.A(_08468_),
    .B(_08480_),
    .C(_08493_),
    .Y(_08494_));
 sky130_fd_sc_hd__nor2_8 _15738_ (.A(_08368_),
    .B(_08435_),
    .Y(_08495_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1059 ();
 sky130_fd_sc_hd__a22oi_4 _15740_ (.A1(net804),
    .A2(_08450_),
    .B1(_08495_),
    .B2(_08494_),
    .Y(_08497_));
 sky130_fd_sc_hd__xnor2_1 _15741_ (.A(net696),
    .B(_08497_),
    .Y(_08498_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1058 ();
 sky130_fd_sc_hd__inv_6 _15743_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .Y(_08500_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1057 ();
 sky130_fd_sc_hd__clkinv_16 _15745_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .Y(_08502_));
 sky130_fd_sc_hd__nor2_8 _15746_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .Y(_08503_));
 sky130_fd_sc_hd__nand3_4 _15747_ (.A(_08500_),
    .B(_08502_),
    .C(_08503_),
    .Y(_08504_));
 sky130_fd_sc_hd__nor2_1 _15748_ (.A(_08494_),
    .B(_08504_),
    .Y(_08505_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1056 ();
 sky130_fd_sc_hd__o22ai_1 _15750_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[39] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[7] ),
    .B2(_08503_),
    .Y(_08507_));
 sky130_fd_sc_hd__a2111oi_1 _15751_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(net767),
    .B1(_08505_),
    .C1(_08507_),
    .D1(_08295_),
    .Y(_08508_));
 sky130_fd_sc_hd__a21oi_2 _15752_ (.A1(_08290_),
    .A2(_08498_),
    .B1(_08508_),
    .Y(_08509_));
 sky130_fd_sc_hd__xnor2_4 _15753_ (.A(_08380_),
    .B(_08509_),
    .Y(_08510_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1055 ();
 sky130_fd_sc_hd__clkinv_16 _15755_ (.A(\gen_regfile_ff.register_file_i.raddr_a_i[4] ),
    .Y(_08512_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1053 ();
 sky130_fd_sc_hd__mux4_2 _15758_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[646] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[678] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[710] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[742] ),
    .S0(net417),
    .S1(net404),
    .X(_08515_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1051 ();
 sky130_fd_sc_hd__mux4_4 _15761_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[902] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[934] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[966] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[998] ),
    .S0(net416),
    .S1(net1235),
    .X(_08518_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1050 ();
 sky130_fd_sc_hd__a22oi_4 _15763_ (.A1(net609),
    .A2(_08515_),
    .B1(_08518_),
    .B2(net1227),
    .Y(_08520_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1049 ();
 sky130_fd_sc_hd__mux4_1 _15765_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[518] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[550] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[582] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[614] ),
    .S0(net418),
    .S1(net404),
    .X(_08522_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1048 ();
 sky130_fd_sc_hd__mux4_2 _15767_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[774] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[806] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[838] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[870] ),
    .S0(net416),
    .S1(net1113),
    .X(_08524_));
 sky130_fd_sc_hd__a22oi_4 _15768_ (.A1(_08342_),
    .A2(_08522_),
    .B1(_08524_),
    .B2(net330),
    .Y(_08525_));
 sky130_fd_sc_hd__nand2_2 _15769_ (.A(_08520_),
    .B(_08525_),
    .Y(_08526_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1046 ();
 sky130_fd_sc_hd__clkinv_16 _15772_ (.A(net394),
    .Y(_08529_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1045 ();
 sky130_fd_sc_hd__mux4_2 _15774_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[134] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[166] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[198] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[230] ),
    .S0(net853),
    .S1(net415),
    .X(_08531_));
 sky130_fd_sc_hd__nor2_1 _15775_ (.A(_08529_),
    .B(_08531_),
    .Y(_08532_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1044 ();
 sky130_fd_sc_hd__mux2_1 _15777_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[70] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[102] ),
    .S(net1130),
    .X(_08534_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1043 ();
 sky130_fd_sc_hd__a221oi_4 _15779_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[38] ),
    .A2(net542),
    .B1(_08534_),
    .B2(net413),
    .C1(net400),
    .Y(_08536_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1041 ();
 sky130_fd_sc_hd__mux4_2 _15782_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[390] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[422] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[454] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[486] ),
    .S0(net416),
    .S1(net1113),
    .X(_08539_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1040 ();
 sky130_fd_sc_hd__mux4_1 _15784_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[262] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[294] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[326] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[358] ),
    .S0(net416),
    .S1(net1070),
    .X(_08541_));
 sky130_fd_sc_hd__a22oi_4 _15785_ (.A1(net1226),
    .A2(_08539_),
    .B1(_08541_),
    .B2(net531),
    .Y(_08542_));
 sky130_fd_sc_hd__o311ai_2 _15786_ (.A1(net977),
    .A2(_08532_),
    .A3(_08536_),
    .B1(_08542_),
    .C1(_08512_),
    .Y(_08543_));
 sky130_fd_sc_hd__o21ai_4 _15787_ (.A1(_08512_),
    .A2(_08526_),
    .B1(_08543_),
    .Y(_08544_));
 sky130_fd_sc_hd__inv_1 _15788_ (.A(\cs_registers_i.pc_id_i[6] ),
    .Y(_08545_));
 sky130_fd_sc_hd__mux2i_1 _15789_ (.A0(net1285),
    .A1(_08545_),
    .S(net942),
    .Y(_08546_));
 sky130_fd_sc_hd__a22o_4 _15790_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[6] ),
    .A2(_08368_),
    .B1(_08372_),
    .B2(_08546_),
    .X(_08547_));
 sky130_fd_sc_hd__nand2_1 _15791_ (.A(_08295_),
    .B(_08547_),
    .Y(_08548_));
 sky130_fd_sc_hd__nand3_1 _15792_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[38] ),
    .B(_08272_),
    .C(_08377_),
    .Y(_08549_));
 sky130_fd_sc_hd__nand2_2 _15793_ (.A(_08548_),
    .B(_08549_),
    .Y(_08550_));
 sky130_fd_sc_hd__inv_1 _15794_ (.A(_08550_),
    .Y(_08551_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1038 ();
 sky130_fd_sc_hd__mux4_1 _15797_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[644] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[676] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[708] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[740] ),
    .S0(net418),
    .S1(net409),
    .X(_08554_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1036 ();
 sky130_fd_sc_hd__mux4_1 _15800_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[900] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[932] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[964] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[996] ),
    .S0(net418),
    .S1(net409),
    .X(_08557_));
 sky130_fd_sc_hd__a22oi_4 _15801_ (.A1(net612),
    .A2(_08554_),
    .B1(_08557_),
    .B2(net565),
    .Y(_08558_));
 sky130_fd_sc_hd__mux4_1 _15802_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[516] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[548] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[580] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[612] ),
    .S0(net418),
    .S1(net409),
    .X(_08559_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1035 ();
 sky130_fd_sc_hd__mux4_2 _15804_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[772] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[804] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[836] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[868] ),
    .S0(net418),
    .S1(net404),
    .X(_08561_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1034 ();
 sky130_fd_sc_hd__a22oi_4 _15806_ (.A1(_08342_),
    .A2(_08559_),
    .B1(_08561_),
    .B2(net330),
    .Y(_08563_));
 sky130_fd_sc_hd__nand2_1 _15807_ (.A(_08558_),
    .B(_08563_),
    .Y(_08564_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1033 ();
 sky130_fd_sc_hd__mux4_4 _15809_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[132] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[164] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[196] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[228] ),
    .S0(net440),
    .S1(net415),
    .X(_08566_));
 sky130_fd_sc_hd__nor2_2 _15810_ (.A(_08529_),
    .B(_08566_),
    .Y(_08567_));
 sky130_fd_sc_hd__mux2_1 _15811_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[68] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[100] ),
    .S(net989),
    .X(_08568_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1032 ();
 sky130_fd_sc_hd__a221oi_4 _15813_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[36] ),
    .A2(net542),
    .B1(_08568_),
    .B2(net1072),
    .C1(net399),
    .Y(_08570_));
 sky130_fd_sc_hd__mux4_1 _15814_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[388] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[420] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[452] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[484] ),
    .S0(net1109),
    .S1(net404),
    .X(_08571_));
 sky130_fd_sc_hd__mux4_1 _15815_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[260] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[292] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[324] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[356] ),
    .S0(net1109),
    .S1(net404),
    .X(_08572_));
 sky130_fd_sc_hd__a22oi_4 _15816_ (.A1(net1227),
    .A2(_08571_),
    .B1(_08572_),
    .B2(net330),
    .Y(_08573_));
 sky130_fd_sc_hd__o311ai_4 _15817_ (.A1(net978),
    .A2(_08567_),
    .A3(_08570_),
    .B1(_08573_),
    .C1(_08512_),
    .Y(_08574_));
 sky130_fd_sc_hd__o21ai_4 _15818_ (.A1(_08564_),
    .A2(_08512_),
    .B1(_08574_),
    .Y(_08575_));
 sky130_fd_sc_hd__o32ai_4 _15819_ (.A1(net843),
    .A2(_08227_),
    .A3(_08364_),
    .B1(_08365_),
    .B2(_08366_),
    .Y(_08576_));
 sky130_fd_sc_hd__nor2_2 _15820_ (.A(_08307_),
    .B(_08576_),
    .Y(_08577_));
 sky130_fd_sc_hd__nand2_1 _15821_ (.A(_08306_),
    .B(_08576_),
    .Y(_08578_));
 sky130_fd_sc_hd__o211a_1 _15822_ (.A1(_08306_),
    .A2(_08367_),
    .B1(_08299_),
    .C1(_08300_),
    .X(_08579_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1031 ();
 sky130_fd_sc_hd__nand2_8 _15824_ (.A(_08206_),
    .B(_08235_),
    .Y(_08581_));
 sky130_fd_sc_hd__nor2_1 _15825_ (.A(_08512_),
    .B(_08581_),
    .Y(_08582_));
 sky130_fd_sc_hd__o22ai_1 _15826_ (.A1(\cs_registers_i.pc_id_i[4] ),
    .A2(_08578_),
    .B1(_08579_),
    .B2(_08582_),
    .Y(_08583_));
 sky130_fd_sc_hd__nor2_1 _15827_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[4] ),
    .B(_08305_),
    .Y(_08584_));
 sky130_fd_sc_hd__a221o_4 _15828_ (.A1(net1455),
    .A2(_08577_),
    .B1(_08583_),
    .B2(_08305_),
    .C1(_08584_),
    .X(_08585_));
 sky130_fd_sc_hd__nor3_4 _15829_ (.A(_08293_),
    .B(_08294_),
    .C(_08265_),
    .Y(_08586_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1030 ();
 sky130_fd_sc_hd__nand3_1 _15831_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[36] ),
    .B(net1106),
    .C(_08377_),
    .Y(_08588_));
 sky130_fd_sc_hd__o21ai_2 _15832_ (.A1(_08272_),
    .A2(_08585_),
    .B1(_08588_),
    .Y(_08589_));
 sky130_fd_sc_hd__nor4bb_4 _15833_ (.A(net387),
    .B(net395),
    .C_N(net384),
    .D_N(net407),
    .Y(_08590_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1029 ();
 sky130_fd_sc_hd__mux2i_1 _15835_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[579] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[611] ),
    .S(net1008),
    .Y(_08592_));
 sky130_fd_sc_hd__and4b_4 _15836_ (.A_N(net384),
    .B(net387),
    .C(net395),
    .D(net1185),
    .X(_08593_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1028 ();
 sky130_fd_sc_hd__mux2i_1 _15838_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[451] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[483] ),
    .S(net938),
    .Y(_08595_));
 sky130_fd_sc_hd__a22oi_2 _15839_ (.A1(net535),
    .A2(_08592_),
    .B1(_08593_),
    .B2(_08595_),
    .Y(_08596_));
 sky130_fd_sc_hd__nor4b_4 _15840_ (.A(net384),
    .B(net395),
    .C(net1185),
    .D_N(net387),
    .Y(_08597_));
 sky130_fd_sc_hd__mux2i_1 _15841_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[259] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[291] ),
    .S(net422),
    .Y(_08598_));
 sky130_fd_sc_hd__nor4b_4 _15842_ (.A(net407),
    .B(net395),
    .C(net1082),
    .D_N(net384),
    .Y(_08599_));
 sky130_fd_sc_hd__mux2i_1 _15843_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[515] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[547] ),
    .S(net1008),
    .Y(_08600_));
 sky130_fd_sc_hd__a22oi_2 _15844_ (.A1(net1003),
    .A2(_08598_),
    .B1(net862),
    .B2(_08600_),
    .Y(_08601_));
 sky130_fd_sc_hd__and4b_4 _15845_ (.A_N(net387),
    .B(net395),
    .C(net1185),
    .D(net384),
    .X(_08602_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1026 ();
 sky130_fd_sc_hd__mux2i_1 _15848_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[707] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[739] ),
    .S(net422),
    .Y(_08605_));
 sky130_fd_sc_hd__nor4bb_4 _15849_ (.A(net387),
    .B(net407),
    .C_N(net395),
    .D_N(net384),
    .Y(_08606_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1025 ();
 sky130_fd_sc_hd__mux2i_1 _15851_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[643] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[675] ),
    .S(net1008),
    .Y(_08608_));
 sky130_fd_sc_hd__a22oi_2 _15852_ (.A1(_08602_),
    .A2(_08605_),
    .B1(net757),
    .B2(_08608_),
    .Y(_08609_));
 sky130_fd_sc_hd__nor4bb_4 _15853_ (.A(net384),
    .B(net395),
    .C_N(net387),
    .D_N(net407),
    .Y(_08610_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1024 ();
 sky130_fd_sc_hd__mux2i_1 _15855_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[323] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[355] ),
    .S(net422),
    .Y(_08612_));
 sky130_fd_sc_hd__nor4bb_4 _15856_ (.A(net384),
    .B(net407),
    .C_N(net395),
    .D_N(net387),
    .Y(_08613_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1023 ();
 sky130_fd_sc_hd__mux2i_1 _15858_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[387] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[419] ),
    .S(net1008),
    .Y(_08615_));
 sky130_fd_sc_hd__a22oi_2 _15859_ (.A1(net549),
    .A2(_08612_),
    .B1(net570),
    .B2(_08615_),
    .Y(_08616_));
 sky130_fd_sc_hd__nand4_4 _15860_ (.A(_08596_),
    .B(_08601_),
    .C(_08609_),
    .D(_08616_),
    .Y(_08617_));
 sky130_fd_sc_hd__nor2_8 _15861_ (.A(_08512_),
    .B(_08309_),
    .Y(_08618_));
 sky130_fd_sc_hd__mux4_1 _15862_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[771] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[803] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[835] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[867] ),
    .S0(net1311),
    .S1(net406),
    .X(_08619_));
 sky130_fd_sc_hd__nand2_1 _15863_ (.A(_08529_),
    .B(_08619_),
    .Y(_08620_));
 sky130_fd_sc_hd__mux4_1 _15864_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[899] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[931] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[963] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[995] ),
    .S0(net1311),
    .S1(net406),
    .X(_08621_));
 sky130_fd_sc_hd__nand2_1 _15865_ (.A(net393),
    .B(_08621_),
    .Y(_08622_));
 sky130_fd_sc_hd__mux2i_1 _15866_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[195] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[227] ),
    .S(net436),
    .Y(_08623_));
 sky130_fd_sc_hd__mux2i_1 _15867_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[131] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[163] ),
    .S(net436),
    .Y(_08624_));
 sky130_fd_sc_hd__mux2i_1 _15868_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[67] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[99] ),
    .S(net436),
    .Y(_08625_));
 sky130_fd_sc_hd__nand2_1 _15869_ (.A(net436),
    .B(\gen_regfile_ff.register_file_i.rf_reg[35] ),
    .Y(_08626_));
 sky130_fd_sc_hd__clkinv_4 _15870_ (.A(net786),
    .Y(_08627_));
 sky130_fd_sc_hd__mux4_2 _15871_ (.A0(_08623_),
    .A1(_08624_),
    .A2(_08625_),
    .A3(_08626_),
    .S0(_08627_),
    .S1(_08529_),
    .X(_08628_));
 sky130_fd_sc_hd__a32o_2 _15872_ (.A1(_08618_),
    .A2(_08620_),
    .A3(_08622_),
    .B1(_08628_),
    .B2(_08179_),
    .X(_08629_));
 sky130_fd_sc_hd__or2_4 _15873_ (.A(_08629_),
    .B(_08617_),
    .X(_08630_));
 sky130_fd_sc_hd__nor2_1 _15874_ (.A(\cs_registers_i.pc_id_i[3] ),
    .B(_08578_),
    .Y(_08631_));
 sky130_fd_sc_hd__and2_4 _15875_ (.A(_08206_),
    .B(_08235_),
    .X(_08632_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1022 ();
 sky130_fd_sc_hd__a21oi_1 _15877_ (.A1(net587),
    .A2(_08632_),
    .B1(_08579_),
    .Y(_08634_));
 sky130_fd_sc_hd__a2111oi_4 _15878_ (.A1(_08577_),
    .A2(_08630_),
    .B1(_08631_),
    .C1(_08634_),
    .D1(_08368_),
    .Y(_08635_));
 sky130_fd_sc_hd__a21oi_4 _15879_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[3] ),
    .A2(_08368_),
    .B1(_08635_),
    .Y(_08636_));
 sky130_fd_sc_hd__a21oi_1 _15880_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[35] ),
    .A2(_08377_),
    .B1(_08295_),
    .Y(_08637_));
 sky130_fd_sc_hd__a21oi_2 _15881_ (.A1(_08636_),
    .A2(_08295_),
    .B1(_08637_),
    .Y(_08638_));
 sky130_fd_sc_hd__nand2_4 _15882_ (.A(_08305_),
    .B(_08435_),
    .Y(_08639_));
 sky130_fd_sc_hd__o211a_4 _15883_ (.A1(_08440_),
    .A2(_08441_),
    .B1(_08305_),
    .C1(_08443_),
    .X(_08640_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1021 ();
 sky130_fd_sc_hd__a211oi_2 _15885_ (.A1(_08362_),
    .A2(_08409_),
    .B1(_08438_),
    .C1(_08368_),
    .Y(_08642_));
 sky130_fd_sc_hd__a41oi_4 _15886_ (.A1(_08445_),
    .A2(_08443_),
    .A3(_08446_),
    .A4(_08447_),
    .B1(_08368_),
    .Y(_08643_));
 sky130_fd_sc_hd__xnor2_2 _15887_ (.A(_08642_),
    .B(_08643_),
    .Y(_08644_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1020 ();
 sky130_fd_sc_hd__nor2_2 _15889_ (.A(_08439_),
    .B(_08643_),
    .Y(_08646_));
 sky130_fd_sc_hd__a32oi_4 _15890_ (.A1(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .A2(_08640_),
    .A3(_08644_),
    .B1(_08646_),
    .B2(net548),
    .Y(_08647_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1012 ();
 sky130_fd_sc_hd__mux4_1 _15899_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[291] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[355] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[419] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[483] ),
    .S0(net359),
    .S1(net340),
    .X(_08656_));
 sky130_fd_sc_hd__nand2_1 _15900_ (.A(net373),
    .B(_08656_),
    .Y(_08657_));
 sky130_fd_sc_hd__inv_12 _15901_ (.A(net1029),
    .Y(_08658_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1011 ();
 sky130_fd_sc_hd__mux4_1 _15903_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[259] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[323] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[387] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[451] ),
    .S0(net359),
    .S1(net340),
    .X(_08660_));
 sky130_fd_sc_hd__nand2_1 _15904_ (.A(_08658_),
    .B(_08660_),
    .Y(_08661_));
 sky130_fd_sc_hd__nand3_4 _15905_ (.A(net336),
    .B(_08657_),
    .C(_08661_),
    .Y(_08662_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1008 ();
 sky130_fd_sc_hd__mux2_1 _15909_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[67] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[195] ),
    .S(net341),
    .X(_08666_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1006 ();
 sky130_fd_sc_hd__nor2b_4 _15912_ (.A(net356),
    .B_N(net342),
    .Y(_08669_));
 sky130_fd_sc_hd__a22oi_2 _15913_ (.A1(net1077),
    .A2(_08666_),
    .B1(_08669_),
    .B2(\gen_regfile_ff.register_file_i.rf_reg[131] ),
    .Y(_08670_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1004 ();
 sky130_fd_sc_hd__mux2_1 _15916_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[35] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[99] ),
    .S(net365),
    .X(_08673_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1003 ();
 sky130_fd_sc_hd__mux2_1 _15918_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[163] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[227] ),
    .S(net365),
    .X(_08675_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1002 ();
 sky130_fd_sc_hd__a221oi_2 _15920_ (.A1(net328),
    .A2(_08673_),
    .B1(_08675_),
    .B2(net1153),
    .C1(net336),
    .Y(_08677_));
 sky130_fd_sc_hd__o21ai_4 _15921_ (.A1(net373),
    .A2(_08670_),
    .B1(_08677_),
    .Y(_08678_));
 sky130_fd_sc_hd__nand2b_4 _15922_ (.A_N(net335),
    .B(net333),
    .Y(_08679_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_999 ();
 sky130_fd_sc_hd__mux4_1 _15926_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[547] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[611] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[675] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[739] ),
    .S0(net352),
    .S1(net340),
    .X(_08683_));
 sky130_fd_sc_hd__mux4_1 _15927_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[515] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[579] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[643] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[707] ),
    .S0(net352),
    .S1(net340),
    .X(_08684_));
 sky130_fd_sc_hd__mux2i_4 _15928_ (.A0(_08683_),
    .A1(_08684_),
    .S(_08658_),
    .Y(_08685_));
 sky130_fd_sc_hd__mux4_1 _15929_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[771] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[803] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[835] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[867] ),
    .S0(net1310),
    .S1(net364),
    .X(_08686_));
 sky130_fd_sc_hd__and3b_4 _15930_ (.A_N(net339),
    .B(net337),
    .C(net332),
    .X(_08687_));
 sky130_fd_sc_hd__and3_4 _15931_ (.A(net333),
    .B(net335),
    .C(net342),
    .X(_08688_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_998 ();
 sky130_fd_sc_hd__mux4_1 _15933_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[899] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[931] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[963] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[995] ),
    .S0(net1310),
    .S1(net364),
    .X(_08690_));
 sky130_fd_sc_hd__a22oi_4 _15934_ (.A1(_08686_),
    .A2(_08687_),
    .B1(_08688_),
    .B2(_08690_),
    .Y(_08691_));
 sky130_fd_sc_hd__o21ai_1 _15935_ (.A1(_08679_),
    .A2(_08685_),
    .B1(_08691_),
    .Y(_08692_));
 sky130_fd_sc_hd__a31oi_4 _15936_ (.A1(_08662_),
    .A2(_08161_),
    .A3(_08678_),
    .B1(_08692_),
    .Y(_08693_));
 sky130_fd_sc_hd__o22ai_4 _15937_ (.A1(_08639_),
    .A2(_08647_),
    .B1(_08436_),
    .B2(_08693_),
    .Y(_08694_));
 sky130_fd_sc_hd__xor2_1 _15938_ (.A(net694),
    .B(_08694_),
    .X(_08695_));
 sky130_fd_sc_hd__nor3_4 _15939_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .C(_08377_),
    .Y(_08696_));
 sky130_fd_sc_hd__o22ai_1 _15940_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[35] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[3] ),
    .B2(_08503_),
    .Y(_08697_));
 sky130_fd_sc_hd__a221o_1 _15941_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(_08630_),
    .B1(_08693_),
    .B2(_08696_),
    .C1(_08697_),
    .X(_08698_));
 sky130_fd_sc_hd__nor2_1 _15942_ (.A(_08295_),
    .B(_08698_),
    .Y(_08699_));
 sky130_fd_sc_hd__a21oi_1 _15943_ (.A1(_08290_),
    .A2(_08695_),
    .B1(_08699_),
    .Y(_08700_));
 sky130_fd_sc_hd__or2_4 _15944_ (.A(_08638_),
    .B(_08700_),
    .X(_08701_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_997 ();
 sky130_fd_sc_hd__a32oi_4 _15946_ (.A1(net448),
    .A2(_08640_),
    .A3(_08644_),
    .B1(_08646_),
    .B2(net755),
    .Y(_08703_));
 sky130_fd_sc_hd__mux2i_1 _15947_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[804] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[868] ),
    .S(net345),
    .Y(_08704_));
 sky130_fd_sc_hd__nand2_4 _15948_ (.A(net377),
    .B(net338),
    .Y(_08705_));
 sky130_fd_sc_hd__nor2b_1 _15949_ (.A(net346),
    .B_N(\gen_regfile_ff.register_file_i.rf_reg[932] ),
    .Y(_08706_));
 sky130_fd_sc_hd__a211oi_1 _15950_ (.A1(net346),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[996] ),
    .B1(_08705_),
    .C1(_08706_),
    .Y(_08707_));
 sky130_fd_sc_hd__nand2_8 _15951_ (.A(net332),
    .B(net337),
    .Y(_08708_));
 sky130_fd_sc_hd__mux2i_1 _15952_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[900] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[964] ),
    .S(net346),
    .Y(_08709_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_996 ();
 sky130_fd_sc_hd__mux2i_1 _15954_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[772] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[836] ),
    .S(net345),
    .Y(_08711_));
 sky130_fd_sc_hd__a22o_1 _15955_ (.A1(net327),
    .A2(_08709_),
    .B1(_08711_),
    .B2(net1043),
    .X(_08712_));
 sky130_fd_sc_hd__a2111oi_4 _15956_ (.A1(_08453_),
    .A2(_08704_),
    .B1(_08707_),
    .C1(_08708_),
    .D1(_08712_),
    .Y(_08713_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_994 ();
 sky130_fd_sc_hd__mux2i_1 _15959_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[516] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[580] ),
    .S(net346),
    .Y(_08716_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_993 ();
 sky130_fd_sc_hd__mux2i_1 _15961_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[548] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[612] ),
    .S(net346),
    .Y(_08718_));
 sky130_fd_sc_hd__a22oi_1 _15962_ (.A1(net1046),
    .A2(_08716_),
    .B1(_08718_),
    .B2(_08453_),
    .Y(_08719_));
 sky130_fd_sc_hd__mux2i_1 _15963_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[676] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[740] ),
    .S(net345),
    .Y(_08720_));
 sky130_fd_sc_hd__mux2i_1 _15964_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[644] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[708] ),
    .S(net345),
    .Y(_08721_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_992 ();
 sky130_fd_sc_hd__a22oi_1 _15966_ (.A1(_08152_),
    .A2(_08720_),
    .B1(_08721_),
    .B2(net327),
    .Y(_08723_));
 sky130_fd_sc_hd__and3_1 _15967_ (.A(_08462_),
    .B(_08719_),
    .C(_08723_),
    .X(_08724_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_991 ();
 sky130_fd_sc_hd__mux2_1 _15969_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[36] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[100] ),
    .S(net367),
    .X(_08726_));
 sky130_fd_sc_hd__a221oi_2 _15970_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[68] ),
    .A2(_08484_),
    .B1(_08726_),
    .B2(net380),
    .C1(net343),
    .Y(_08727_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_989 ();
 sky130_fd_sc_hd__mux4_1 _15973_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[132] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[164] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[196] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[228] ),
    .S0(net379),
    .S1(net511),
    .X(_08730_));
 sky130_fd_sc_hd__nor2_8 _15974_ (.A(net334),
    .B(net337),
    .Y(_08731_));
 sky130_fd_sc_hd__o21ai_2 _15975_ (.A1(_08481_),
    .A2(_08730_),
    .B1(_08731_),
    .Y(_08732_));
 sky130_fd_sc_hd__nor2_4 _15976_ (.A(_08727_),
    .B(_08732_),
    .Y(_08733_));
 sky130_fd_sc_hd__nor2b_4 _15977_ (.A(net333),
    .B_N(net335),
    .Y(_08734_));
 sky130_fd_sc_hd__mux2i_1 _15978_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[388] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[452] ),
    .S(net345),
    .Y(_08735_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_988 ();
 sky130_fd_sc_hd__mux2i_1 _15980_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[260] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[324] ),
    .S(net345),
    .Y(_08737_));
 sky130_fd_sc_hd__a22oi_1 _15981_ (.A1(net327),
    .A2(_08735_),
    .B1(_08737_),
    .B2(net1043),
    .Y(_08738_));
 sky130_fd_sc_hd__mux2i_1 _15982_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[292] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[356] ),
    .S(net345),
    .Y(_08739_));
 sky130_fd_sc_hd__mux2i_1 _15983_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[420] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[484] ),
    .S(net345),
    .Y(_08740_));
 sky130_fd_sc_hd__a22oi_1 _15984_ (.A1(_08453_),
    .A2(_08739_),
    .B1(_08740_),
    .B2(_08152_),
    .Y(_08741_));
 sky130_fd_sc_hd__and3_1 _15985_ (.A(net706),
    .B(_08738_),
    .C(_08741_),
    .X(_08742_));
 sky130_fd_sc_hd__nor4_4 _15986_ (.A(_08713_),
    .B(_08742_),
    .C(_08733_),
    .D(_08724_),
    .Y(_08743_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_987 ();
 sky130_fd_sc_hd__o22a_4 _15988_ (.A1(_08639_),
    .A2(_08703_),
    .B1(net308),
    .B2(_08436_),
    .X(_08745_));
 sky130_fd_sc_hd__xnor2_2 _15989_ (.A(net695),
    .B(_08745_),
    .Y(_08746_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_986 ();
 sky130_fd_sc_hd__nand2_1 _15991_ (.A(_08696_),
    .B(net308),
    .Y(_08748_));
 sky130_fd_sc_hd__o221ai_1 _15992_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[36] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[4] ),
    .B2(_08503_),
    .C1(_08748_),
    .Y(_08749_));
 sky130_fd_sc_hd__a211oi_2 _15993_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(net1456),
    .B1(_08749_),
    .C1(_08290_),
    .Y(_08750_));
 sky130_fd_sc_hd__a21oi_2 _15994_ (.A1(net1134),
    .A2(_08746_),
    .B1(_08750_),
    .Y(_08751_));
 sky130_fd_sc_hd__maj3_2 _15995_ (.A(_08751_),
    .B(_08589_),
    .C(_08701_),
    .X(_08752_));
 sky130_fd_sc_hd__nand2b_1 _15996_ (.A_N(_08643_),
    .B(net551),
    .Y(_08753_));
 sky130_fd_sc_hd__nand3b_1 _15997_ (.A_N(\id_stage_i.controller_i.instr_is_compressed_i ),
    .B(_08444_),
    .C(_08643_),
    .Y(_08754_));
 sky130_fd_sc_hd__a21oi_2 _15998_ (.A1(_08753_),
    .A2(_08754_),
    .B1(_08439_),
    .Y(_08755_));
 sky130_fd_sc_hd__and3_1 _15999_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .B(_08640_),
    .C(_08644_),
    .X(_08756_));
 sky130_fd_sc_hd__mux2i_1 _16000_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[770] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[834] ),
    .S(net360),
    .Y(_08757_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_985 ();
 sky130_fd_sc_hd__mux2i_1 _16002_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[898] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[962] ),
    .S(net360),
    .Y(_08759_));
 sky130_fd_sc_hd__a221oi_2 _16003_ (.A1(net325),
    .A2(_08757_),
    .B1(_08759_),
    .B2(net1119),
    .C1(_08708_),
    .Y(_08760_));
 sky130_fd_sc_hd__mux4_1 _16004_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[802] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[866] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[930] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[994] ),
    .S0(net360),
    .S1(net340),
    .X(_08761_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_984 ();
 sky130_fd_sc_hd__nand2b_1 _16006_ (.A_N(_08761_),
    .B(net373),
    .Y(_08763_));
 sky130_fd_sc_hd__nand2_2 _16007_ (.A(_08760_),
    .B(_08763_),
    .Y(_08764_));
 sky130_fd_sc_hd__mux2_1 _16008_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[66] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[194] ),
    .S(net340),
    .X(_08765_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_981 ();
 sky130_fd_sc_hd__a221oi_1 _16012_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[130] ),
    .A2(_08669_),
    .B1(_08765_),
    .B2(net1141),
    .C1(net1154),
    .Y(_08769_));
 sky130_fd_sc_hd__mux4_1 _16013_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[34] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[98] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[162] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[226] ),
    .S0(net363),
    .S1(net340),
    .X(_08770_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_980 ();
 sky130_fd_sc_hd__o21ai_0 _16015_ (.A1(_08658_),
    .A2(_08770_),
    .B1(_08731_),
    .Y(_08772_));
 sky130_fd_sc_hd__nor2_2 _16016_ (.A(_08769_),
    .B(_08772_),
    .Y(_08773_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_978 ();
 sky130_fd_sc_hd__mux2i_1 _16019_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[514] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[578] ),
    .S(net350),
    .Y(_08776_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_977 ();
 sky130_fd_sc_hd__mux2i_1 _16021_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[546] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[610] ),
    .S(net350),
    .Y(_08778_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_976 ();
 sky130_fd_sc_hd__a22oi_1 _16023_ (.A1(net325),
    .A2(_08776_),
    .B1(_08778_),
    .B2(net329),
    .Y(_08780_));
 sky130_fd_sc_hd__mux2i_1 _16024_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[642] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[706] ),
    .S(net350),
    .Y(_08781_));
 sky130_fd_sc_hd__mux2i_1 _16025_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[674] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[738] ),
    .S(net350),
    .Y(_08782_));
 sky130_fd_sc_hd__a22oi_1 _16026_ (.A1(net1474),
    .A2(_08781_),
    .B1(_08782_),
    .B2(net1024),
    .Y(_08783_));
 sky130_fd_sc_hd__and3_4 _16027_ (.A(_08462_),
    .B(_08780_),
    .C(_08783_),
    .X(_08784_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_974 ();
 sky130_fd_sc_hd__mux2i_1 _16030_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[386] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[450] ),
    .S(net351),
    .Y(_08787_));
 sky130_fd_sc_hd__mux2i_1 _16031_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[258] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[322] ),
    .S(net351),
    .Y(_08788_));
 sky130_fd_sc_hd__a22oi_1 _16032_ (.A1(net1474),
    .A2(_08787_),
    .B1(_08788_),
    .B2(net325),
    .Y(_08789_));
 sky130_fd_sc_hd__mux2i_1 _16033_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[290] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[354] ),
    .S(net351),
    .Y(_08790_));
 sky130_fd_sc_hd__mux2i_1 _16034_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[418] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[482] ),
    .S(net351),
    .Y(_08791_));
 sky130_fd_sc_hd__a22oi_1 _16035_ (.A1(net329),
    .A2(_08790_),
    .B1(_08791_),
    .B2(net1024),
    .Y(_08792_));
 sky130_fd_sc_hd__and3_2 _16036_ (.A(net704),
    .B(_08789_),
    .C(_08792_),
    .X(_08793_));
 sky130_fd_sc_hd__nor3_4 _16037_ (.A(_08773_),
    .B(_08784_),
    .C(_08793_),
    .Y(_08794_));
 sky130_fd_sc_hd__nand2_8 _16038_ (.A(_08764_),
    .B(_08794_),
    .Y(_08795_));
 sky130_fd_sc_hd__o32ai_4 _16039_ (.A1(_08639_),
    .A2(_08755_),
    .A3(_08756_),
    .B1(_08436_),
    .B2(_08795_),
    .Y(_08796_));
 sky130_fd_sc_hd__xnor2_1 _16040_ (.A(net296),
    .B(_08796_),
    .Y(_08797_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_973 ();
 sky130_fd_sc_hd__nor2b_4 _16042_ (.A(net405),
    .B_N(net393),
    .Y(_08799_));
 sky130_fd_sc_hd__mux2i_1 _16043_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[898] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[930] ),
    .S(net429),
    .Y(_08800_));
 sky130_fd_sc_hd__mux2i_1 _16044_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[770] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[802] ),
    .S(net429),
    .Y(_08801_));
 sky130_fd_sc_hd__a22oi_1 _16045_ (.A1(net624),
    .A2(_08800_),
    .B1(_08801_),
    .B2(net1195),
    .Y(_08802_));
 sky130_fd_sc_hd__and2_4 _16046_ (.A(net397),
    .B(net403),
    .X(_08803_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_972 ();
 sky130_fd_sc_hd__mux2i_1 _16048_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[962] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[994] ),
    .S(net1122),
    .Y(_08805_));
 sky130_fd_sc_hd__mux2i_1 _16049_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[834] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[866] ),
    .S(net430),
    .Y(_08806_));
 sky130_fd_sc_hd__nor2b_4 _16050_ (.A(net393),
    .B_N(net406),
    .Y(_08807_));
 sky130_fd_sc_hd__a22oi_1 _16051_ (.A1(_08803_),
    .A2(_08805_),
    .B1(_08806_),
    .B2(net615),
    .Y(_08808_));
 sky130_fd_sc_hd__nand2_8 _16052_ (.A(net383),
    .B(net1108),
    .Y(_08809_));
 sky130_fd_sc_hd__a21oi_2 _16053_ (.A1(_08802_),
    .A2(_08808_),
    .B1(_08809_),
    .Y(_08810_));
 sky130_fd_sc_hd__nand2b_4 _16054_ (.A_N(net403),
    .B(net397),
    .Y(_08811_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_971 ();
 sky130_fd_sc_hd__mux2i_1 _16056_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[130] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[162] ),
    .S(net433),
    .Y(_08813_));
 sky130_fd_sc_hd__nor2_1 _16057_ (.A(_08811_),
    .B(_08813_),
    .Y(_08814_));
 sky130_fd_sc_hd__nand2_8 _16058_ (.A(net397),
    .B(net403),
    .Y(_08815_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_970 ();
 sky130_fd_sc_hd__mux2i_1 _16060_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[194] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[226] ),
    .S(net433),
    .Y(_08817_));
 sky130_fd_sc_hd__mux2i_1 _16061_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[66] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[98] ),
    .S(net433),
    .Y(_08818_));
 sky130_fd_sc_hd__nand2b_4 _16062_ (.A_N(net397),
    .B(net403),
    .Y(_08819_));
 sky130_fd_sc_hd__o22ai_1 _16063_ (.A1(_08815_),
    .A2(_08817_),
    .B1(_08818_),
    .B2(_08819_),
    .Y(_08820_));
 sky130_fd_sc_hd__or2_4 _16064_ (.A(net385),
    .B(net389),
    .X(_08821_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_969 ();
 sky130_fd_sc_hd__a31o_1 _16066_ (.A1(net433),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[34] ),
    .A3(net1195),
    .B1(_08821_),
    .X(_08823_));
 sky130_fd_sc_hd__nor3_2 _16067_ (.A(_08814_),
    .B(_08820_),
    .C(_08823_),
    .Y(_08824_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_968 ();
 sky130_fd_sc_hd__mux2i_4 _16069_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[514] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[546] ),
    .S(net421),
    .Y(_08826_));
 sky130_fd_sc_hd__mux2i_1 _16070_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[450] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[482] ),
    .S(net901),
    .Y(_08827_));
 sky130_fd_sc_hd__a22oi_4 _16071_ (.A1(_08826_),
    .A2(net586),
    .B1(_08827_),
    .B2(_08593_),
    .Y(_08828_));
 sky130_fd_sc_hd__mux2i_1 _16072_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[258] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[290] ),
    .S(net421),
    .Y(_08829_));
 sky130_fd_sc_hd__mux2i_1 _16073_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[706] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[738] ),
    .S(net1283),
    .Y(_08830_));
 sky130_fd_sc_hd__a22oi_2 _16074_ (.A1(_08829_),
    .A2(net556),
    .B1(_08830_),
    .B2(_08602_),
    .Y(_08831_));
 sky130_fd_sc_hd__mux2i_1 _16075_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[386] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[418] ),
    .S(net421),
    .Y(_08832_));
 sky130_fd_sc_hd__mux2i_1 _16076_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[322] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[354] ),
    .S(net1283),
    .Y(_08833_));
 sky130_fd_sc_hd__a22oi_4 _16077_ (.A1(net569),
    .A2(_08832_),
    .B1(_08833_),
    .B2(net550),
    .Y(_08834_));
 sky130_fd_sc_hd__mux2i_1 _16078_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[642] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[674] ),
    .S(net421),
    .Y(_08835_));
 sky130_fd_sc_hd__mux2i_1 _16079_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[578] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[610] ),
    .S(net1283),
    .Y(_08836_));
 sky130_fd_sc_hd__a22oi_4 _16080_ (.A1(net758),
    .A2(_08835_),
    .B1(_08836_),
    .B2(net536),
    .Y(_08837_));
 sky130_fd_sc_hd__nand4_4 _16081_ (.A(_08837_),
    .B(_08831_),
    .C(_08828_),
    .D(_08834_),
    .Y(_08838_));
 sky130_fd_sc_hd__or3_4 _16082_ (.A(_08838_),
    .B(_08824_),
    .C(_08810_),
    .X(_08839_));
 sky130_fd_sc_hd__o22ai_1 _16083_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[34] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[2] ),
    .B2(_08503_),
    .Y(_08840_));
 sky130_fd_sc_hd__a21oi_2 _16084_ (.A1(_08839_),
    .A2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .B1(_08840_),
    .Y(_08841_));
 sky130_fd_sc_hd__o21ai_0 _16085_ (.A1(_08504_),
    .A2(_08795_),
    .B1(_08841_),
    .Y(_08842_));
 sky130_fd_sc_hd__nand2_1 _16086_ (.A(_08272_),
    .B(_08842_),
    .Y(_08843_));
 sky130_fd_sc_hd__o21ai_2 _16087_ (.A1(_08272_),
    .A2(_08797_),
    .B1(_08843_),
    .Y(_08844_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_966 ();
 sky130_fd_sc_hd__a21oi_1 _16090_ (.A1(net661),
    .A2(_08632_),
    .B1(_08579_),
    .Y(_08847_));
 sky130_fd_sc_hd__nor2_1 _16091_ (.A(\cs_registers_i.pc_id_i[2] ),
    .B(_08578_),
    .Y(_08848_));
 sky130_fd_sc_hd__a2111oi_4 _16092_ (.A1(_08839_),
    .A2(_08577_),
    .B1(_08847_),
    .C1(_08848_),
    .D1(_08368_),
    .Y(_08849_));
 sky130_fd_sc_hd__a21oi_4 _16093_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[2] ),
    .A2(_08368_),
    .B1(_08849_),
    .Y(_08850_));
 sky130_fd_sc_hd__a21oi_1 _16094_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[34] ),
    .A2(_08377_),
    .B1(_08295_),
    .Y(_08851_));
 sky130_fd_sc_hd__a21oi_4 _16095_ (.A1(_08850_),
    .A2(net1134),
    .B1(_08851_),
    .Y(_08852_));
 sky130_fd_sc_hd__or2_1 _16096_ (.A(_08852_),
    .B(_08844_),
    .X(_08853_));
 sky130_fd_sc_hd__inv_1 _16097_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[0] ),
    .Y(_08854_));
 sky130_fd_sc_hd__nand2_1 _16098_ (.A(net571),
    .B(_08632_),
    .Y(_08855_));
 sky130_fd_sc_hd__mux2i_4 _16099_ (.A0(_08854_),
    .A1(_08855_),
    .S(net940),
    .Y(_08856_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_962 ();
 sky130_fd_sc_hd__mux2i_1 _16104_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[896] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[928] ),
    .S(net433),
    .Y(_08861_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_960 ();
 sky130_fd_sc_hd__mux2i_1 _16107_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[768] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[800] ),
    .S(net433),
    .Y(_08864_));
 sky130_fd_sc_hd__a22oi_2 _16108_ (.A1(net323),
    .A2(_08861_),
    .B1(_08864_),
    .B2(net1195),
    .Y(_08865_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_959 ();
 sky130_fd_sc_hd__mux2i_1 _16110_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[960] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[992] ),
    .S(net433),
    .Y(_08867_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_957 ();
 sky130_fd_sc_hd__mux2i_1 _16113_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[832] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[864] ),
    .S(net433),
    .Y(_08870_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_956 ();
 sky130_fd_sc_hd__a22oi_2 _16115_ (.A1(_08803_),
    .A2(_08867_),
    .B1(_08870_),
    .B2(net614),
    .Y(_08872_));
 sky130_fd_sc_hd__a21oi_4 _16116_ (.A1(_08865_),
    .A2(_08872_),
    .B1(_08809_),
    .Y(_08873_));
 sky130_fd_sc_hd__mux2i_1 _16117_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[704] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[736] ),
    .S(net428),
    .Y(_08874_));
 sky130_fd_sc_hd__mux2i_1 _16118_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[640] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[672] ),
    .S(net428),
    .Y(_08875_));
 sky130_fd_sc_hd__a22oi_4 _16119_ (.A1(_08602_),
    .A2(_08874_),
    .B1(_08875_),
    .B2(net1002),
    .Y(_08876_));
 sky130_fd_sc_hd__mux2i_2 _16120_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[512] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[544] ),
    .S(net428),
    .Y(_08877_));
 sky130_fd_sc_hd__mux2i_1 _16121_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[320] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[352] ),
    .S(net1122),
    .Y(_08878_));
 sky130_fd_sc_hd__a22oi_2 _16122_ (.A1(_08877_),
    .A2(_08599_),
    .B1(_08878_),
    .B2(net875),
    .Y(_08879_));
 sky130_fd_sc_hd__mux2i_1 _16123_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[256] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[288] ),
    .S(net1122),
    .Y(_08880_));
 sky130_fd_sc_hd__mux2i_1 _16124_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[448] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[480] ),
    .S(net428),
    .Y(_08881_));
 sky130_fd_sc_hd__a22oi_2 _16125_ (.A1(_08597_),
    .A2(_08880_),
    .B1(_08881_),
    .B2(_08593_),
    .Y(_08882_));
 sky130_fd_sc_hd__mux2i_2 _16126_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[576] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[608] ),
    .S(net428),
    .Y(_08883_));
 sky130_fd_sc_hd__mux2i_2 _16127_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[384] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[416] ),
    .S(net428),
    .Y(_08884_));
 sky130_fd_sc_hd__a22oi_2 _16128_ (.A1(net955),
    .A2(_08883_),
    .B1(_08884_),
    .B2(net1118),
    .Y(_08885_));
 sky130_fd_sc_hd__nand4_4 _16129_ (.A(_08879_),
    .B(_08876_),
    .C(_08882_),
    .D(_08885_),
    .Y(_08886_));
 sky130_fd_sc_hd__mux2i_1 _16130_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[64] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[96] ),
    .S(net434),
    .Y(_08887_));
 sky130_fd_sc_hd__mux2i_1 _16131_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[128] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[160] ),
    .S(net434),
    .Y(_08888_));
 sky130_fd_sc_hd__o22ai_2 _16132_ (.A1(_08819_),
    .A2(_08887_),
    .B1(_08888_),
    .B2(_08811_),
    .Y(_08889_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_954 ();
 sky130_fd_sc_hd__mux2_1 _16135_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[192] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[224] ),
    .S(net434),
    .X(_08892_));
 sky130_fd_sc_hd__a32o_1 _16136_ (.A1(net434),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[32] ),
    .A3(net1197),
    .B1(_08803_),
    .B2(_08892_),
    .X(_08893_));
 sky130_fd_sc_hd__nor3_4 _16137_ (.A(_08821_),
    .B(_08889_),
    .C(_08893_),
    .Y(_08894_));
 sky130_fd_sc_hd__nor3_4 _16138_ (.A(_08886_),
    .B(_08873_),
    .C(_08894_),
    .Y(_08895_));
 sky130_fd_sc_hd__nor3b_4 _16139_ (.A(net1115),
    .B(net310),
    .C_N(net495),
    .Y(_08896_));
 sky130_fd_sc_hd__a21oi_4 _16140_ (.A1(net1115),
    .A2(_08856_),
    .B1(_08896_),
    .Y(_08897_));
 sky130_fd_sc_hd__nand2_1 _16141_ (.A(_08642_),
    .B(_08640_),
    .Y(_08898_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_953 ();
 sky130_fd_sc_hd__mux2i_2 _16143_ (.A0(net1133),
    .A1(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .S(_08643_),
    .Y(_08900_));
 sky130_fd_sc_hd__nand4b_4 _16144_ (.A_N(net376),
    .B(net339),
    .C(net332),
    .D(net335),
    .Y(_08901_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_949 ();
 sky130_fd_sc_hd__mux2i_2 _16149_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[896] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[960] ),
    .S(net361),
    .Y(_08906_));
 sky130_fd_sc_hd__mux2i_2 _16150_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[800] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[864] ),
    .S(net362),
    .Y(_08907_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_948 ();
 sky130_fd_sc_hd__o22ai_4 _16152_ (.A1(net934),
    .A2(_08906_),
    .B1(_08907_),
    .B2(net930),
    .Y(_08909_));
 sky130_fd_sc_hd__nand4_4 _16153_ (.A(net376),
    .B(net335),
    .C(net332),
    .D(net339),
    .Y(_08910_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_947 ();
 sky130_fd_sc_hd__mux2i_2 _16155_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[928] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[992] ),
    .S(net361),
    .Y(_08912_));
 sky130_fd_sc_hd__mux2i_2 _16156_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[768] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[832] ),
    .S(net362),
    .Y(_08913_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_946 ();
 sky130_fd_sc_hd__o22ai_4 _16158_ (.A1(net1210),
    .A2(_08912_),
    .B1(_08913_),
    .B2(net506),
    .Y(_08915_));
 sky130_fd_sc_hd__nor2_4 _16159_ (.A(_08909_),
    .B(_08915_),
    .Y(_08916_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_943 ();
 sky130_fd_sc_hd__mux4_1 _16163_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[128] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[160] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[192] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[224] ),
    .S0(net374),
    .S1(net363),
    .X(_08920_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_941 ();
 sky130_fd_sc_hd__mux2_1 _16166_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[32] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[96] ),
    .S(net363),
    .X(_08923_));
 sky130_fd_sc_hd__a221o_1 _16167_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[64] ),
    .A2(net324),
    .B1(_08923_),
    .B2(net1133),
    .C1(net341),
    .X(_08924_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_940 ();
 sky130_fd_sc_hd__o211ai_4 _16169_ (.A1(_08481_),
    .A2(_08920_),
    .B1(_08924_),
    .C1(_08731_),
    .Y(_08926_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_936 ();
 sky130_fd_sc_hd__mux2i_1 _16174_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[544] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[608] ),
    .S(net357),
    .Y(_08931_));
 sky130_fd_sc_hd__mux2i_1 _16175_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[640] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[704] ),
    .S(net357),
    .Y(_08932_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_934 ();
 sky130_fd_sc_hd__a22oi_2 _16178_ (.A1(_08931_),
    .A2(net329),
    .B1(_08932_),
    .B2(net326),
    .Y(_08935_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_933 ();
 sky130_fd_sc_hd__mux2i_1 _16180_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[512] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[576] ),
    .S(net357),
    .Y(_08937_));
 sky130_fd_sc_hd__mux2i_1 _16181_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[672] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[736] ),
    .S(net357),
    .Y(_08938_));
 sky130_fd_sc_hd__a22oi_2 _16182_ (.A1(_08937_),
    .A2(net325),
    .B1(_08938_),
    .B2(net1024),
    .Y(_08939_));
 sky130_fd_sc_hd__nand3_4 _16183_ (.A(_08462_),
    .B(_08939_),
    .C(_08935_),
    .Y(_08940_));
 sky130_fd_sc_hd__mux2i_1 _16184_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[384] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[448] ),
    .S(net357),
    .Y(_08941_));
 sky130_fd_sc_hd__mux2i_1 _16185_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[256] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[320] ),
    .S(net357),
    .Y(_08942_));
 sky130_fd_sc_hd__a22oi_2 _16186_ (.A1(net326),
    .A2(_08941_),
    .B1(_08942_),
    .B2(net325),
    .Y(_08943_));
 sky130_fd_sc_hd__mux2i_2 _16187_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[288] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[352] ),
    .S(net357),
    .Y(_08944_));
 sky130_fd_sc_hd__mux2i_1 _16188_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[416] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[480] ),
    .S(net357),
    .Y(_08945_));
 sky130_fd_sc_hd__a22oi_2 _16189_ (.A1(net329),
    .A2(_08944_),
    .B1(_08945_),
    .B2(net1024),
    .Y(_08946_));
 sky130_fd_sc_hd__nand3_4 _16190_ (.A(_08946_),
    .B(_08943_),
    .C(net704),
    .Y(_08947_));
 sky130_fd_sc_hd__and4_4 _16191_ (.A(_08916_),
    .B(_08926_),
    .C(_08940_),
    .D(_08947_),
    .X(_08948_));
 sky130_fd_sc_hd__o32ai_4 _16192_ (.A1(_08898_),
    .A2(_08639_),
    .A3(_08900_),
    .B1(_08436_),
    .B2(_08948_),
    .Y(_08949_));
 sky130_fd_sc_hd__nand4_4 _16193_ (.A(_08916_),
    .B(_08926_),
    .C(_08940_),
    .D(_08947_),
    .Y(_08950_));
 sky130_fd_sc_hd__o22ai_1 _16194_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[32] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[0] ),
    .B2(_08503_),
    .Y(_08951_));
 sky130_fd_sc_hd__nor2_1 _16195_ (.A(_08295_),
    .B(_08951_),
    .Y(_08952_));
 sky130_fd_sc_hd__o221ai_4 _16196_ (.A1(_08500_),
    .A2(net495),
    .B1(_08504_),
    .B2(_08950_),
    .C1(_08952_),
    .Y(_08953_));
 sky130_fd_sc_hd__nand2_1 _16197_ (.A(_08949_),
    .B(_08953_),
    .Y(_08954_));
 sky130_fd_sc_hd__a22o_1 _16198_ (.A1(_08897_),
    .A2(_08949_),
    .B1(_08954_),
    .B2(net296),
    .X(_08955_));
 sky130_fd_sc_hd__a21oi_1 _16199_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[32] ),
    .A2(_08377_),
    .B1(_08953_),
    .Y(_08956_));
 sky130_fd_sc_hd__a21oi_4 _16200_ (.A1(_08295_),
    .A2(_08955_),
    .B1(_08956_),
    .Y(_08957_));
 sky130_fd_sc_hd__nand2b_1 _16201_ (.A_N(_08643_),
    .B(net372),
    .Y(_08958_));
 sky130_fd_sc_hd__nand3_1 _16202_ (.A(\id_stage_i.controller_i.instr_is_compressed_i ),
    .B(_08444_),
    .C(_08643_),
    .Y(_08959_));
 sky130_fd_sc_hd__a21oi_1 _16203_ (.A1(_08958_),
    .A2(_08959_),
    .B1(_08439_),
    .Y(_08960_));
 sky130_fd_sc_hd__and3_1 _16204_ (.A(net1021),
    .B(_08640_),
    .C(_08644_),
    .X(_08961_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_931 ();
 sky130_fd_sc_hd__mux4_2 _16207_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[129] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[161] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[193] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[225] ),
    .S0(net374),
    .S1(net363),
    .X(_08964_));
 sky130_fd_sc_hd__mux2_1 _16208_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[33] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[97] ),
    .S(net363),
    .X(_08965_));
 sky130_fd_sc_hd__a221o_1 _16209_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[65] ),
    .A2(net324),
    .B1(net374),
    .B2(_08965_),
    .C1(net341),
    .X(_08966_));
 sky130_fd_sc_hd__o211ai_4 _16210_ (.A1(_08964_),
    .A2(_08481_),
    .B1(_08966_),
    .C1(_08731_),
    .Y(_08967_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_929 ();
 sky130_fd_sc_hd__mux2i_1 _16213_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[513] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[577] ),
    .S(net360),
    .Y(_08970_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_927 ();
 sky130_fd_sc_hd__mux2i_1 _16216_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[545] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[609] ),
    .S(net360),
    .Y(_08973_));
 sky130_fd_sc_hd__a22oi_1 _16217_ (.A1(_08970_),
    .A2(net325),
    .B1(_08973_),
    .B2(net328),
    .Y(_08974_));
 sky130_fd_sc_hd__mux2i_1 _16218_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[641] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[705] ),
    .S(net360),
    .Y(_08975_));
 sky130_fd_sc_hd__mux2i_1 _16219_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[673] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[737] ),
    .S(net360),
    .Y(_08976_));
 sky130_fd_sc_hd__a22oi_1 _16220_ (.A1(net326),
    .A2(_08975_),
    .B1(_08976_),
    .B2(_08152_),
    .Y(_08977_));
 sky130_fd_sc_hd__nand3_2 _16221_ (.A(_08462_),
    .B(_08977_),
    .C(_08974_),
    .Y(_08978_));
 sky130_fd_sc_hd__mux2i_1 _16222_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[769] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[833] ),
    .S(net360),
    .Y(_08979_));
 sky130_fd_sc_hd__mux2i_1 _16223_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[897] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[961] ),
    .S(net360),
    .Y(_08980_));
 sky130_fd_sc_hd__a22oi_1 _16224_ (.A1(net325),
    .A2(_08979_),
    .B1(_08980_),
    .B2(net326),
    .Y(_08981_));
 sky130_fd_sc_hd__mux2i_1 _16225_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[801] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[865] ),
    .S(net360),
    .Y(_08982_));
 sky130_fd_sc_hd__nand2_1 _16226_ (.A(net328),
    .B(_08982_),
    .Y(_08983_));
 sky130_fd_sc_hd__mux2i_1 _16227_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[929] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[993] ),
    .S(net360),
    .Y(_08984_));
 sky130_fd_sc_hd__a21oi_1 _16228_ (.A1(_08152_),
    .A2(_08984_),
    .B1(_08708_),
    .Y(_08985_));
 sky130_fd_sc_hd__nand3_2 _16229_ (.A(_08981_),
    .B(_08985_),
    .C(_08983_),
    .Y(_08986_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_926 ();
 sky130_fd_sc_hd__mux2i_1 _16231_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[289] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[353] ),
    .S(net360),
    .Y(_08988_));
 sky130_fd_sc_hd__mux2i_1 _16232_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[257] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[321] ),
    .S(net360),
    .Y(_08989_));
 sky130_fd_sc_hd__a22oi_1 _16233_ (.A1(net328),
    .A2(_08988_),
    .B1(_08989_),
    .B2(net325),
    .Y(_08990_));
 sky130_fd_sc_hd__mux2i_1 _16234_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[417] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[481] ),
    .S(net360),
    .Y(_08991_));
 sky130_fd_sc_hd__mux2i_1 _16235_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[385] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[449] ),
    .S(net360),
    .Y(_08992_));
 sky130_fd_sc_hd__a22oi_1 _16236_ (.A1(_08152_),
    .A2(_08991_),
    .B1(_08992_),
    .B2(net326),
    .Y(_08993_));
 sky130_fd_sc_hd__nand3_2 _16237_ (.A(_08993_),
    .B(_08990_),
    .C(net700),
    .Y(_08994_));
 sky130_fd_sc_hd__and4_4 _16238_ (.A(_08967_),
    .B(_08994_),
    .C(_08986_),
    .D(_08978_),
    .X(_08995_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_924 ();
 sky130_fd_sc_hd__nand2_4 _16241_ (.A(_08495_),
    .B(_08995_),
    .Y(_08998_));
 sky130_fd_sc_hd__o31a_4 _16242_ (.A1(_08495_),
    .A2(_08960_),
    .A3(_08961_),
    .B1(_08998_),
    .X(_08999_));
 sky130_fd_sc_hd__xnor2_1 _16243_ (.A(net296),
    .B(_08999_),
    .Y(_09000_));
 sky130_fd_sc_hd__nand2b_1 _16244_ (.A_N(net395),
    .B(net1082),
    .Y(_09001_));
 sky130_fd_sc_hd__mux4_2 _16245_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[257] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[289] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[321] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[353] ),
    .S0(net430),
    .S1(net406),
    .X(_09002_));
 sky130_fd_sc_hd__nor2_1 _16246_ (.A(_09001_),
    .B(_09002_),
    .Y(_09003_));
 sky130_fd_sc_hd__nand3_1 _16247_ (.A(net1082),
    .B(net395),
    .C(net406),
    .Y(_09004_));
 sky130_fd_sc_hd__nor2b_1 _16248_ (.A(net1122),
    .B_N(\gen_regfile_ff.register_file_i.rf_reg[449] ),
    .Y(_09005_));
 sky130_fd_sc_hd__a211oi_1 _16249_ (.A1(net1122),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[481] ),
    .B1(_09004_),
    .C1(_09005_),
    .Y(_09006_));
 sky130_fd_sc_hd__nand2_1 _16250_ (.A(net1082),
    .B(net395),
    .Y(_09007_));
 sky130_fd_sc_hd__nor2b_1 _16251_ (.A(net430),
    .B_N(\gen_regfile_ff.register_file_i.rf_reg[385] ),
    .Y(_09008_));
 sky130_fd_sc_hd__a2111oi_2 _16252_ (.A1(net912),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[417] ),
    .B1(_09007_),
    .C1(_09008_),
    .D1(net406),
    .Y(_09009_));
 sky130_fd_sc_hd__or4_4 _16253_ (.A(net384),
    .B(_09009_),
    .C(_09006_),
    .D(_09003_),
    .X(_09010_));
 sky130_fd_sc_hd__mux2i_1 _16254_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[193] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[225] ),
    .S(net434),
    .Y(_09011_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_923 ();
 sky130_fd_sc_hd__mux2i_1 _16256_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[129] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[161] ),
    .S(net434),
    .Y(_09013_));
 sky130_fd_sc_hd__a22oi_1 _16257_ (.A1(_08803_),
    .A2(_09011_),
    .B1(_09013_),
    .B2(net323),
    .Y(_09014_));
 sky130_fd_sc_hd__mux2i_1 _16258_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[65] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[97] ),
    .S(net434),
    .Y(_09015_));
 sky130_fd_sc_hd__nand3b_1 _16259_ (.A_N(net402),
    .B(\gen_regfile_ff.register_file_i.rf_reg[33] ),
    .C(net434),
    .Y(_09016_));
 sky130_fd_sc_hd__o211ai_2 _16260_ (.A1(_08627_),
    .A2(_09015_),
    .B1(_09016_),
    .C1(_08529_),
    .Y(_09017_));
 sky130_fd_sc_hd__a21oi_2 _16261_ (.A1(_09017_),
    .A2(_09014_),
    .B1(net389),
    .Y(_09018_));
 sky130_fd_sc_hd__mux2i_1 _16262_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[769] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[801] ),
    .S(net432),
    .Y(_09019_));
 sky130_fd_sc_hd__mux2i_1 _16263_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[897] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[929] ),
    .S(net432),
    .Y(_09020_));
 sky130_fd_sc_hd__a22oi_2 _16264_ (.A1(net1195),
    .A2(_09019_),
    .B1(_09020_),
    .B2(net624),
    .Y(_09021_));
 sky130_fd_sc_hd__mux2i_2 _16265_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[833] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[865] ),
    .S(net432),
    .Y(_09022_));
 sky130_fd_sc_hd__mux2i_1 _16266_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[961] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[993] ),
    .S(net432),
    .Y(_09023_));
 sky130_fd_sc_hd__a22oi_2 _16267_ (.A1(net614),
    .A2(_09022_),
    .B1(_09023_),
    .B2(_08803_),
    .Y(_09024_));
 sky130_fd_sc_hd__nand3_4 _16268_ (.A(_08618_),
    .B(_09021_),
    .C(_09024_),
    .Y(_09025_));
 sky130_fd_sc_hd__mux2i_1 _16269_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[641] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[673] ),
    .S(net432),
    .Y(_09026_));
 sky130_fd_sc_hd__nand2_1 _16270_ (.A(net624),
    .B(_09026_),
    .Y(_09027_));
 sky130_fd_sc_hd__mux2i_1 _16271_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[577] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[609] ),
    .S(net432),
    .Y(_09028_));
 sky130_fd_sc_hd__mux2i_1 _16272_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[513] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[545] ),
    .S(net432),
    .Y(_09029_));
 sky130_fd_sc_hd__a22oi_1 _16273_ (.A1(net614),
    .A2(_09028_),
    .B1(_09029_),
    .B2(net1195),
    .Y(_09030_));
 sky130_fd_sc_hd__mux2i_1 _16274_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[705] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[737] ),
    .S(net432),
    .Y(_09031_));
 sky130_fd_sc_hd__nand2b_4 _16275_ (.A_N(net1082),
    .B(net383),
    .Y(_09032_));
 sky130_fd_sc_hd__a21oi_1 _16276_ (.A1(_08803_),
    .A2(_09031_),
    .B1(_09032_),
    .Y(_09033_));
 sky130_fd_sc_hd__nand3_2 _16277_ (.A(_09027_),
    .B(_09030_),
    .C(_09033_),
    .Y(_09034_));
 sky130_fd_sc_hd__o211ai_4 _16278_ (.A1(_09018_),
    .A2(_09010_),
    .B1(_09025_),
    .C1(_09034_),
    .Y(_09035_));
 sky130_fd_sc_hd__o22ai_1 _16279_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[33] ),
    .A2(_08502_),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[1] ),
    .B2(_08503_),
    .Y(_09036_));
 sky130_fd_sc_hd__a21oi_2 _16280_ (.A1(_08696_),
    .A2(net981),
    .B1(_09036_),
    .Y(_09037_));
 sky130_fd_sc_hd__o211ai_2 _16281_ (.A1(_08500_),
    .A2(net559),
    .B1(_09037_),
    .C1(net314),
    .Y(_09038_));
 sky130_fd_sc_hd__o21a_2 _16282_ (.A1(net314),
    .A2(_09000_),
    .B1(_09038_),
    .X(_09039_));
 sky130_fd_sc_hd__nor3_2 _16283_ (.A(_08307_),
    .B(_08576_),
    .C(net559),
    .Y(_09040_));
 sky130_fd_sc_hd__nor2_1 _16284_ (.A(_08627_),
    .B(_08581_),
    .Y(_09041_));
 sky130_fd_sc_hd__o22ai_1 _16285_ (.A1(\cs_registers_i.pc_id_i[1] ),
    .A2(_08578_),
    .B1(_08579_),
    .B2(_09041_),
    .Y(_09042_));
 sky130_fd_sc_hd__nor3_2 _16286_ (.A(_08368_),
    .B(_09040_),
    .C(_09042_),
    .Y(_09043_));
 sky130_fd_sc_hd__a21oi_4 _16287_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[1] ),
    .A2(_08368_),
    .B1(_09043_),
    .Y(_09044_));
 sky130_fd_sc_hd__a21oi_1 _16288_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[33] ),
    .A2(_08377_),
    .B1(_08295_),
    .Y(_09045_));
 sky130_fd_sc_hd__a21oi_4 _16289_ (.A1(_09044_),
    .A2(_08295_),
    .B1(_09045_),
    .Y(_09046_));
 sky130_fd_sc_hd__maj3_2 _16290_ (.A(_08957_),
    .B(_09039_),
    .C(_09046_),
    .X(_09047_));
 sky130_fd_sc_hd__and2_1 _16291_ (.A(_08638_),
    .B(_08700_),
    .X(_09048_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_922 ();
 sky130_fd_sc_hd__o21a_1 _16293_ (.A1(_08272_),
    .A2(_08585_),
    .B1(_08588_),
    .X(_09050_));
 sky130_fd_sc_hd__a211oi_2 _16294_ (.A1(_08746_),
    .A2(_08290_),
    .B1(_08750_),
    .C1(_09050_),
    .Y(_09051_));
 sky130_fd_sc_hd__and2_0 _16295_ (.A(_08844_),
    .B(_08852_),
    .X(_09052_));
 sky130_fd_sc_hd__a2111o_2 _16296_ (.A1(_09047_),
    .A2(_08853_),
    .B1(_09048_),
    .C1(_09051_),
    .D1(_09052_),
    .X(_09053_));
 sky130_fd_sc_hd__or4b_4 _16297_ (.A(net333),
    .B(net376),
    .C(net338),
    .D_N(net335),
    .X(_09054_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_921 ();
 sky130_fd_sc_hd__mux2i_1 _16299_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[261] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[325] ),
    .S(net370),
    .Y(_09056_));
 sky130_fd_sc_hd__mux2i_1 _16300_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[805] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[869] ),
    .S(net370),
    .Y(_09057_));
 sky130_fd_sc_hd__o22ai_1 _16301_ (.A1(net807),
    .A2(_09056_),
    .B1(_09057_),
    .B2(net523),
    .Y(_09058_));
 sky130_fd_sc_hd__mux2i_1 _16302_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[773] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[837] ),
    .S(net370),
    .Y(_09059_));
 sky130_fd_sc_hd__nand4bb_4 _16303_ (.A_N(net333),
    .B_N(net338),
    .C(net376),
    .D(net335),
    .Y(_09060_));
 sky130_fd_sc_hd__mux2i_1 _16304_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[293] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[357] ),
    .S(net370),
    .Y(_09061_));
 sky130_fd_sc_hd__o22ai_1 _16305_ (.A1(net501),
    .A2(_09059_),
    .B1(_09060_),
    .B2(_09061_),
    .Y(_09062_));
 sky130_fd_sc_hd__nor2_2 _16306_ (.A(_09058_),
    .B(_09062_),
    .Y(_09063_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_920 ();
 sky130_fd_sc_hd__mux4_2 _16308_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[133] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[165] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[197] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[229] ),
    .S0(net379),
    .S1(net371),
    .X(_09065_));
 sky130_fd_sc_hd__mux2_1 _16309_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[37] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[101] ),
    .S(net367),
    .X(_09066_));
 sky130_fd_sc_hd__a221o_1 _16310_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[69] ),
    .A2(_08484_),
    .B1(_09066_),
    .B2(net1220),
    .C1(net343),
    .X(_09067_));
 sky130_fd_sc_hd__o211ai_4 _16311_ (.A1(_08481_),
    .A2(_09065_),
    .B1(_09067_),
    .C1(_08731_),
    .Y(_09068_));
 sky130_fd_sc_hd__mux4_1 _16312_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[901] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[933] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[965] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[997] ),
    .S0(net379),
    .S1(net371),
    .X(_09069_));
 sky130_fd_sc_hd__nor2_1 _16313_ (.A(net334),
    .B(net379),
    .Y(_09070_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_919 ();
 sky130_fd_sc_hd__mux2i_1 _16315_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[389] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[453] ),
    .S(net371),
    .Y(_09072_));
 sky130_fd_sc_hd__nor2b_1 _16316_ (.A(net334),
    .B_N(net379),
    .Y(_09073_));
 sky130_fd_sc_hd__mux2i_1 _16317_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[421] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[485] ),
    .S(net371),
    .Y(_09074_));
 sky130_fd_sc_hd__nand2_2 _16318_ (.A(net337),
    .B(net339),
    .Y(_09075_));
 sky130_fd_sc_hd__a221oi_2 _16319_ (.A1(_09070_),
    .A2(_09072_),
    .B1(_09073_),
    .B2(_09074_),
    .C1(_09075_),
    .Y(_09076_));
 sky130_fd_sc_hd__o21ai_2 _16320_ (.A1(_08161_),
    .A2(_09069_),
    .B1(_09076_),
    .Y(_09077_));
 sky130_fd_sc_hd__mux2i_1 _16321_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[549] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[613] ),
    .S(net1142),
    .Y(_09078_));
 sky130_fd_sc_hd__mux2i_1 _16322_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[645] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[709] ),
    .S(net346),
    .Y(_09079_));
 sky130_fd_sc_hd__a22oi_1 _16323_ (.A1(net889),
    .A2(_09078_),
    .B1(_09079_),
    .B2(net589),
    .Y(_09080_));
 sky130_fd_sc_hd__mux2i_1 _16324_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[517] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[581] ),
    .S(net1142),
    .Y(_09081_));
 sky130_fd_sc_hd__mux2i_1 _16325_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[677] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[741] ),
    .S(net1142),
    .Y(_09082_));
 sky130_fd_sc_hd__a22oi_1 _16326_ (.A1(net1046),
    .A2(_09081_),
    .B1(_09082_),
    .B2(_08152_),
    .Y(_09083_));
 sky130_fd_sc_hd__nand3_1 _16327_ (.A(_08462_),
    .B(_09080_),
    .C(_09083_),
    .Y(_09084_));
 sky130_fd_sc_hd__nand4_4 _16328_ (.A(_09063_),
    .B(_09068_),
    .C(_09077_),
    .D(_09084_),
    .Y(_09085_));
 sky130_fd_sc_hd__a22oi_4 _16329_ (.A1(net581),
    .A2(_08450_),
    .B1(_08495_),
    .B2(_09085_),
    .Y(_09086_));
 sky130_fd_sc_hd__xnor2_1 _16330_ (.A(net695),
    .B(_09086_),
    .Y(_09087_));
 sky130_fd_sc_hd__mux4_1 _16331_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[645] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[677] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[709] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[741] ),
    .S0(net420),
    .S1(net1112),
    .X(_09088_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_918 ();
 sky130_fd_sc_hd__mux4_2 _16333_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[901] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[933] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[965] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[997] ),
    .S0(net419),
    .S1(net412),
    .X(_09090_));
 sky130_fd_sc_hd__a22oi_2 _16334_ (.A1(net1247),
    .A2(_09088_),
    .B1(_09090_),
    .B2(_08324_),
    .Y(_09091_));
 sky130_fd_sc_hd__mux4_1 _16335_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[517] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[549] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[581] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[613] ),
    .S0(net420),
    .S1(net410),
    .X(_09092_));
 sky130_fd_sc_hd__mux4_1 _16336_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[773] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[805] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[837] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[869] ),
    .S0(net416),
    .S1(net1235),
    .X(_09093_));
 sky130_fd_sc_hd__a22oi_2 _16337_ (.A1(_08342_),
    .A2(_09092_),
    .B1(_09093_),
    .B2(net330),
    .Y(_09094_));
 sky130_fd_sc_hd__nand2_1 _16338_ (.A(_09091_),
    .B(_09094_),
    .Y(_09095_));
 sky130_fd_sc_hd__mux4_2 _16339_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[133] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[165] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[197] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[229] ),
    .S0(net440),
    .S1(net414),
    .X(_09096_));
 sky130_fd_sc_hd__nor2_2 _16340_ (.A(_08529_),
    .B(_09096_),
    .Y(_09097_));
 sky130_fd_sc_hd__mux2_1 _16341_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[69] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[101] ),
    .S(net439),
    .X(_09098_));
 sky130_fd_sc_hd__a221oi_4 _16342_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[37] ),
    .A2(_08321_),
    .B1(_09098_),
    .B2(net1072),
    .C1(net399),
    .Y(_09099_));
 sky130_fd_sc_hd__mux4_2 _16343_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[389] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[421] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[453] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[485] ),
    .S0(net419),
    .S1(net412),
    .X(_09100_));
 sky130_fd_sc_hd__mux4_1 _16344_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[261] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[293] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[325] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[357] ),
    .S0(net416),
    .S1(net1113),
    .X(_09101_));
 sky130_fd_sc_hd__a22oi_4 _16345_ (.A1(_08324_),
    .A2(_09100_),
    .B1(_09101_),
    .B2(net330),
    .Y(_09102_));
 sky130_fd_sc_hd__o311ai_4 _16346_ (.A1(net975),
    .A2(_09097_),
    .A3(_09099_),
    .B1(_09102_),
    .C1(_08512_),
    .Y(_09103_));
 sky130_fd_sc_hd__o21ai_4 _16347_ (.A1(_09095_),
    .A2(_08512_),
    .B1(_09103_),
    .Y(_09104_));
 sky130_fd_sc_hd__nor2_1 _16348_ (.A(_08504_),
    .B(_09085_),
    .Y(_09105_));
 sky130_fd_sc_hd__o22ai_2 _16349_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[37] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[5] ),
    .B2(_08503_),
    .Y(_09106_));
 sky130_fd_sc_hd__a2111oi_4 _16350_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(net796),
    .B1(_09106_),
    .C1(_09105_),
    .D1(_08295_),
    .Y(_09107_));
 sky130_fd_sc_hd__inv_1 _16351_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[5] ),
    .Y(_09108_));
 sky130_fd_sc_hd__mux2_1 _16352_ (.A0(_09108_),
    .A1(_09104_),
    .S(_08372_),
    .X(_09109_));
 sky130_fd_sc_hd__nand3_1 _16353_ (.A(\cs_registers_i.pc_id_i[5] ),
    .B(_08372_),
    .C(net941),
    .Y(_09110_));
 sky130_fd_sc_hd__o21ai_4 _16354_ (.A1(_09109_),
    .A2(net941),
    .B1(_09110_),
    .Y(_09111_));
 sky130_fd_sc_hd__and3_1 _16355_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[37] ),
    .B(net1106),
    .C(_08377_),
    .X(_09112_));
 sky130_fd_sc_hd__a21oi_1 _16356_ (.A1(_08295_),
    .A2(_09111_),
    .B1(_09112_),
    .Y(_09113_));
 sky130_fd_sc_hd__a211oi_4 _16357_ (.A1(_09087_),
    .A2(_08295_),
    .B1(_09107_),
    .C1(_09113_),
    .Y(_09114_));
 sky130_fd_sc_hd__a21o_1 _16358_ (.A1(_08295_),
    .A2(_09111_),
    .B1(_09112_),
    .X(_09115_));
 sky130_fd_sc_hd__a21oi_1 _16359_ (.A1(_08290_),
    .A2(_09087_),
    .B1(_09107_),
    .Y(_09116_));
 sky130_fd_sc_hd__nor2_1 _16360_ (.A(_09115_),
    .B(_09116_),
    .Y(_09117_));
 sky130_fd_sc_hd__nor2_2 _16361_ (.A(_09114_),
    .B(_09117_),
    .Y(_09118_));
 sky130_fd_sc_hd__a31oi_4 _16362_ (.A1(net1278),
    .A2(net880),
    .A3(_09118_),
    .B1(_09114_),
    .Y(_09119_));
 sky130_fd_sc_hd__mux4_2 _16363_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[134] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[166] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[198] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[230] ),
    .S0(net381),
    .S1(net513),
    .X(_09120_));
 sky130_fd_sc_hd__mux2_1 _16364_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[38] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[102] ),
    .S(net366),
    .X(_09121_));
 sky130_fd_sc_hd__a221o_1 _16365_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[70] ),
    .A2(_08484_),
    .B1(_09121_),
    .B2(net380),
    .C1(net343),
    .X(_09122_));
 sky130_fd_sc_hd__o211ai_4 _16366_ (.A1(_08481_),
    .A2(_09120_),
    .B1(_09122_),
    .C1(_08731_),
    .Y(_09123_));
 sky130_fd_sc_hd__mux2i_1 _16367_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[550] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[614] ),
    .S(net344),
    .Y(_09124_));
 sky130_fd_sc_hd__mux2i_1 _16368_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[646] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[710] ),
    .S(net344),
    .Y(_09125_));
 sky130_fd_sc_hd__a22oi_2 _16369_ (.A1(net1201),
    .A2(_09124_),
    .B1(_09125_),
    .B2(net1013),
    .Y(_09126_));
 sky130_fd_sc_hd__mux2i_1 _16370_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[518] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[582] ),
    .S(net344),
    .Y(_09127_));
 sky130_fd_sc_hd__mux2i_1 _16371_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[678] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[742] ),
    .S(net344),
    .Y(_09128_));
 sky130_fd_sc_hd__a22oi_2 _16372_ (.A1(net1043),
    .A2(_09127_),
    .B1(_09128_),
    .B2(net1153),
    .Y(_09129_));
 sky130_fd_sc_hd__nand3_4 _16373_ (.A(_08462_),
    .B(_09126_),
    .C(_09129_),
    .Y(_09130_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_917 ();
 sky130_fd_sc_hd__mux2i_1 _16375_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[422] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[486] ),
    .S(net368),
    .Y(_09132_));
 sky130_fd_sc_hd__mux2i_1 _16376_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[390] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[454] ),
    .S(net368),
    .Y(_09133_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_916 ();
 sky130_fd_sc_hd__o22ai_2 _16378_ (.A1(net866),
    .A2(_09132_),
    .B1(_09133_),
    .B2(net895),
    .Y(_09135_));
 sky130_fd_sc_hd__mux2i_1 _16379_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[902] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[966] ),
    .S(net368),
    .Y(_09136_));
 sky130_fd_sc_hd__mux2i_1 _16380_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[806] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[870] ),
    .S(net368),
    .Y(_09137_));
 sky130_fd_sc_hd__o22ai_2 _16381_ (.A1(net605),
    .A2(_09136_),
    .B1(_09137_),
    .B2(net525),
    .Y(_09138_));
 sky130_fd_sc_hd__mux2i_1 _16382_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[774] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[838] ),
    .S(net368),
    .Y(_09139_));
 sky130_fd_sc_hd__mux2i_1 _16383_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[294] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[358] ),
    .S(net368),
    .Y(_09140_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_915 ();
 sky130_fd_sc_hd__o22ai_2 _16385_ (.A1(net504),
    .A2(_09139_),
    .B1(_09140_),
    .B2(net764),
    .Y(_09142_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_914 ();
 sky130_fd_sc_hd__mux2i_1 _16387_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[262] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[326] ),
    .S(net368),
    .Y(_09144_));
 sky130_fd_sc_hd__mux2i_1 _16388_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[934] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[998] ),
    .S(net368),
    .Y(_09145_));
 sky130_fd_sc_hd__o22ai_4 _16389_ (.A1(net770),
    .A2(_09144_),
    .B1(_09145_),
    .B2(net633),
    .Y(_09146_));
 sky130_fd_sc_hd__nor4_4 _16390_ (.A(_09135_),
    .B(_09138_),
    .C(_09146_),
    .D(_09142_),
    .Y(_09147_));
 sky130_fd_sc_hd__nand3_4 _16391_ (.A(_09123_),
    .B(_09130_),
    .C(net498),
    .Y(_09148_));
 sky130_fd_sc_hd__a22oi_4 _16392_ (.A1(net666),
    .A2(_08450_),
    .B1(_08495_),
    .B2(_09148_),
    .Y(_09149_));
 sky130_fd_sc_hd__xnor2_2 _16393_ (.A(net696),
    .B(_09149_),
    .Y(_09150_));
 sky130_fd_sc_hd__nor2_1 _16394_ (.A(_08504_),
    .B(_09148_),
    .Y(_09151_));
 sky130_fd_sc_hd__o22ai_1 _16395_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[38] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[6] ),
    .B2(_08503_),
    .Y(_09152_));
 sky130_fd_sc_hd__a211oi_2 _16396_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(net572),
    .B1(_09152_),
    .C1(_09151_),
    .Y(_09153_));
 sky130_fd_sc_hd__mux2i_4 _16397_ (.A0(_09150_),
    .A1(_09153_),
    .S(net1101),
    .Y(_09154_));
 sky130_fd_sc_hd__inv_1 _16398_ (.A(_09154_),
    .Y(_09155_));
 sky130_fd_sc_hd__maj3_1 _16399_ (.A(_08551_),
    .B(_09119_),
    .C(_09155_),
    .X(_09156_));
 sky130_fd_sc_hd__xnor2_4 _16400_ (.A(_09156_),
    .B(_08510_),
    .Y(_09157_));
 sky130_fd_sc_hd__clkinv_8 _16401_ (.A(net1022),
    .Y(net178));
 sky130_fd_sc_hd__xnor2_2 _16402_ (.A(_08550_),
    .B(_09154_),
    .Y(_09158_));
 sky130_fd_sc_hd__xnor2_4 _16403_ (.A(_09158_),
    .B(_09119_),
    .Y(_09159_));
 sky130_fd_sc_hd__inv_4 _16404_ (.A(_09159_),
    .Y(net177));
 sky130_fd_sc_hd__xnor2_1 _16405_ (.A(_09115_),
    .B(_09116_),
    .Y(_09160_));
 sky130_fd_sc_hd__nor3_2 _16406_ (.A(_08510_),
    .B(_09160_),
    .C(_09158_),
    .Y(_09161_));
 sky130_fd_sc_hd__mux2i_2 _16407_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[520] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[552] ),
    .S(net733),
    .Y(_09162_));
 sky130_fd_sc_hd__mux2i_1 _16408_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[648] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[680] ),
    .S(net733),
    .Y(_09163_));
 sky130_fd_sc_hd__a22oi_1 _16409_ (.A1(net864),
    .A2(_09162_),
    .B1(_09163_),
    .B2(net620),
    .Y(_09164_));
 sky130_fd_sc_hd__mux2i_1 _16410_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[456] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[488] ),
    .S(net733),
    .Y(_09165_));
 sky130_fd_sc_hd__mux2i_2 _16411_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[584] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[616] ),
    .S(net733),
    .Y(_09166_));
 sky130_fd_sc_hd__a22oi_1 _16412_ (.A1(_08593_),
    .A2(_09165_),
    .B1(_09166_),
    .B2(net717),
    .Y(_09167_));
 sky130_fd_sc_hd__mux2i_1 _16413_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[264] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[296] ),
    .S(net733),
    .Y(_09168_));
 sky130_fd_sc_hd__mux2i_1 _16414_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[712] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[744] ),
    .S(net733),
    .Y(_09169_));
 sky130_fd_sc_hd__a22oi_1 _16415_ (.A1(net558),
    .A2(_09168_),
    .B1(_09169_),
    .B2(_08602_),
    .Y(_09170_));
 sky130_fd_sc_hd__mux2i_1 _16416_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[328] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[360] ),
    .S(net733),
    .Y(_09171_));
 sky130_fd_sc_hd__mux2i_1 _16417_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[392] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[424] ),
    .S(net733),
    .Y(_09172_));
 sky130_fd_sc_hd__a22oi_1 _16418_ (.A1(net714),
    .A2(_09171_),
    .B1(_09172_),
    .B2(net567),
    .Y(_09173_));
 sky130_fd_sc_hd__and4_4 _16419_ (.A(_09167_),
    .B(_09173_),
    .C(_09170_),
    .D(_09164_),
    .X(_09174_));
 sky130_fd_sc_hd__mux4_1 _16420_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[136] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[168] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[200] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[232] ),
    .S0(net436),
    .S1(net401),
    .X(_09175_));
 sky130_fd_sc_hd__nand2_1 _16421_ (.A(net396),
    .B(_09175_),
    .Y(_09176_));
 sky130_fd_sc_hd__mux2i_1 _16422_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[72] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[104] ),
    .S(net436),
    .Y(_09177_));
 sky130_fd_sc_hd__a21oi_1 _16423_ (.A1(net436),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[40] ),
    .B1(net401),
    .Y(_09178_));
 sky130_fd_sc_hd__a211o_1 _16424_ (.A1(net401),
    .A2(_09177_),
    .B1(_09178_),
    .C1(net396),
    .X(_09179_));
 sky130_fd_sc_hd__mux4_1 _16425_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[904] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[936] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[968] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1000] ),
    .S0(net938),
    .S1(net1078),
    .X(_09180_));
 sky130_fd_sc_hd__mux4_1 _16426_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[776] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[808] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[840] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[872] ),
    .S0(net938),
    .S1(net1078),
    .X(_09181_));
 sky130_fd_sc_hd__mux2i_4 _16427_ (.A0(_09180_),
    .A1(_09181_),
    .S(_08529_),
    .Y(_09182_));
 sky130_fd_sc_hd__a32oi_4 _16428_ (.A1(_08179_),
    .A2(_09176_),
    .A3(_09179_),
    .B1(_09182_),
    .B2(_08618_),
    .Y(_09183_));
 sky130_fd_sc_hd__nand2_8 _16429_ (.A(_09174_),
    .B(_09183_),
    .Y(_09184_));
 sky130_fd_sc_hd__inv_1 _16430_ (.A(\cs_registers_i.pc_id_i[8] ),
    .Y(_09185_));
 sky130_fd_sc_hd__mux2i_1 _16431_ (.A0(_09184_),
    .A1(_09185_),
    .S(net310),
    .Y(_09186_));
 sky130_fd_sc_hd__a22o_4 _16432_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[8] ),
    .A2(_08368_),
    .B1(_09186_),
    .B2(_08372_),
    .X(_09187_));
 sky130_fd_sc_hd__nand2_1 _16433_ (.A(net1134),
    .B(_09187_),
    .Y(_09188_));
 sky130_fd_sc_hd__nand3_1 _16434_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[40] ),
    .B(_08272_),
    .C(_08377_),
    .Y(_09189_));
 sky130_fd_sc_hd__nand2_1 _16435_ (.A(_09188_),
    .B(_09189_),
    .Y(_09190_));
 sky130_fd_sc_hd__inv_1 _16436_ (.A(_09190_),
    .Y(_09191_));
 sky130_fd_sc_hd__mux4_1 _16437_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[136] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[168] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[200] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[232] ),
    .S0(net373),
    .S1(net1141),
    .X(_09192_));
 sky130_fd_sc_hd__nor2_1 _16438_ (.A(_08481_),
    .B(_09192_),
    .Y(_09193_));
 sky130_fd_sc_hd__mux2_1 _16439_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[40] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[104] ),
    .S(net1141),
    .X(_09194_));
 sky130_fd_sc_hd__a221oi_2 _16440_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[72] ),
    .A2(net324),
    .B1(_09194_),
    .B2(net373),
    .C1(net341),
    .Y(_09195_));
 sky130_fd_sc_hd__mux2i_1 _16441_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[552] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[616] ),
    .S(net349),
    .Y(_09196_));
 sky130_fd_sc_hd__nand2_1 _16442_ (.A(net1201),
    .B(_09196_),
    .Y(_09197_));
 sky130_fd_sc_hd__mux2i_1 _16443_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[680] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[744] ),
    .S(net349),
    .Y(_09198_));
 sky130_fd_sc_hd__mux2i_1 _16444_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[520] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[584] ),
    .S(net349),
    .Y(_09199_));
 sky130_fd_sc_hd__a22oi_2 _16445_ (.A1(net1024),
    .A2(_09198_),
    .B1(_09199_),
    .B2(net650),
    .Y(_09200_));
 sky130_fd_sc_hd__mux2i_1 _16446_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[648] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[712] ),
    .S(net349),
    .Y(_09201_));
 sky130_fd_sc_hd__a21oi_1 _16447_ (.A1(net1013),
    .A2(_09201_),
    .B1(_08679_),
    .Y(_09202_));
 sky130_fd_sc_hd__nand3_4 _16448_ (.A(_09197_),
    .B(_09200_),
    .C(_09202_),
    .Y(_09203_));
 sky130_fd_sc_hd__mux2i_1 _16449_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[808] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[872] ),
    .S(net352),
    .Y(_09204_));
 sky130_fd_sc_hd__mux2i_1 _16450_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[904] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[968] ),
    .S(net351),
    .Y(_09205_));
 sky130_fd_sc_hd__o22ai_2 _16451_ (.A1(net518),
    .A2(_09204_),
    .B1(_09205_),
    .B2(net601),
    .Y(_09206_));
 sky130_fd_sc_hd__mux2i_1 _16452_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[936] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1000] ),
    .S(net351),
    .Y(_09207_));
 sky130_fd_sc_hd__mux2i_1 _16453_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[296] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[360] ),
    .S(net351),
    .Y(_09208_));
 sky130_fd_sc_hd__o22ai_2 _16454_ (.A1(net629),
    .A2(_09207_),
    .B1(_09208_),
    .B2(net759),
    .Y(_09209_));
 sky130_fd_sc_hd__mux2i_1 _16455_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[776] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[840] ),
    .S(net352),
    .Y(_09210_));
 sky130_fd_sc_hd__mux2i_2 _16456_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[392] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[456] ),
    .S(net349),
    .Y(_09211_));
 sky130_fd_sc_hd__o22ai_2 _16457_ (.A1(net508),
    .A2(_09210_),
    .B1(_09211_),
    .B2(net892),
    .Y(_09212_));
 sky130_fd_sc_hd__mux2i_2 _16458_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[424] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[488] ),
    .S(net349),
    .Y(_09213_));
 sky130_fd_sc_hd__mux2i_1 _16459_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[264] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[328] ),
    .S(net351),
    .Y(_09214_));
 sky130_fd_sc_hd__o22ai_2 _16460_ (.A1(net870),
    .A2(_09213_),
    .B1(_09214_),
    .B2(net772),
    .Y(_09215_));
 sky130_fd_sc_hd__nor4_4 _16461_ (.A(_09215_),
    .B(_09209_),
    .C(_09206_),
    .D(_09212_),
    .Y(_09216_));
 sky130_fd_sc_hd__o311a_4 _16462_ (.A1(_08163_),
    .A2(_09193_),
    .A3(_09195_),
    .B1(_09203_),
    .C1(_09216_),
    .X(_09217_));
 sky130_fd_sc_hd__o22ai_1 _16463_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[40] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[8] ),
    .B2(_08503_),
    .Y(_09218_));
 sky130_fd_sc_hd__a221o_1 _16464_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(_09184_),
    .B1(_09217_),
    .B2(_08696_),
    .C1(_09218_),
    .X(_09219_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_913 ();
 sky130_fd_sc_hd__nor2_1 _16466_ (.A(_08436_),
    .B(_09217_),
    .Y(_09221_));
 sky130_fd_sc_hd__a21oi_4 _16467_ (.A1(net814),
    .A2(_08450_),
    .B1(_09221_),
    .Y(_09222_));
 sky130_fd_sc_hd__xnor2_1 _16468_ (.A(net694),
    .B(_09222_),
    .Y(_09223_));
 sky130_fd_sc_hd__nand2_1 _16469_ (.A(net1134),
    .B(_09223_),
    .Y(_09224_));
 sky130_fd_sc_hd__o21ai_2 _16470_ (.A1(net1134),
    .A2(_09219_),
    .B1(_09224_),
    .Y(_09225_));
 sky130_fd_sc_hd__nand2_1 _16471_ (.A(_09191_),
    .B(_09225_),
    .Y(_09226_));
 sky130_fd_sc_hd__nand4_4 _16472_ (.A(_09053_),
    .B(_08752_),
    .C(_09161_),
    .D(_09226_),
    .Y(_09227_));
 sky130_fd_sc_hd__and2_0 _16473_ (.A(_08380_),
    .B(_08509_),
    .X(_09228_));
 sky130_fd_sc_hd__maj3_2 _16474_ (.A(_08550_),
    .B(_09114_),
    .C(_09154_),
    .X(_09229_));
 sky130_fd_sc_hd__or2_0 _16475_ (.A(_08380_),
    .B(_08509_),
    .X(_09230_));
 sky130_fd_sc_hd__o21ai_2 _16476_ (.A1(_09228_),
    .A2(_09229_),
    .B1(_09230_),
    .Y(_09231_));
 sky130_fd_sc_hd__maj3_2 _16477_ (.A(_09231_),
    .B(_09225_),
    .C(_09191_),
    .X(_09232_));
 sky130_fd_sc_hd__nand2_4 _16478_ (.A(_09232_),
    .B(_09227_),
    .Y(_09233_));
 sky130_fd_sc_hd__mux2i_1 _16479_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[809] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[873] ),
    .S(net359),
    .Y(_09234_));
 sky130_fd_sc_hd__mux2i_1 _16480_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[905] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[969] ),
    .S(net359),
    .Y(_09235_));
 sky130_fd_sc_hd__o22ai_1 _16481_ (.A1(net1280),
    .A2(_09234_),
    .B1(_09235_),
    .B2(net934),
    .Y(_09236_));
 sky130_fd_sc_hd__mux2i_1 _16482_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[777] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[841] ),
    .S(net359),
    .Y(_09237_));
 sky130_fd_sc_hd__mux2i_1 _16483_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[937] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1001] ),
    .S(net359),
    .Y(_09238_));
 sky130_fd_sc_hd__o22ai_1 _16484_ (.A1(net506),
    .A2(_09237_),
    .B1(_09238_),
    .B2(_08910_),
    .Y(_09239_));
 sky130_fd_sc_hd__nor2_1 _16485_ (.A(_09236_),
    .B(_09239_),
    .Y(_09240_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_912 ();
 sky130_fd_sc_hd__mux4_1 _16487_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[137] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[169] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[201] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[233] ),
    .S0(net375),
    .S1(net365),
    .X(_09242_));
 sky130_fd_sc_hd__mux2_1 _16488_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[41] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[105] ),
    .S(net365),
    .X(_09243_));
 sky130_fd_sc_hd__a221o_1 _16489_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[73] ),
    .A2(net324),
    .B1(_09243_),
    .B2(net1154),
    .C1(net343),
    .X(_09244_));
 sky130_fd_sc_hd__o211ai_4 _16490_ (.A1(_08481_),
    .A2(_09242_),
    .B1(_09244_),
    .C1(_08731_),
    .Y(_09245_));
 sky130_fd_sc_hd__mux2i_1 _16491_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[297] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[361] ),
    .S(net353),
    .Y(_09246_));
 sky130_fd_sc_hd__mux2i_1 _16492_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[265] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[329] ),
    .S(net353),
    .Y(_09247_));
 sky130_fd_sc_hd__a22oi_1 _16493_ (.A1(net328),
    .A2(_09246_),
    .B1(_09247_),
    .B2(net325),
    .Y(_09248_));
 sky130_fd_sc_hd__mux2i_1 _16494_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[425] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[489] ),
    .S(net353),
    .Y(_09249_));
 sky130_fd_sc_hd__mux2i_1 _16495_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[393] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[457] ),
    .S(net353),
    .Y(_09250_));
 sky130_fd_sc_hd__a22oi_1 _16496_ (.A1(net1024),
    .A2(_09249_),
    .B1(_09250_),
    .B2(net326),
    .Y(_09251_));
 sky130_fd_sc_hd__nand3_2 _16497_ (.A(net700),
    .B(_09248_),
    .C(_09251_),
    .Y(_09252_));
 sky130_fd_sc_hd__mux2i_1 _16498_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[553] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[617] ),
    .S(net353),
    .Y(_09253_));
 sky130_fd_sc_hd__mux2i_1 _16499_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[649] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[713] ),
    .S(net353),
    .Y(_09254_));
 sky130_fd_sc_hd__a22oi_1 _16500_ (.A1(net328),
    .A2(_09253_),
    .B1(_09254_),
    .B2(net1119),
    .Y(_09255_));
 sky130_fd_sc_hd__mux2i_1 _16501_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[521] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[585] ),
    .S(net353),
    .Y(_09256_));
 sky130_fd_sc_hd__mux2i_1 _16502_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[681] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[745] ),
    .S(net353),
    .Y(_09257_));
 sky130_fd_sc_hd__a22oi_1 _16503_ (.A1(net325),
    .A2(_09256_),
    .B1(_09257_),
    .B2(net1024),
    .Y(_09258_));
 sky130_fd_sc_hd__nand3_2 _16504_ (.A(_08462_),
    .B(_09255_),
    .C(_09258_),
    .Y(_09259_));
 sky130_fd_sc_hd__nand4_4 _16505_ (.A(_09240_),
    .B(_09245_),
    .C(_09252_),
    .D(_09259_),
    .Y(_09260_));
 sky130_fd_sc_hd__a22o_4 _16506_ (.A1(net674),
    .A2(_08450_),
    .B1(_09260_),
    .B2(_08495_),
    .X(_09261_));
 sky130_fd_sc_hd__xor2_1 _16507_ (.A(net297),
    .B(_09261_),
    .X(_09262_));
 sky130_fd_sc_hd__mux4_1 _16508_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[777] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[809] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[841] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[873] ),
    .S0(net1311),
    .S1(net406),
    .X(_09263_));
 sky130_fd_sc_hd__nand3b_4 _16509_ (.A_N(net396),
    .B(net1108),
    .C(net384),
    .Y(_09264_));
 sky130_fd_sc_hd__nand3_4 _16510_ (.A(net384),
    .B(net388),
    .C(net396),
    .Y(_09265_));
 sky130_fd_sc_hd__mux4_1 _16511_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[905] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[937] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[969] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1001] ),
    .S0(net1123),
    .S1(net406),
    .X(_09266_));
 sky130_fd_sc_hd__o22ai_1 _16512_ (.A1(_09263_),
    .A2(_09264_),
    .B1(_09265_),
    .B2(_09266_),
    .Y(_09267_));
 sky130_fd_sc_hd__mux4_2 _16513_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[137] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[169] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[201] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[233] ),
    .S0(net438),
    .S1(net402),
    .X(_09268_));
 sky130_fd_sc_hd__mux2i_1 _16514_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[73] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[105] ),
    .S(net435),
    .Y(_09269_));
 sky130_fd_sc_hd__a21oi_1 _16515_ (.A1(net435),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[41] ),
    .B1(net401),
    .Y(_09270_));
 sky130_fd_sc_hd__a211oi_2 _16516_ (.A1(net401),
    .A2(_09269_),
    .B1(_09270_),
    .C1(net398),
    .Y(_09271_));
 sky130_fd_sc_hd__a211oi_4 _16517_ (.A1(net398),
    .A2(_09268_),
    .B1(_09271_),
    .C1(_08821_),
    .Y(_09272_));
 sky130_fd_sc_hd__mux4_1 _16518_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[521] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[553] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[585] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[617] ),
    .S0(net424),
    .S1(net406),
    .X(_09273_));
 sky130_fd_sc_hd__mux4_1 _16519_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[265] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[297] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[329] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[361] ),
    .S0(net424),
    .S1(net406),
    .X(_09274_));
 sky130_fd_sc_hd__nand2b_4 _16520_ (.A_N(net383),
    .B(net1082),
    .Y(_09275_));
 sky130_fd_sc_hd__o22ai_1 _16521_ (.A1(_09032_),
    .A2(_09273_),
    .B1(_09274_),
    .B2(_09275_),
    .Y(_09276_));
 sky130_fd_sc_hd__mux4_1 _16522_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[393] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[425] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[457] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[489] ),
    .S0(net424),
    .S1(net406),
    .X(_09277_));
 sky130_fd_sc_hd__nand3b_1 _16523_ (.A_N(net383),
    .B(net1082),
    .C(net395),
    .Y(_09278_));
 sky130_fd_sc_hd__nand3b_4 _16524_ (.A_N(net388),
    .B(net393),
    .C(net383),
    .Y(_09279_));
 sky130_fd_sc_hd__mux4_1 _16525_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[649] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[681] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[713] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[745] ),
    .S0(net424),
    .S1(net406),
    .X(_09280_));
 sky130_fd_sc_hd__o22ai_1 _16526_ (.A1(_09277_),
    .A2(_09278_),
    .B1(_09279_),
    .B2(_09280_),
    .Y(_09281_));
 sky130_fd_sc_hd__a21o_1 _16527_ (.A1(_08529_),
    .A2(_09276_),
    .B1(_09281_),
    .X(_09282_));
 sky130_fd_sc_hd__or3_4 _16528_ (.A(_09282_),
    .B(_09272_),
    .C(_09267_),
    .X(_09283_));
 sky130_fd_sc_hd__o22ai_1 _16529_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[41] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[9] ),
    .B2(_08503_),
    .Y(_09284_));
 sky130_fd_sc_hd__nor2_1 _16530_ (.A(_08504_),
    .B(_09260_),
    .Y(_09285_));
 sky130_fd_sc_hd__a2111oi_2 _16531_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(_09283_),
    .B1(_09284_),
    .C1(_09285_),
    .D1(_08295_),
    .Y(_09286_));
 sky130_fd_sc_hd__a21oi_1 _16532_ (.A1(_08290_),
    .A2(_09262_),
    .B1(_09286_),
    .Y(_09287_));
 sky130_fd_sc_hd__inv_1 _16533_ (.A(\cs_registers_i.pc_id_i[9] ),
    .Y(_09288_));
 sky130_fd_sc_hd__mux2i_1 _16534_ (.A0(_09283_),
    .A1(_09288_),
    .S(net943),
    .Y(_09289_));
 sky130_fd_sc_hd__a22o_4 _16535_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[9] ),
    .A2(_08368_),
    .B1(_08372_),
    .B2(_09289_),
    .X(_09290_));
 sky130_fd_sc_hd__and3_1 _16536_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[41] ),
    .B(_08272_),
    .C(_08377_),
    .X(_09291_));
 sky130_fd_sc_hd__a21oi_4 _16537_ (.A1(_08290_),
    .A2(_09290_),
    .B1(_09291_),
    .Y(_09292_));
 sky130_fd_sc_hd__xor2_2 _16538_ (.A(_09287_),
    .B(_09292_),
    .X(_09293_));
 sky130_fd_sc_hd__xnor2_4 _16539_ (.A(_09293_),
    .B(_09233_),
    .Y(net180));
 sky130_fd_sc_hd__a21o_2 _16540_ (.A1(_08853_),
    .A2(_09047_),
    .B1(_09052_),
    .X(_09294_));
 sky130_fd_sc_hd__a21oi_4 _16541_ (.A1(_08701_),
    .A2(_09294_),
    .B1(_09048_),
    .Y(_09295_));
 sky130_fd_sc_hd__xnor2_2 _16542_ (.A(_08589_),
    .B(_08751_),
    .Y(_09296_));
 sky130_fd_sc_hd__or4_1 _16543_ (.A(_08510_),
    .B(_09160_),
    .C(_09158_),
    .D(_09296_),
    .X(_09297_));
 sky130_fd_sc_hd__maj3_1 _16544_ (.A(_09115_),
    .B(_09116_),
    .C(net1306),
    .X(_09298_));
 sky130_fd_sc_hd__maj3_1 _16545_ (.A(_08550_),
    .B(_09154_),
    .C(_09298_),
    .X(_09299_));
 sky130_fd_sc_hd__o21ai_2 _16546_ (.A1(_09228_),
    .A2(_09299_),
    .B1(_09230_),
    .Y(_09300_));
 sky130_fd_sc_hd__o21ai_2 _16547_ (.A1(_09295_),
    .A2(_09297_),
    .B1(_09300_),
    .Y(_09301_));
 sky130_fd_sc_hd__xnor2_2 _16548_ (.A(_09190_),
    .B(_09225_),
    .Y(_09302_));
 sky130_fd_sc_hd__xnor2_4 _16549_ (.A(_09302_),
    .B(_09301_),
    .Y(_09303_));
 sky130_fd_sc_hd__inv_12 _16550_ (.A(net1065),
    .Y(net179));
 sky130_fd_sc_hd__nand2_2 _16551_ (.A(net826),
    .B(_08640_),
    .Y(_09304_));
 sky130_fd_sc_hd__or3_1 _16552_ (.A(_08658_),
    .B(_08640_),
    .C(_08643_),
    .X(_09305_));
 sky130_fd_sc_hd__a21oi_1 _16553_ (.A1(_09304_),
    .A2(_09305_),
    .B1(_08439_),
    .Y(_09306_));
 sky130_fd_sc_hd__nand3_1 _16554_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .B(_08439_),
    .C(_08640_),
    .Y(_09307_));
 sky130_fd_sc_hd__nor2_1 _16555_ (.A(_08643_),
    .B(_09307_),
    .Y(_09308_));
 sky130_fd_sc_hd__mux2i_1 _16556_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[299] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[363] ),
    .S(net344),
    .Y(_09309_));
 sky130_fd_sc_hd__mux2i_1 _16557_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[267] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[331] ),
    .S(net344),
    .Y(_09310_));
 sky130_fd_sc_hd__a22oi_1 _16558_ (.A1(net329),
    .A2(_09309_),
    .B1(_09310_),
    .B2(net1044),
    .Y(_09311_));
 sky130_fd_sc_hd__mux2i_1 _16559_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[427] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[491] ),
    .S(net368),
    .Y(_09312_));
 sky130_fd_sc_hd__mux2i_1 _16560_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[395] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[459] ),
    .S(net368),
    .Y(_09313_));
 sky130_fd_sc_hd__a22oi_1 _16561_ (.A1(net1024),
    .A2(_09312_),
    .B1(_09313_),
    .B2(net327),
    .Y(_09314_));
 sky130_fd_sc_hd__and3_1 _16562_ (.A(net707),
    .B(_09311_),
    .C(_09314_),
    .X(_09315_));
 sky130_fd_sc_hd__mux2i_1 _16563_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[555] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[619] ),
    .S(net344),
    .Y(_09316_));
 sky130_fd_sc_hd__mux2i_1 _16564_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[651] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[715] ),
    .S(net344),
    .Y(_09317_));
 sky130_fd_sc_hd__a22oi_1 _16565_ (.A1(net329),
    .A2(_09316_),
    .B1(_09317_),
    .B2(net1474),
    .Y(_09318_));
 sky130_fd_sc_hd__mux2i_1 _16566_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[523] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[587] ),
    .S(net344),
    .Y(_09319_));
 sky130_fd_sc_hd__mux2i_1 _16567_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[683] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[747] ),
    .S(net344),
    .Y(_09320_));
 sky130_fd_sc_hd__a22oi_1 _16568_ (.A1(net1043),
    .A2(_09319_),
    .B1(_09320_),
    .B2(net1024),
    .Y(_09321_));
 sky130_fd_sc_hd__and3_1 _16569_ (.A(_08462_),
    .B(_09318_),
    .C(_09321_),
    .X(_09322_));
 sky130_fd_sc_hd__mux2_1 _16570_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[43] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[107] ),
    .S(net367),
    .X(_09323_));
 sky130_fd_sc_hd__a221oi_4 _16571_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[75] ),
    .A2(net324),
    .B1(_09323_),
    .B2(net1220),
    .C1(net339),
    .Y(_09324_));
 sky130_fd_sc_hd__mux4_1 _16572_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[139] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[171] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[203] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[235] ),
    .S0(net378),
    .S1(net367),
    .X(_09325_));
 sky130_fd_sc_hd__o21ai_4 _16573_ (.A1(_08481_),
    .A2(_09325_),
    .B1(_08731_),
    .Y(_09326_));
 sky130_fd_sc_hd__mux4_1 _16574_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[907] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[939] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[971] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1003] ),
    .S0(net376),
    .S1(net345),
    .X(_09327_));
 sky130_fd_sc_hd__mux4_1 _16575_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[779] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[811] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[843] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[875] ),
    .S0(net376),
    .S1(net345),
    .X(_09328_));
 sky130_fd_sc_hd__a22oi_2 _16576_ (.A1(_08688_),
    .A2(_09327_),
    .B1(_09328_),
    .B2(_08687_),
    .Y(_09329_));
 sky130_fd_sc_hd__o21ai_4 _16577_ (.A1(_09324_),
    .A2(_09326_),
    .B1(_09329_),
    .Y(_09330_));
 sky130_fd_sc_hd__nor3_4 _16578_ (.A(_09322_),
    .B(_09315_),
    .C(_09330_),
    .Y(_09331_));
 sky130_fd_sc_hd__nand2_1 _16579_ (.A(_08495_),
    .B(net307),
    .Y(_09332_));
 sky130_fd_sc_hd__o31ai_4 _16580_ (.A1(_08495_),
    .A2(_09306_),
    .A3(_09308_),
    .B1(_09332_),
    .Y(_09333_));
 sky130_fd_sc_hd__xnor2_4 _16581_ (.A(net297),
    .B(_09333_),
    .Y(_09334_));
 sky130_fd_sc_hd__mux4_2 _16582_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[907] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[939] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[971] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1003] ),
    .S0(net1109),
    .S1(net404),
    .X(_09335_));
 sky130_fd_sc_hd__mux4_2 _16583_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[779] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[811] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[843] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[875] ),
    .S0(net1109),
    .S1(net404),
    .X(_09336_));
 sky130_fd_sc_hd__mux4_1 _16584_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[651] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[683] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[715] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[747] ),
    .S0(net417),
    .S1(net404),
    .X(_09337_));
 sky130_fd_sc_hd__mux4_1 _16585_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[523] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[555] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[587] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[619] ),
    .S0(net417),
    .S1(net404),
    .X(_09338_));
 sky130_fd_sc_hd__a22o_4 _16586_ (.A1(net609),
    .A2(_09337_),
    .B1(_09338_),
    .B2(_08342_),
    .X(_09339_));
 sky130_fd_sc_hd__a221oi_4 _16587_ (.A1(_08324_),
    .A2(_09335_),
    .B1(_09336_),
    .B2(net330),
    .C1(_09339_),
    .Y(_09340_));
 sky130_fd_sc_hd__mux4_1 _16588_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[139] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[171] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[203] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[235] ),
    .S0(net420),
    .S1(net414),
    .X(_09341_));
 sky130_fd_sc_hd__nor2_1 _16589_ (.A(_08529_),
    .B(_09341_),
    .Y(_09342_));
 sky130_fd_sc_hd__mux2_1 _16590_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[75] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[107] ),
    .S(net989),
    .X(_09343_));
 sky130_fd_sc_hd__a221oi_1 _16591_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[43] ),
    .A2(_08321_),
    .B1(_09343_),
    .B2(net1072),
    .C1(net399),
    .Y(_09344_));
 sky130_fd_sc_hd__mux4_2 _16592_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[395] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[427] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[459] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[491] ),
    .S0(net417),
    .S1(net1113),
    .X(_09345_));
 sky130_fd_sc_hd__mux4_1 _16593_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[267] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[299] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[331] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[363] ),
    .S0(net417),
    .S1(net404),
    .X(_09346_));
 sky130_fd_sc_hd__a22oi_4 _16594_ (.A1(net1226),
    .A2(_09345_),
    .B1(_09346_),
    .B2(net530),
    .Y(_09347_));
 sky130_fd_sc_hd__o31a_2 _16595_ (.A1(net975),
    .A2(_09342_),
    .A3(_09344_),
    .B1(_09347_),
    .X(_09348_));
 sky130_fd_sc_hd__mux2i_4 _16596_ (.A0(_09340_),
    .A1(_09348_),
    .S(_08512_),
    .Y(_09349_));
 sky130_fd_sc_hd__o22ai_1 _16597_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[43] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[11] ),
    .B2(_08503_),
    .Y(_09350_));
 sky130_fd_sc_hd__a21oi_1 _16598_ (.A1(_08696_),
    .A2(net307),
    .B1(_09350_),
    .Y(_09351_));
 sky130_fd_sc_hd__o211ai_1 _16599_ (.A1(_08500_),
    .A2(net1187),
    .B1(_09351_),
    .C1(net313),
    .Y(_09352_));
 sky130_fd_sc_hd__a21boi_4 _16600_ (.A1(net1134),
    .A2(_09334_),
    .B1_N(_09352_),
    .Y(_09353_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_911 ();
 sky130_fd_sc_hd__mux2i_1 _16602_ (.A0(_09349_),
    .A1(\cs_registers_i.pc_id_i[11] ),
    .S(_08370_),
    .Y(_09355_));
 sky130_fd_sc_hd__nor2_1 _16603_ (.A(_08307_),
    .B(_09355_),
    .Y(_09356_));
 sky130_fd_sc_hd__a21oi_4 _16604_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[11] ),
    .A2(_08368_),
    .B1(_09356_),
    .Y(_09357_));
 sky130_fd_sc_hd__a21oi_1 _16605_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[43] ),
    .A2(_08377_),
    .B1(_08295_),
    .Y(_09358_));
 sky130_fd_sc_hd__a21oi_4 _16606_ (.A1(_09357_),
    .A2(net1134),
    .B1(_09358_),
    .Y(_09359_));
 sky130_fd_sc_hd__xor2_4 _16607_ (.A(_09353_),
    .B(_09359_),
    .X(_09360_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_910 ();
 sky130_fd_sc_hd__mux4_1 _16609_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[650] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[682] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[714] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[746] ),
    .S0(net417),
    .S1(net404),
    .X(_09362_));
 sky130_fd_sc_hd__mux4_1 _16610_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[522] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[554] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[586] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[618] ),
    .S0(net1135),
    .S1(net404),
    .X(_09363_));
 sky130_fd_sc_hd__a22oi_4 _16611_ (.A1(net609),
    .A2(_09362_),
    .B1(_09363_),
    .B2(_08342_),
    .Y(_09364_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_909 ();
 sky130_fd_sc_hd__mux4_2 _16613_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[906] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[938] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[970] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1002] ),
    .S0(net419),
    .S1(net412),
    .X(_09366_));
 sky130_fd_sc_hd__mux4_1 _16614_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[778] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[810] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[842] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[874] ),
    .S0(net416),
    .S1(net1070),
    .X(_09367_));
 sky130_fd_sc_hd__a22oi_4 _16615_ (.A1(net1226),
    .A2(_09366_),
    .B1(_09367_),
    .B2(net330),
    .Y(_09368_));
 sky130_fd_sc_hd__nand3_2 _16616_ (.A(net386),
    .B(_09364_),
    .C(_09368_),
    .Y(_09369_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_908 ();
 sky130_fd_sc_hd__mux4_1 _16618_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[138] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[170] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[202] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[234] ),
    .S0(net420),
    .S1(net414),
    .X(_09371_));
 sky130_fd_sc_hd__nor2_2 _16619_ (.A(_08529_),
    .B(_09371_),
    .Y(_09372_));
 sky130_fd_sc_hd__mux2_1 _16620_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[74] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[106] ),
    .S(net989),
    .X(_09373_));
 sky130_fd_sc_hd__a221oi_4 _16621_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[42] ),
    .A2(net538),
    .B1(_09373_),
    .B2(net1072),
    .C1(net399),
    .Y(_09374_));
 sky130_fd_sc_hd__mux4_2 _16622_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[394] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[426] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[458] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[490] ),
    .S0(net419),
    .S1(net412),
    .X(_09375_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_907 ();
 sky130_fd_sc_hd__mux4_1 _16624_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[266] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[298] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[330] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[362] ),
    .S0(net416),
    .S1(net1070),
    .X(_09377_));
 sky130_fd_sc_hd__a22oi_4 _16625_ (.A1(net1226),
    .A2(_09375_),
    .B1(_09377_),
    .B2(net330),
    .Y(_09378_));
 sky130_fd_sc_hd__o311ai_4 _16626_ (.A1(net1152),
    .A2(_09372_),
    .A3(_09374_),
    .B1(_09378_),
    .C1(_08512_),
    .Y(_09379_));
 sky130_fd_sc_hd__nand2_8 _16627_ (.A(_09369_),
    .B(_09379_),
    .Y(_09380_));
 sky130_fd_sc_hd__inv_1 _16628_ (.A(\cs_registers_i.pc_id_i[10] ),
    .Y(_09381_));
 sky130_fd_sc_hd__mux2_1 _16629_ (.A0(_09380_),
    .A1(_09381_),
    .S(net943),
    .X(_09382_));
 sky130_fd_sc_hd__nand2_1 _16630_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[10] ),
    .B(_08307_),
    .Y(_09383_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_906 ();
 sky130_fd_sc_hd__o22ai_4 _16632_ (.A1(_08307_),
    .A2(_09382_),
    .B1(_09383_),
    .B2(net944),
    .Y(_09385_));
 sky130_fd_sc_hd__nand2_1 _16633_ (.A(_08295_),
    .B(_09385_),
    .Y(_09386_));
 sky130_fd_sc_hd__nand3_1 _16634_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[42] ),
    .B(_08272_),
    .C(_08377_),
    .Y(_09387_));
 sky130_fd_sc_hd__nand2_1 _16635_ (.A(_09386_),
    .B(_09387_),
    .Y(_09388_));
 sky130_fd_sc_hd__mux4_2 _16636_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[138] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[170] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[202] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[234] ),
    .S0(net379),
    .S1(net371),
    .X(_09389_));
 sky130_fd_sc_hd__mux2_1 _16637_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[42] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[106] ),
    .S(net356),
    .X(_09390_));
 sky130_fd_sc_hd__a221o_1 _16638_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[74] ),
    .A2(net324),
    .B1(_09390_),
    .B2(net1220),
    .C1(net342),
    .X(_09391_));
 sky130_fd_sc_hd__o211ai_4 _16639_ (.A1(_08481_),
    .A2(_09389_),
    .B1(_09391_),
    .C1(_08731_),
    .Y(_09392_));
 sky130_fd_sc_hd__mux2i_1 _16640_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[266] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[330] ),
    .S(net370),
    .Y(_09393_));
 sky130_fd_sc_hd__mux2i_1 _16641_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[906] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[970] ),
    .S(net369),
    .Y(_09394_));
 sky130_fd_sc_hd__o22ai_2 _16642_ (.A1(net808),
    .A2(_09393_),
    .B1(_09394_),
    .B2(net605),
    .Y(_09395_));
 sky130_fd_sc_hd__mux2i_1 _16643_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[938] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1002] ),
    .S(net369),
    .Y(_09396_));
 sky130_fd_sc_hd__mux2i_1 _16644_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[810] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[874] ),
    .S(net370),
    .Y(_09397_));
 sky130_fd_sc_hd__o22ai_2 _16645_ (.A1(net633),
    .A2(_09396_),
    .B1(_09397_),
    .B2(net525),
    .Y(_09398_));
 sky130_fd_sc_hd__mux2i_1 _16646_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[426] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[490] ),
    .S(net369),
    .Y(_09399_));
 sky130_fd_sc_hd__mux2i_1 _16647_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[778] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[842] ),
    .S(net370),
    .Y(_09400_));
 sky130_fd_sc_hd__o22ai_2 _16648_ (.A1(net866),
    .A2(_09399_),
    .B1(_09400_),
    .B2(net504),
    .Y(_09401_));
 sky130_fd_sc_hd__mux2i_1 _16649_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[298] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[362] ),
    .S(net370),
    .Y(_09402_));
 sky130_fd_sc_hd__mux2i_1 _16650_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[394] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[458] ),
    .S(net369),
    .Y(_09403_));
 sky130_fd_sc_hd__o22ai_2 _16651_ (.A1(net764),
    .A2(_09402_),
    .B1(_09403_),
    .B2(net895),
    .Y(_09404_));
 sky130_fd_sc_hd__nor4_4 _16652_ (.A(_09395_),
    .B(_09398_),
    .C(_09401_),
    .D(_09404_),
    .Y(_09405_));
 sky130_fd_sc_hd__mux2i_1 _16653_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[554] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[618] ),
    .S(net344),
    .Y(_09406_));
 sky130_fd_sc_hd__mux2i_1 _16654_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[650] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[714] ),
    .S(net344),
    .Y(_09407_));
 sky130_fd_sc_hd__a22oi_2 _16655_ (.A1(net1201),
    .A2(_09406_),
    .B1(_09407_),
    .B2(net1013),
    .Y(_09408_));
 sky130_fd_sc_hd__mux2i_1 _16656_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[522] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[586] ),
    .S(net344),
    .Y(_09409_));
 sky130_fd_sc_hd__mux2i_1 _16657_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[682] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[746] ),
    .S(net344),
    .Y(_09410_));
 sky130_fd_sc_hd__a22oi_2 _16658_ (.A1(net650),
    .A2(_09409_),
    .B1(_09410_),
    .B2(net1153),
    .Y(_09411_));
 sky130_fd_sc_hd__nand3_4 _16659_ (.A(_08462_),
    .B(_09408_),
    .C(_09411_),
    .Y(_09412_));
 sky130_fd_sc_hd__nand3_4 _16660_ (.A(_09392_),
    .B(_09412_),
    .C(net1079),
    .Y(_09413_));
 sky130_fd_sc_hd__a22oi_4 _16661_ (.A1(net919),
    .A2(_08450_),
    .B1(_08495_),
    .B2(_09413_),
    .Y(_09414_));
 sky130_fd_sc_hd__xnor2_2 _16662_ (.A(net694),
    .B(_09414_),
    .Y(_09415_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_905 ();
 sky130_fd_sc_hd__nor2_1 _16664_ (.A(_08504_),
    .B(_09413_),
    .Y(_09417_));
 sky130_fd_sc_hd__o22ai_1 _16665_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[42] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[10] ),
    .B2(_08503_),
    .Y(_09418_));
 sky130_fd_sc_hd__a211oi_1 _16666_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(_09380_),
    .B1(_09417_),
    .C1(_09418_),
    .Y(_09419_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_904 ();
 sky130_fd_sc_hd__mux2i_4 _16668_ (.A0(_09415_),
    .A1(_09419_),
    .S(net1105),
    .Y(_09421_));
 sky130_fd_sc_hd__xnor2_2 _16669_ (.A(_09388_),
    .B(_09421_),
    .Y(_09422_));
 sky130_fd_sc_hd__nor2_2 _16670_ (.A(_09293_),
    .B(_09422_),
    .Y(_09423_));
 sky130_fd_sc_hd__a211oi_2 _16671_ (.A1(_08295_),
    .A2(_09262_),
    .B1(_09286_),
    .C1(_09292_),
    .Y(_09424_));
 sky130_fd_sc_hd__maj3_2 _16672_ (.A(_09424_),
    .B(_09388_),
    .C(_09421_),
    .X(_09425_));
 sky130_fd_sc_hd__a21oi_4 _16673_ (.A1(_09423_),
    .A2(_09233_),
    .B1(_09425_),
    .Y(_09426_));
 sky130_fd_sc_hd__xor2_4 _16674_ (.A(_09360_),
    .B(_09426_),
    .X(_09427_));
 sky130_fd_sc_hd__inv_4 _16675_ (.A(net1590),
    .Y(net152));
 sky130_fd_sc_hd__nand2b_1 _16676_ (.A_N(_09287_),
    .B(_09292_),
    .Y(_09428_));
 sky130_fd_sc_hd__a21oi_2 _16677_ (.A1(_09233_),
    .A2(_09428_),
    .B1(_09424_),
    .Y(_09429_));
 sky130_fd_sc_hd__xor2_4 _16678_ (.A(_09422_),
    .B(_09429_),
    .X(net151));
 sky130_fd_sc_hd__mux4_1 _16679_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[909] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[941] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[973] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1005] ),
    .S0(net1123),
    .S1(net401),
    .X(_09430_));
 sky130_fd_sc_hd__mux4_1 _16680_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[781] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[813] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[845] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[877] ),
    .S0(net1123),
    .S1(net401),
    .X(_09431_));
 sky130_fd_sc_hd__o22ai_1 _16681_ (.A1(_09265_),
    .A2(_09430_),
    .B1(_09431_),
    .B2(_09264_),
    .Y(_09432_));
 sky130_fd_sc_hd__mux4_1 _16682_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[141] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[173] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[205] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[237] ),
    .S0(net435),
    .S1(net402),
    .X(_09433_));
 sky130_fd_sc_hd__mux2i_1 _16683_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[77] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[109] ),
    .S(net434),
    .Y(_09434_));
 sky130_fd_sc_hd__a21oi_1 _16684_ (.A1(net434),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[45] ),
    .B1(net401),
    .Y(_09435_));
 sky130_fd_sc_hd__a211oi_1 _16685_ (.A1(net401),
    .A2(_09434_),
    .B1(_09435_),
    .C1(net396),
    .Y(_09436_));
 sky130_fd_sc_hd__a211oi_2 _16686_ (.A1(net396),
    .A2(_09433_),
    .B1(_09436_),
    .C1(_08821_),
    .Y(_09437_));
 sky130_fd_sc_hd__mux4_4 _16687_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[525] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[557] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[589] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[621] ),
    .S0(net421),
    .S1(net1185),
    .X(_09438_));
 sky130_fd_sc_hd__mux4_1 _16688_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[269] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[301] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[333] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[365] ),
    .S0(net429),
    .S1(net1078),
    .X(_09439_));
 sky130_fd_sc_hd__o22ai_4 _16689_ (.A1(_09032_),
    .A2(_09438_),
    .B1(_09439_),
    .B2(_09275_),
    .Y(_09440_));
 sky130_fd_sc_hd__mux4_4 _16690_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[397] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[429] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[461] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[493] ),
    .S0(net428),
    .S1(net1078),
    .X(_09441_));
 sky130_fd_sc_hd__mux4_4 _16691_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[653] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[685] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[717] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[749] ),
    .S0(net1283),
    .S1(net1078),
    .X(_09442_));
 sky130_fd_sc_hd__o22ai_2 _16692_ (.A1(_09278_),
    .A2(_09441_),
    .B1(_09442_),
    .B2(_09279_),
    .Y(_09443_));
 sky130_fd_sc_hd__a21o_1 _16693_ (.A1(_09440_),
    .A2(_08529_),
    .B1(_09443_),
    .X(_09444_));
 sky130_fd_sc_hd__or3_4 _16694_ (.A(_09444_),
    .B(_09437_),
    .C(_09432_),
    .X(_09445_));
 sky130_fd_sc_hd__nor2_4 _16695_ (.A(net310),
    .B(net849),
    .Y(_09446_));
 sky130_fd_sc_hd__a21oi_2 _16696_ (.A1(\cs_registers_i.pc_id_i[13] ),
    .A2(net310),
    .B1(_09446_),
    .Y(_09447_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_903 ();
 sky130_fd_sc_hd__nand2_1 _16698_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[13] ),
    .B(_08368_),
    .Y(_09449_));
 sky130_fd_sc_hd__o21ai_4 _16699_ (.A1(net1116),
    .A2(_09447_),
    .B1(_09449_),
    .Y(_09450_));
 sky130_fd_sc_hd__and3_1 _16700_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[45] ),
    .B(_08272_),
    .C(_08377_),
    .X(_09451_));
 sky130_fd_sc_hd__a21o_1 _16701_ (.A1(_09450_),
    .A2(_08290_),
    .B1(_09451_),
    .X(_09452_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_901 ();
 sky130_fd_sc_hd__and2_4 _16704_ (.A(_08439_),
    .B(_08643_),
    .X(_09455_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_900 ();
 sky130_fd_sc_hd__or2_2 _16706_ (.A(_09455_),
    .B(_09304_),
    .X(_09457_));
 sky130_fd_sc_hd__nor3_2 _16707_ (.A(_08439_),
    .B(_08640_),
    .C(_08643_),
    .Y(_09458_));
 sky130_fd_sc_hd__o21ai_1 _16708_ (.A1(_09455_),
    .A2(_09458_),
    .B1(net445),
    .Y(_09459_));
 sky130_fd_sc_hd__mux2i_1 _16709_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[269] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[333] ),
    .S(net1093),
    .Y(_09460_));
 sky130_fd_sc_hd__mux2i_1 _16710_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[301] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[365] ),
    .S(net1093),
    .Y(_09461_));
 sky130_fd_sc_hd__a22oi_2 _16711_ (.A1(net325),
    .A2(_09460_),
    .B1(_09461_),
    .B2(net1201),
    .Y(_09462_));
 sky130_fd_sc_hd__mux2i_1 _16712_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[397] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[461] ),
    .S(net351),
    .Y(_09463_));
 sky130_fd_sc_hd__mux2i_1 _16713_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[429] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[493] ),
    .S(net351),
    .Y(_09464_));
 sky130_fd_sc_hd__a22oi_2 _16714_ (.A1(net1119),
    .A2(_09463_),
    .B1(_09464_),
    .B2(net1153),
    .Y(_09465_));
 sky130_fd_sc_hd__nand3_4 _16715_ (.A(net705),
    .B(_09462_),
    .C(_09465_),
    .Y(_09466_));
 sky130_fd_sc_hd__mux2i_1 _16716_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[557] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[621] ),
    .S(net350),
    .Y(_09467_));
 sky130_fd_sc_hd__mux2i_1 _16717_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[653] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[717] ),
    .S(net350),
    .Y(_09468_));
 sky130_fd_sc_hd__a22oi_2 _16718_ (.A1(net1201),
    .A2(_09467_),
    .B1(_09468_),
    .B2(net1013),
    .Y(_09469_));
 sky130_fd_sc_hd__mux2i_1 _16719_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[525] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[589] ),
    .S(net350),
    .Y(_09470_));
 sky130_fd_sc_hd__mux2i_1 _16720_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[685] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[749] ),
    .S(net350),
    .Y(_09471_));
 sky130_fd_sc_hd__a22oi_2 _16721_ (.A1(net325),
    .A2(_09470_),
    .B1(_09471_),
    .B2(net1153),
    .Y(_09472_));
 sky130_fd_sc_hd__nand3_4 _16722_ (.A(net698),
    .B(_09469_),
    .C(_09472_),
    .Y(_09473_));
 sky130_fd_sc_hd__mux2_1 _16723_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[45] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[109] ),
    .S(net1141),
    .X(_09474_));
 sky130_fd_sc_hd__a221o_1 _16724_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[77] ),
    .A2(net324),
    .B1(_09474_),
    .B2(net983),
    .C1(net340),
    .X(_09475_));
 sky130_fd_sc_hd__mux4_1 _16725_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[141] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[173] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[205] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[237] ),
    .S0(net374),
    .S1(net1077),
    .X(_09476_));
 sky130_fd_sc_hd__nand2b_1 _16726_ (.A_N(_09476_),
    .B(net341),
    .Y(_09477_));
 sky130_fd_sc_hd__mux4_1 _16727_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[909] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[941] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[973] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1005] ),
    .S0(net373),
    .S1(net362),
    .X(_09478_));
 sky130_fd_sc_hd__mux4_1 _16728_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[781] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[813] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[845] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[877] ),
    .S0(net373),
    .S1(net362),
    .X(_09479_));
 sky130_fd_sc_hd__a22o_1 _16729_ (.A1(_08688_),
    .A2(_09478_),
    .B1(_09479_),
    .B2(_08687_),
    .X(_09480_));
 sky130_fd_sc_hd__a31oi_4 _16730_ (.A1(_08731_),
    .A2(_09475_),
    .A3(_09477_),
    .B1(_09480_),
    .Y(_09481_));
 sky130_fd_sc_hd__nand3_4 _16731_ (.A(_09466_),
    .B(_09473_),
    .C(_09481_),
    .Y(_09482_));
 sky130_fd_sc_hd__nor2_2 _16732_ (.A(_08436_),
    .B(_09482_),
    .Y(_09483_));
 sky130_fd_sc_hd__a31oi_4 _16733_ (.A1(_08436_),
    .A2(_09457_),
    .A3(_09459_),
    .B1(_09483_),
    .Y(_09484_));
 sky130_fd_sc_hd__xor2_1 _16734_ (.A(net296),
    .B(_09484_),
    .X(_09485_));
 sky130_fd_sc_hd__and3_2 _16735_ (.A(_09466_),
    .B(_09473_),
    .C(_09481_),
    .X(_09486_));
 sky130_fd_sc_hd__o22ai_1 _16736_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[45] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[13] ),
    .B2(_08503_),
    .Y(_09487_));
 sky130_fd_sc_hd__a221o_1 _16737_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(net833),
    .B1(_09486_),
    .B2(_08696_),
    .C1(_09487_),
    .X(_09488_));
 sky130_fd_sc_hd__nor2_1 _16738_ (.A(net1134),
    .B(_09488_),
    .Y(_09489_));
 sky130_fd_sc_hd__a21oi_2 _16739_ (.A1(net1134),
    .A2(_09485_),
    .B1(_09489_),
    .Y(_09490_));
 sky130_fd_sc_hd__xor2_2 _16740_ (.A(_09490_),
    .B(_09452_),
    .X(_09491_));
 sky130_fd_sc_hd__inv_2 _16741_ (.A(_09491_),
    .Y(_09492_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_899 ();
 sky130_fd_sc_hd__or2_2 _16743_ (.A(_09455_),
    .B(_09458_),
    .X(_09494_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_898 ();
 sky130_fd_sc_hd__nor2_2 _16745_ (.A(_09455_),
    .B(_09304_),
    .Y(_09496_));
 sky130_fd_sc_hd__a21oi_1 _16746_ (.A1(net491),
    .A2(_09494_),
    .B1(_09496_),
    .Y(_09497_));
 sky130_fd_sc_hd__mux2i_1 _16747_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[556] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[620] ),
    .S(net354),
    .Y(_09498_));
 sky130_fd_sc_hd__nand2_1 _16748_ (.A(net328),
    .B(_09498_),
    .Y(_09499_));
 sky130_fd_sc_hd__mux2i_1 _16749_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[684] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[748] ),
    .S(net353),
    .Y(_09500_));
 sky130_fd_sc_hd__mux2i_1 _16750_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[524] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[588] ),
    .S(net354),
    .Y(_09501_));
 sky130_fd_sc_hd__a22oi_1 _16751_ (.A1(net1153),
    .A2(_09500_),
    .B1(_09501_),
    .B2(net325),
    .Y(_09502_));
 sky130_fd_sc_hd__mux2i_1 _16752_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[652] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[716] ),
    .S(net353),
    .Y(_09503_));
 sky130_fd_sc_hd__a21oi_1 _16753_ (.A1(net1014),
    .A2(_09503_),
    .B1(_08679_),
    .Y(_09504_));
 sky130_fd_sc_hd__and3_1 _16754_ (.A(_09499_),
    .B(_09502_),
    .C(_09504_),
    .X(_09505_));
 sky130_fd_sc_hd__mux2i_1 _16755_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[300] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[364] ),
    .S(net355),
    .Y(_09506_));
 sky130_fd_sc_hd__mux2i_1 _16756_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[268] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[332] ),
    .S(net355),
    .Y(_09507_));
 sky130_fd_sc_hd__o22ai_1 _16757_ (.A1(_09060_),
    .A2(_09506_),
    .B1(_09507_),
    .B2(net772),
    .Y(_09508_));
 sky130_fd_sc_hd__mux2i_1 _16758_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[428] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[492] ),
    .S(net355),
    .Y(_09509_));
 sky130_fd_sc_hd__mux2i_1 _16759_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[812] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[876] ),
    .S(net355),
    .Y(_09510_));
 sky130_fd_sc_hd__o22ai_1 _16760_ (.A1(_08469_),
    .A2(_09509_),
    .B1(_09510_),
    .B2(net517),
    .Y(_09511_));
 sky130_fd_sc_hd__mux2i_1 _16761_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[396] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[460] ),
    .S(net355),
    .Y(_09512_));
 sky130_fd_sc_hd__mux2i_1 _16762_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[908] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[972] ),
    .S(net355),
    .Y(_09513_));
 sky130_fd_sc_hd__o22ai_1 _16763_ (.A1(_08474_),
    .A2(_09512_),
    .B1(_09513_),
    .B2(_08901_),
    .Y(_09514_));
 sky130_fd_sc_hd__mux2i_1 _16764_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[940] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1004] ),
    .S(net355),
    .Y(_09515_));
 sky130_fd_sc_hd__mux2i_1 _16765_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[780] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[844] ),
    .S(net355),
    .Y(_09516_));
 sky130_fd_sc_hd__o22ai_1 _16766_ (.A1(_08910_),
    .A2(_09515_),
    .B1(_09516_),
    .B2(net507),
    .Y(_09517_));
 sky130_fd_sc_hd__or4_4 _16767_ (.A(_09508_),
    .B(_09511_),
    .C(_09514_),
    .D(_09517_),
    .X(_09518_));
 sky130_fd_sc_hd__mux4_1 _16768_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[140] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[172] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[204] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[236] ),
    .S0(net1154),
    .S1(net1120),
    .X(_09519_));
 sky130_fd_sc_hd__nor2_1 _16769_ (.A(_08481_),
    .B(_09519_),
    .Y(_09520_));
 sky130_fd_sc_hd__mux2_1 _16770_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[44] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[108] ),
    .S(net1120),
    .X(_09521_));
 sky130_fd_sc_hd__a221oi_2 _16771_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[76] ),
    .A2(net324),
    .B1(_09521_),
    .B2(net983),
    .C1(net343),
    .Y(_09522_));
 sky130_fd_sc_hd__nor3_4 _16772_ (.A(_08163_),
    .B(_09520_),
    .C(_09522_),
    .Y(_09523_));
 sky130_fd_sc_hd__or3_4 _16773_ (.A(_09505_),
    .B(_09518_),
    .C(_09523_),
    .X(_09524_));
 sky130_fd_sc_hd__nand2_1 _16774_ (.A(_08495_),
    .B(_09524_),
    .Y(_09525_));
 sky130_fd_sc_hd__o21ai_2 _16775_ (.A1(_08495_),
    .A2(_09497_),
    .B1(_09525_),
    .Y(_09526_));
 sky130_fd_sc_hd__xor2_2 _16776_ (.A(net297),
    .B(_09526_),
    .X(_09527_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_897 ();
 sky130_fd_sc_hd__mux2_1 _16778_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[140] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[172] ),
    .S(net753),
    .X(_09529_));
 sky130_fd_sc_hd__nor2b_4 _16779_ (.A(net397),
    .B_N(net1084),
    .Y(_09530_));
 sky130_fd_sc_hd__a22oi_2 _16780_ (.A1(net398),
    .A2(_09529_),
    .B1(_09530_),
    .B2(\gen_regfile_ff.register_file_i.rf_reg[44] ),
    .Y(_09531_));
 sky130_fd_sc_hd__mux4_1 _16781_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[76] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[108] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[204] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[236] ),
    .S0(net753),
    .S1(net398),
    .X(_09532_));
 sky130_fd_sc_hd__nand2_1 _16782_ (.A(net403),
    .B(_09532_),
    .Y(_09533_));
 sky130_fd_sc_hd__o211ai_4 _16783_ (.A1(net402),
    .A2(_09531_),
    .B1(_09533_),
    .C1(_08179_),
    .Y(_09534_));
 sky130_fd_sc_hd__mux2_1 _16784_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[908] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[940] ),
    .S(net1016),
    .X(_09535_));
 sky130_fd_sc_hd__nand2b_1 _16785_ (.A_N(\gen_regfile_ff.register_file_i.rf_reg[1004] ),
    .B(net799),
    .Y(_09536_));
 sky130_fd_sc_hd__o221ai_2 _16786_ (.A1(net799),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[972] ),
    .B1(_09535_),
    .B2(net405),
    .C1(_09536_),
    .Y(_09537_));
 sky130_fd_sc_hd__mux2_1 _16787_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[780] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[812] ),
    .S(net427),
    .X(_09538_));
 sky130_fd_sc_hd__mux2_1 _16788_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[844] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[876] ),
    .S(net865),
    .X(_09539_));
 sky130_fd_sc_hd__o211ai_2 _16789_ (.A1(net405),
    .A2(_09538_),
    .B1(_09539_),
    .C1(_08529_),
    .Y(_09540_));
 sky130_fd_sc_hd__a221oi_2 _16790_ (.A1(net323),
    .A2(_09535_),
    .B1(_09538_),
    .B2(_08187_),
    .C1(_08809_),
    .Y(_09541_));
 sky130_fd_sc_hd__o211ai_4 _16791_ (.A1(_08529_),
    .A2(_09537_),
    .B1(_09540_),
    .C1(_09541_),
    .Y(_09542_));
 sky130_fd_sc_hd__nand3b_4 _16792_ (.A_N(net383),
    .B(net1108),
    .C(net406),
    .Y(_09543_));
 sky130_fd_sc_hd__mux4_1 _16793_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[332] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[364] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[460] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[492] ),
    .S0(net1016),
    .S1(net393),
    .X(_09544_));
 sky130_fd_sc_hd__mux4_1 _16794_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[268] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[300] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[396] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[428] ),
    .S0(net1016),
    .S1(net393),
    .X(_09545_));
 sky130_fd_sc_hd__or3b_4 _16795_ (.A(net383),
    .B(net1083),
    .C_N(net388),
    .X(_09546_));
 sky130_fd_sc_hd__o22ai_2 _16796_ (.A1(_09543_),
    .A2(_09544_),
    .B1(_09545_),
    .B2(_09546_),
    .Y(_09547_));
 sky130_fd_sc_hd__mux4_1 _16797_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[652] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[684] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[716] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[748] ),
    .S0(net424),
    .S1(net1083),
    .X(_09548_));
 sky130_fd_sc_hd__mux4_1 _16798_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[524] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[556] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[588] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[620] ),
    .S0(net1016),
    .S1(net1204),
    .X(_09549_));
 sky130_fd_sc_hd__or3b_4 _16799_ (.A(net1108),
    .B(net393),
    .C_N(net383),
    .X(_09550_));
 sky130_fd_sc_hd__o22ai_1 _16800_ (.A1(_09279_),
    .A2(_09548_),
    .B1(_09549_),
    .B2(_09550_),
    .Y(_09551_));
 sky130_fd_sc_hd__nor2_2 _16801_ (.A(_09547_),
    .B(_09551_),
    .Y(_09552_));
 sky130_fd_sc_hd__nand3_4 _16802_ (.A(_09534_),
    .B(_09542_),
    .C(_09552_),
    .Y(_09553_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_896 ();
 sky130_fd_sc_hd__o22ai_1 _16804_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[44] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[12] ),
    .B2(_08503_),
    .Y(_09555_));
 sky130_fd_sc_hd__nor2_1 _16805_ (.A(_08504_),
    .B(_09524_),
    .Y(_09556_));
 sky130_fd_sc_hd__a2111oi_2 _16806_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(_09553_),
    .B1(_09555_),
    .C1(_09556_),
    .D1(net1134),
    .Y(_09557_));
 sky130_fd_sc_hd__a21oi_4 _16807_ (.A1(net1134),
    .A2(_09527_),
    .B1(_09557_),
    .Y(_09558_));
 sky130_fd_sc_hd__nor2_1 _16808_ (.A(_08370_),
    .B(_09553_),
    .Y(_09559_));
 sky130_fd_sc_hd__a21oi_1 _16809_ (.A1(\cs_registers_i.pc_id_i[12] ),
    .A2(_08370_),
    .B1(_09559_),
    .Y(_09560_));
 sky130_fd_sc_hd__nand2_1 _16810_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[12] ),
    .B(_08368_),
    .Y(_09561_));
 sky130_fd_sc_hd__o21ai_4 _16811_ (.A1(net1115),
    .A2(_09560_),
    .B1(_09561_),
    .Y(_09562_));
 sky130_fd_sc_hd__nand2_1 _16812_ (.A(net1134),
    .B(_09562_),
    .Y(_09563_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_895 ();
 sky130_fd_sc_hd__nand3_1 _16814_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[44] ),
    .B(_08272_),
    .C(_08377_),
    .Y(_09565_));
 sky130_fd_sc_hd__nand2_2 _16815_ (.A(_09563_),
    .B(_09565_),
    .Y(_09566_));
 sky130_fd_sc_hd__xnor2_4 _16816_ (.A(_09558_),
    .B(_09566_),
    .Y(_09567_));
 sky130_fd_sc_hd__nand2_1 _16817_ (.A(_09360_),
    .B(_09423_),
    .Y(_09568_));
 sky130_fd_sc_hd__a21o_4 _16818_ (.A1(_09232_),
    .A2(_09227_),
    .B1(_09568_),
    .X(_09569_));
 sky130_fd_sc_hd__and2_1 _16819_ (.A(_09353_),
    .B(_09359_),
    .X(_09570_));
 sky130_fd_sc_hd__a21oi_2 _16820_ (.A1(_09558_),
    .A2(_09566_),
    .B1(_09570_),
    .Y(_09571_));
 sky130_fd_sc_hd__o21ai_0 _16821_ (.A1(_09353_),
    .A2(_09359_),
    .B1(_09425_),
    .Y(_09572_));
 sky130_fd_sc_hd__nor2_1 _16822_ (.A(_09558_),
    .B(_09566_),
    .Y(_09573_));
 sky130_fd_sc_hd__a21o_1 _16823_ (.A1(_09571_),
    .A2(_09572_),
    .B1(_09573_),
    .X(_09574_));
 sky130_fd_sc_hd__o21ai_2 _16824_ (.A1(_09567_),
    .A2(_09569_),
    .B1(_09574_),
    .Y(_09575_));
 sky130_fd_sc_hd__xnor2_4 _16825_ (.A(_09575_),
    .B(_09492_),
    .Y(net154));
 sky130_fd_sc_hd__nor2_1 _16826_ (.A(_09353_),
    .B(_09359_),
    .Y(_09576_));
 sky130_fd_sc_hd__o21bai_4 _16827_ (.A1(_09576_),
    .A2(_09426_),
    .B1_N(_09570_),
    .Y(_09577_));
 sky130_fd_sc_hd__xnor2_4 _16828_ (.A(_09577_),
    .B(_09567_),
    .Y(net153));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_894 ();
 sky130_fd_sc_hd__a21oi_1 _16830_ (.A1(net443),
    .A2(_09494_),
    .B1(_09496_),
    .Y(_09579_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_893 ();
 sky130_fd_sc_hd__mux4_1 _16832_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[142] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[174] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[206] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[238] ),
    .S0(net1476),
    .S1(net988),
    .X(_09581_));
 sky130_fd_sc_hd__mux2_1 _16833_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[46] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[110] ),
    .S(net366),
    .X(_09582_));
 sky130_fd_sc_hd__a221o_1 _16834_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[78] ),
    .A2(net324),
    .B1(_09582_),
    .B2(net1476),
    .C1(net342),
    .X(_09583_));
 sky130_fd_sc_hd__o211ai_4 _16835_ (.A1(_08481_),
    .A2(_09581_),
    .B1(_09583_),
    .C1(_08731_),
    .Y(_09584_));
 sky130_fd_sc_hd__mux4_1 _16836_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[910] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[942] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[974] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1006] ),
    .S0(net379),
    .S1(net371),
    .X(_09585_));
 sky130_fd_sc_hd__nand2_1 _16837_ (.A(net334),
    .B(_09585_),
    .Y(_09586_));
 sky130_fd_sc_hd__mux4_1 _16838_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[398] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[430] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[462] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[494] ),
    .S0(net379),
    .S1(net371),
    .X(_09587_));
 sky130_fd_sc_hd__nand2_1 _16839_ (.A(_08161_),
    .B(_09587_),
    .Y(_09588_));
 sky130_fd_sc_hd__a21o_2 _16840_ (.A1(_09586_),
    .A2(_09588_),
    .B1(_09075_),
    .X(_09589_));
 sky130_fd_sc_hd__mux2i_2 _16841_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[782] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[846] ),
    .S(net370),
    .Y(_09590_));
 sky130_fd_sc_hd__mux2i_2 _16842_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[814] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[878] ),
    .S(net370),
    .Y(_09591_));
 sky130_fd_sc_hd__o22ai_4 _16843_ (.A1(net503),
    .A2(_09590_),
    .B1(_09591_),
    .B2(net524),
    .Y(_09592_));
 sky130_fd_sc_hd__mux2i_1 _16844_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[302] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[366] ),
    .S(net1142),
    .Y(_09593_));
 sky130_fd_sc_hd__nor2_1 _16845_ (.A(_09060_),
    .B(_09593_),
    .Y(_09594_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_892 ();
 sky130_fd_sc_hd__mux2i_1 _16847_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[270] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[334] ),
    .S(net1142),
    .Y(_09596_));
 sky130_fd_sc_hd__nor2_1 _16848_ (.A(net883),
    .B(_09596_),
    .Y(_09597_));
 sky130_fd_sc_hd__nor3_2 _16849_ (.A(_09592_),
    .B(_09594_),
    .C(_09597_),
    .Y(_09598_));
 sky130_fd_sc_hd__mux2i_1 _16850_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[558] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[622] ),
    .S(net988),
    .Y(_09599_));
 sky130_fd_sc_hd__mux2i_1 _16851_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[654] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[718] ),
    .S(net988),
    .Y(_09600_));
 sky130_fd_sc_hd__a22oi_1 _16852_ (.A1(net328),
    .A2(_09599_),
    .B1(_09600_),
    .B2(net592),
    .Y(_09601_));
 sky130_fd_sc_hd__mux2i_1 _16853_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[526] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[590] ),
    .S(net364),
    .Y(_09602_));
 sky130_fd_sc_hd__mux2i_1 _16854_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[686] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[750] ),
    .S(net988),
    .Y(_09603_));
 sky130_fd_sc_hd__a22oi_1 _16855_ (.A1(net325),
    .A2(_09602_),
    .B1(_09603_),
    .B2(net1153),
    .Y(_09604_));
 sky130_fd_sc_hd__nand3_1 _16856_ (.A(net698),
    .B(_09601_),
    .C(_09604_),
    .Y(_09605_));
 sky130_fd_sc_hd__nand4_4 _16857_ (.A(_09598_),
    .B(_09589_),
    .C(_09584_),
    .D(_09605_),
    .Y(_09606_));
 sky130_fd_sc_hd__nand2_1 _16858_ (.A(_08495_),
    .B(_09606_),
    .Y(_09607_));
 sky130_fd_sc_hd__o21ai_2 _16859_ (.A1(_08495_),
    .A2(_09579_),
    .B1(_09607_),
    .Y(_09608_));
 sky130_fd_sc_hd__xor2_2 _16860_ (.A(net296),
    .B(_09608_),
    .X(_09609_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_891 ();
 sky130_fd_sc_hd__mux4_1 _16862_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[910] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[942] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[974] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1006] ),
    .S0(net419),
    .S1(net412),
    .X(_09611_));
 sky130_fd_sc_hd__mux4_1 _16863_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[782] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[814] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[846] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[878] ),
    .S0(net420),
    .S1(net1009),
    .X(_09612_));
 sky130_fd_sc_hd__mux2_2 _16864_ (.A0(_09611_),
    .A1(_09612_),
    .S(_08529_),
    .X(_09613_));
 sky130_fd_sc_hd__nand2_1 _16865_ (.A(net1140),
    .B(_09613_),
    .Y(_09614_));
 sky130_fd_sc_hd__mux2i_1 _16866_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[718] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[750] ),
    .S(net962),
    .Y(_09615_));
 sky130_fd_sc_hd__mux2i_1 _16867_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[654] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[686] ),
    .S(net962),
    .Y(_09616_));
 sky130_fd_sc_hd__a22oi_2 _16868_ (.A1(_08803_),
    .A2(_09615_),
    .B1(_09616_),
    .B2(net1149),
    .Y(_09617_));
 sky130_fd_sc_hd__mux2i_1 _16869_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[590] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[622] ),
    .S(net1111),
    .Y(_09618_));
 sky130_fd_sc_hd__mux2i_1 _16870_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[526] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[558] ),
    .S(net962),
    .Y(_09619_));
 sky130_fd_sc_hd__a22oi_1 _16871_ (.A1(net613),
    .A2(_09618_),
    .B1(_09619_),
    .B2(net649),
    .Y(_09620_));
 sky130_fd_sc_hd__nand3_1 _16872_ (.A(_08309_),
    .B(_09617_),
    .C(_09620_),
    .Y(_09621_));
 sky130_fd_sc_hd__mux4_2 _16873_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[398] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[430] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[462] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[494] ),
    .S0(net420),
    .S1(net412),
    .X(_09622_));
 sky130_fd_sc_hd__mux4_1 _16874_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[270] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[302] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[334] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[366] ),
    .S0(net420),
    .S1(net1072),
    .X(_09623_));
 sky130_fd_sc_hd__mux2_2 _16875_ (.A0(_09622_),
    .A1(_09623_),
    .S(_08529_),
    .X(_09624_));
 sky130_fd_sc_hd__mux2_1 _16876_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[206] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[238] ),
    .S(net437),
    .X(_09625_));
 sky130_fd_sc_hd__mux2_1 _16877_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[142] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[174] ),
    .S(net437),
    .X(_09626_));
 sky130_fd_sc_hd__o22ai_2 _16878_ (.A1(_08815_),
    .A2(_09625_),
    .B1(_09626_),
    .B2(_08811_),
    .Y(_09627_));
 sky130_fd_sc_hd__mux2_1 _16879_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[78] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[110] ),
    .S(net1084),
    .X(_09628_));
 sky130_fd_sc_hd__a221oi_4 _16880_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[46] ),
    .A2(net539),
    .B1(_09628_),
    .B2(net413),
    .C1(net400),
    .Y(_09629_));
 sky130_fd_sc_hd__nor3_1 _16881_ (.A(net1282),
    .B(_09627_),
    .C(_09629_),
    .Y(_09630_));
 sky130_fd_sc_hd__a211oi_1 _16882_ (.A1(net1282),
    .A2(_09624_),
    .B1(_09630_),
    .C1(net383),
    .Y(_09631_));
 sky130_fd_sc_hd__a31o_4 _16883_ (.A1(net383),
    .A2(_09614_),
    .A3(_09621_),
    .B1(_09631_),
    .X(_09632_));
 sky130_fd_sc_hd__o22ai_1 _16884_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[46] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[14] ),
    .B2(_08503_),
    .Y(_09633_));
 sky130_fd_sc_hd__nor2_1 _16885_ (.A(_08504_),
    .B(_09606_),
    .Y(_09634_));
 sky130_fd_sc_hd__a2111oi_2 _16886_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(_09632_),
    .B1(_09633_),
    .C1(_09634_),
    .D1(_08295_),
    .Y(_09635_));
 sky130_fd_sc_hd__a21oi_4 _16887_ (.A1(net1134),
    .A2(_09609_),
    .B1(_09635_),
    .Y(_09636_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_890 ();
 sky130_fd_sc_hd__nand2_1 _16889_ (.A(\cs_registers_i.pc_id_i[14] ),
    .B(net310),
    .Y(_09638_));
 sky130_fd_sc_hd__o21ai_0 _16890_ (.A1(net310),
    .A2(_09632_),
    .B1(_09638_),
    .Y(_09639_));
 sky130_fd_sc_hd__a22o_4 _16891_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[14] ),
    .A2(_08368_),
    .B1(_08372_),
    .B2(_09639_),
    .X(_09640_));
 sky130_fd_sc_hd__nand2_1 _16892_ (.A(net1134),
    .B(_09640_),
    .Y(_09641_));
 sky130_fd_sc_hd__nand3_1 _16893_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[46] ),
    .B(_08272_),
    .C(_08377_),
    .Y(_09642_));
 sky130_fd_sc_hd__nand2_2 _16894_ (.A(_09641_),
    .B(_09642_),
    .Y(_09643_));
 sky130_fd_sc_hd__xor2_4 _16895_ (.A(_09636_),
    .B(_09643_),
    .X(_09644_));
 sky130_fd_sc_hd__nor2_4 _16896_ (.A(_09567_),
    .B(_09492_),
    .Y(_09645_));
 sky130_fd_sc_hd__nand2_2 _16897_ (.A(_09644_),
    .B(_09645_),
    .Y(_09646_));
 sky130_fd_sc_hd__nor2_1 _16898_ (.A(_09636_),
    .B(_09643_),
    .Y(_09647_));
 sky130_fd_sc_hd__a22oi_1 _16899_ (.A1(_09452_),
    .A2(_09490_),
    .B1(_09636_),
    .B2(_09643_),
    .Y(_09648_));
 sky130_fd_sc_hd__nand2_1 _16900_ (.A(_09491_),
    .B(_09644_),
    .Y(_09649_));
 sky130_fd_sc_hd__o22a_1 _16901_ (.A1(_09647_),
    .A2(_09648_),
    .B1(_09649_),
    .B2(_09574_),
    .X(_09650_));
 sky130_fd_sc_hd__o21ai_4 _16902_ (.A1(_09646_),
    .A2(_09569_),
    .B1(_09650_),
    .Y(_09651_));
 sky130_fd_sc_hd__mux4_1 _16903_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[143] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[175] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[207] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[239] ),
    .S0(net435),
    .S1(net402),
    .X(_09652_));
 sky130_fd_sc_hd__nand2_1 _16904_ (.A(net396),
    .B(_09652_),
    .Y(_09653_));
 sky130_fd_sc_hd__mux2i_1 _16905_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[79] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[111] ),
    .S(net1129),
    .Y(_09654_));
 sky130_fd_sc_hd__a21oi_1 _16906_ (.A1(net1129),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[47] ),
    .B1(net402),
    .Y(_09655_));
 sky130_fd_sc_hd__a211o_1 _16907_ (.A1(net402),
    .A2(_09654_),
    .B1(_09655_),
    .C1(net396),
    .X(_09656_));
 sky130_fd_sc_hd__mux2i_1 _16908_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[527] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[559] ),
    .S(net901),
    .Y(_09657_));
 sky130_fd_sc_hd__mux2i_1 _16909_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[655] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[687] ),
    .S(net901),
    .Y(_09658_));
 sky130_fd_sc_hd__a22oi_2 _16910_ (.A1(net585),
    .A2(_09657_),
    .B1(_09658_),
    .B2(net618),
    .Y(_09659_));
 sky130_fd_sc_hd__mux2i_1 _16911_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[463] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[495] ),
    .S(net901),
    .Y(_09660_));
 sky130_fd_sc_hd__mux2i_1 _16912_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[591] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[623] ),
    .S(net901),
    .Y(_09661_));
 sky130_fd_sc_hd__a22oi_2 _16913_ (.A1(_08593_),
    .A2(_09660_),
    .B1(_09661_),
    .B2(net536),
    .Y(_09662_));
 sky130_fd_sc_hd__mux2i_1 _16914_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[271] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[303] ),
    .S(net901),
    .Y(_09663_));
 sky130_fd_sc_hd__mux2i_1 _16915_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[719] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[751] ),
    .S(net901),
    .Y(_09664_));
 sky130_fd_sc_hd__a22oi_2 _16916_ (.A1(net556),
    .A2(_09663_),
    .B1(_09664_),
    .B2(_08602_),
    .Y(_09665_));
 sky130_fd_sc_hd__mux2i_1 _16917_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[335] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[367] ),
    .S(net901),
    .Y(_09666_));
 sky130_fd_sc_hd__mux2i_1 _16918_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[399] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[431] ),
    .S(net901),
    .Y(_09667_));
 sky130_fd_sc_hd__a22oi_2 _16919_ (.A1(net550),
    .A2(_09666_),
    .B1(_09667_),
    .B2(net568),
    .Y(_09668_));
 sky130_fd_sc_hd__nand4_4 _16920_ (.A(_09659_),
    .B(_09662_),
    .C(_09665_),
    .D(_09668_),
    .Y(_09669_));
 sky130_fd_sc_hd__mux4_1 _16921_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[911] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[943] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[975] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1007] ),
    .S0(net429),
    .S1(net1078),
    .X(_09670_));
 sky130_fd_sc_hd__nand2_1 _16922_ (.A(net395),
    .B(_09670_),
    .Y(_09671_));
 sky130_fd_sc_hd__mux4_1 _16923_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[783] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[815] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[847] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[879] ),
    .S0(net1175),
    .S1(net1078),
    .X(_09672_));
 sky130_fd_sc_hd__nand2_1 _16924_ (.A(_08529_),
    .B(_09672_),
    .Y(_09673_));
 sky130_fd_sc_hd__and3_4 _16925_ (.A(_08618_),
    .B(_09671_),
    .C(_09673_),
    .X(_09674_));
 sky130_fd_sc_hd__a311oi_4 _16926_ (.A1(_08179_),
    .A2(_09653_),
    .A3(_09656_),
    .B1(_09674_),
    .C1(_09669_),
    .Y(_09675_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_889 ();
 sky130_fd_sc_hd__mux2i_2 _16928_ (.A0(net835),
    .A1(\cs_registers_i.pc_id_i[15] ),
    .S(net310),
    .Y(_09677_));
 sky130_fd_sc_hd__nand2_1 _16929_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[15] ),
    .B(_08368_),
    .Y(_09678_));
 sky130_fd_sc_hd__o21ai_4 _16930_ (.A1(net1115),
    .A2(_09677_),
    .B1(_09678_),
    .Y(_09679_));
 sky130_fd_sc_hd__inv_1 _16931_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[47] ),
    .Y(_09680_));
 sky130_fd_sc_hd__nor3_1 _16932_ (.A(_09680_),
    .B(net1134),
    .C(_08503_),
    .Y(_09681_));
 sky130_fd_sc_hd__a21oi_2 _16933_ (.A1(net1134),
    .A2(_09679_),
    .B1(_09681_),
    .Y(_09682_));
 sky130_fd_sc_hd__mux2_1 _16934_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[47] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[111] ),
    .S(net1077),
    .X(_09683_));
 sky130_fd_sc_hd__a221oi_4 _16935_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[79] ),
    .A2(net324),
    .B1(_09683_),
    .B2(net1133),
    .C1(net341),
    .Y(_09684_));
 sky130_fd_sc_hd__mux4_1 _16936_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[143] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[175] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[207] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[239] ),
    .S0(net374),
    .S1(net1077),
    .X(_09685_));
 sky130_fd_sc_hd__o21ai_4 _16937_ (.A1(_08481_),
    .A2(_09685_),
    .B1(_08731_),
    .Y(_09686_));
 sky130_fd_sc_hd__mux2i_2 _16938_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[399] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[463] ),
    .S(net350),
    .Y(_09687_));
 sky130_fd_sc_hd__mux2i_1 _16939_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[911] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[975] ),
    .S(net358),
    .Y(_09688_));
 sky130_fd_sc_hd__o22ai_1 _16940_ (.A1(net892),
    .A2(_09687_),
    .B1(_09688_),
    .B2(net601),
    .Y(_09689_));
 sky130_fd_sc_hd__mux2i_1 _16941_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[271] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[335] ),
    .S(net351),
    .Y(_09690_));
 sky130_fd_sc_hd__mux2i_1 _16942_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[783] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[847] ),
    .S(net358),
    .Y(_09691_));
 sky130_fd_sc_hd__o22ai_1 _16943_ (.A1(net772),
    .A2(_09690_),
    .B1(_09691_),
    .B2(net510),
    .Y(_09692_));
 sky130_fd_sc_hd__mux2i_1 _16944_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[815] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[879] ),
    .S(net358),
    .Y(_09693_));
 sky130_fd_sc_hd__mux2i_2 _16945_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[431] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[495] ),
    .S(net350),
    .Y(_09694_));
 sky130_fd_sc_hd__o22ai_1 _16946_ (.A1(net522),
    .A2(_09693_),
    .B1(_09694_),
    .B2(net870),
    .Y(_09695_));
 sky130_fd_sc_hd__mux2i_1 _16947_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[943] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1007] ),
    .S(net358),
    .Y(_09696_));
 sky130_fd_sc_hd__mux2i_1 _16948_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[303] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[367] ),
    .S(net358),
    .Y(_09697_));
 sky130_fd_sc_hd__o22ai_1 _16949_ (.A1(net632),
    .A2(_09696_),
    .B1(_09697_),
    .B2(net759),
    .Y(_09698_));
 sky130_fd_sc_hd__nor4_4 _16950_ (.A(_09689_),
    .B(_09698_),
    .C(_09695_),
    .D(_09692_),
    .Y(_09699_));
 sky130_fd_sc_hd__mux2i_1 _16951_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[559] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[623] ),
    .S(net350),
    .Y(_09700_));
 sky130_fd_sc_hd__mux2i_1 _16952_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[655] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[719] ),
    .S(net350),
    .Y(_09701_));
 sky130_fd_sc_hd__a22oi_1 _16953_ (.A1(net1201),
    .A2(_09700_),
    .B1(_09701_),
    .B2(net1013),
    .Y(_09702_));
 sky130_fd_sc_hd__mux2i_1 _16954_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[527] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[591] ),
    .S(net350),
    .Y(_09703_));
 sky130_fd_sc_hd__mux2i_1 _16955_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[687] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[751] ),
    .S(net350),
    .Y(_09704_));
 sky130_fd_sc_hd__a22oi_1 _16956_ (.A1(net650),
    .A2(_09703_),
    .B1(_09704_),
    .B2(net1153),
    .Y(_09705_));
 sky130_fd_sc_hd__nand3_2 _16957_ (.A(net698),
    .B(_09702_),
    .C(_09705_),
    .Y(_09706_));
 sky130_fd_sc_hd__o211ai_4 _16958_ (.A1(_09684_),
    .A2(_09686_),
    .B1(_09699_),
    .C1(_09706_),
    .Y(_09707_));
 sky130_fd_sc_hd__nor2_1 _16959_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[15] ),
    .B(_08503_),
    .Y(_09708_));
 sky130_fd_sc_hd__a21oi_1 _16960_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(_09680_),
    .B1(_09708_),
    .Y(_09709_));
 sky130_fd_sc_hd__o221ai_1 _16961_ (.A1(_08500_),
    .A2(net836),
    .B1(_09707_),
    .B2(_08504_),
    .C1(_09709_),
    .Y(_09710_));
 sky130_fd_sc_hd__a21oi_1 _16962_ (.A1(net1129),
    .A2(_09494_),
    .B1(_09496_),
    .Y(_09711_));
 sky130_fd_sc_hd__nand2_1 _16963_ (.A(_08495_),
    .B(_09707_),
    .Y(_09712_));
 sky130_fd_sc_hd__o21ai_2 _16964_ (.A1(_08495_),
    .A2(_09711_),
    .B1(_09712_),
    .Y(_09713_));
 sky130_fd_sc_hd__xor2_1 _16965_ (.A(net296),
    .B(_09713_),
    .X(_09714_));
 sky130_fd_sc_hd__nor2_1 _16966_ (.A(net312),
    .B(_09714_),
    .Y(_09715_));
 sky130_fd_sc_hd__a21oi_2 _16967_ (.A1(_08272_),
    .A2(_09710_),
    .B1(_09715_),
    .Y(_09716_));
 sky130_fd_sc_hd__xnor2_2 _16968_ (.A(_09682_),
    .B(_09716_),
    .Y(_09717_));
 sky130_fd_sc_hd__xnor2_4 _16969_ (.A(net769),
    .B(_09717_),
    .Y(net156));
 sky130_fd_sc_hd__o21ai_1 _16970_ (.A1(_09353_),
    .A2(_09359_),
    .B1(_09645_),
    .Y(_09718_));
 sky130_fd_sc_hd__nor2_1 _16971_ (.A(_09573_),
    .B(_09571_),
    .Y(_09719_));
 sky130_fd_sc_hd__nor2_1 _16972_ (.A(_09490_),
    .B(_09719_),
    .Y(_09720_));
 sky130_fd_sc_hd__a21oi_1 _16973_ (.A1(_09490_),
    .A2(_09719_),
    .B1(_09452_),
    .Y(_09721_));
 sky130_fd_sc_hd__o22ai_4 _16974_ (.A1(_09718_),
    .A2(_09426_),
    .B1(_09720_),
    .B2(_09721_),
    .Y(_09722_));
 sky130_fd_sc_hd__xor2_4 _16975_ (.A(_09644_),
    .B(_09722_),
    .X(net155));
 sky130_fd_sc_hd__mux4_2 _16976_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[273] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[305] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[337] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[369] ),
    .S0(net429),
    .S1(net406),
    .X(_09723_));
 sky130_fd_sc_hd__nor2_1 _16977_ (.A(_09001_),
    .B(_09723_),
    .Y(_09724_));
 sky130_fd_sc_hd__nor2b_1 _16978_ (.A(net912),
    .B_N(\gen_regfile_ff.register_file_i.rf_reg[465] ),
    .Y(_09725_));
 sky130_fd_sc_hd__a211oi_1 _16979_ (.A1(net912),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[497] ),
    .B1(_09004_),
    .C1(_09725_),
    .Y(_09726_));
 sky130_fd_sc_hd__nor2b_1 _16980_ (.A(net912),
    .B_N(\gen_regfile_ff.register_file_i.rf_reg[401] ),
    .Y(_09727_));
 sky130_fd_sc_hd__a2111oi_0 _16981_ (.A1(net912),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[433] ),
    .B1(_09007_),
    .C1(_09727_),
    .D1(net406),
    .Y(_09728_));
 sky130_fd_sc_hd__or4_4 _16982_ (.A(net384),
    .B(_09724_),
    .C(_09726_),
    .D(_09728_),
    .X(_09729_));
 sky130_fd_sc_hd__mux2i_2 _16983_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[209] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[241] ),
    .S(net435),
    .Y(_09730_));
 sky130_fd_sc_hd__mux2i_2 _16984_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[145] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[177] ),
    .S(net435),
    .Y(_09731_));
 sky130_fd_sc_hd__a22oi_2 _16985_ (.A1(_08803_),
    .A2(_09730_),
    .B1(_09731_),
    .B2(net323),
    .Y(_09732_));
 sky130_fd_sc_hd__mux2_1 _16986_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[81] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[113] ),
    .S(net435),
    .X(_09733_));
 sky130_fd_sc_hd__a221o_1 _16987_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[49] ),
    .A2(net541),
    .B1(_09733_),
    .B2(net401),
    .C1(net396),
    .X(_09734_));
 sky130_fd_sc_hd__a21oi_4 _16988_ (.A1(_09732_),
    .A2(_09734_),
    .B1(net1282),
    .Y(_09735_));
 sky130_fd_sc_hd__mux2i_1 _16989_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[785] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[817] ),
    .S(net1175),
    .Y(_09736_));
 sky130_fd_sc_hd__mux2i_1 _16990_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[913] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[945] ),
    .S(net1175),
    .Y(_09737_));
 sky130_fd_sc_hd__a22oi_2 _16991_ (.A1(net1196),
    .A2(_09736_),
    .B1(_09737_),
    .B2(net626),
    .Y(_09738_));
 sky130_fd_sc_hd__mux2i_1 _16992_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[849] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[881] ),
    .S(net429),
    .Y(_09739_));
 sky130_fd_sc_hd__mux2i_1 _16993_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[977] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1009] ),
    .S(net1175),
    .Y(_09740_));
 sky130_fd_sc_hd__a22oi_2 _16994_ (.A1(net616),
    .A2(_09739_),
    .B1(_09740_),
    .B2(_08803_),
    .Y(_09741_));
 sky130_fd_sc_hd__nand3_4 _16995_ (.A(_08618_),
    .B(_09738_),
    .C(_09741_),
    .Y(_09742_));
 sky130_fd_sc_hd__mux2i_1 _16996_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[657] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[689] ),
    .S(net1556),
    .Y(_09743_));
 sky130_fd_sc_hd__nand2_1 _16997_ (.A(net626),
    .B(_09743_),
    .Y(_09744_));
 sky130_fd_sc_hd__mux2i_1 _16998_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[593] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[625] ),
    .S(net1556),
    .Y(_09745_));
 sky130_fd_sc_hd__mux2i_1 _16999_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[529] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[561] ),
    .S(net1556),
    .Y(_09746_));
 sky130_fd_sc_hd__a22oi_2 _17000_ (.A1(net616),
    .A2(_09745_),
    .B1(_09746_),
    .B2(net1196),
    .Y(_09747_));
 sky130_fd_sc_hd__mux2i_1 _17001_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[721] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[753] ),
    .S(net1556),
    .Y(_09748_));
 sky130_fd_sc_hd__a21oi_1 _17002_ (.A1(_08803_),
    .A2(_09748_),
    .B1(_09032_),
    .Y(_09749_));
 sky130_fd_sc_hd__nand3_4 _17003_ (.A(_09744_),
    .B(_09747_),
    .C(_09749_),
    .Y(_09750_));
 sky130_fd_sc_hd__o211ai_4 _17004_ (.A1(_09735_),
    .A2(_09729_),
    .B1(_09742_),
    .C1(_09750_),
    .Y(_09751_));
 sky130_fd_sc_hd__mux2i_1 _17005_ (.A0(net776),
    .A1(\cs_registers_i.pc_id_i[17] ),
    .S(net310),
    .Y(_09752_));
 sky130_fd_sc_hd__nor2_1 _17006_ (.A(net1117),
    .B(_09752_),
    .Y(_09753_));
 sky130_fd_sc_hd__a21oi_4 _17007_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[17] ),
    .A2(_08368_),
    .B1(_09753_),
    .Y(_09754_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_888 ();
 sky130_fd_sc_hd__a21oi_1 _17009_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[49] ),
    .A2(_08377_),
    .B1(net1134),
    .Y(_09756_));
 sky130_fd_sc_hd__a21oi_2 _17010_ (.A1(_09754_),
    .A2(net1134),
    .B1(_09756_),
    .Y(_09757_));
 sky130_fd_sc_hd__inv_2 _17011_ (.A(_09757_),
    .Y(_09758_));
 sky130_fd_sc_hd__mux2_1 _17012_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[49] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[113] ),
    .S(net365),
    .X(_09759_));
 sky130_fd_sc_hd__a221oi_1 _17013_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[81] ),
    .A2(net324),
    .B1(_09759_),
    .B2(net374),
    .C1(net341),
    .Y(_09760_));
 sky130_fd_sc_hd__mux4_1 _17014_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[145] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[177] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[209] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[241] ),
    .S0(net374),
    .S1(net365),
    .X(_09761_));
 sky130_fd_sc_hd__o21ai_0 _17015_ (.A1(_08481_),
    .A2(_09761_),
    .B1(_08731_),
    .Y(_09762_));
 sky130_fd_sc_hd__nor2_2 _17016_ (.A(_09760_),
    .B(_09762_),
    .Y(_09763_));
 sky130_fd_sc_hd__mux2i_1 _17017_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[913] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[977] ),
    .S(net358),
    .Y(_09764_));
 sky130_fd_sc_hd__mux2i_1 _17018_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[945] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1009] ),
    .S(net358),
    .Y(_09765_));
 sky130_fd_sc_hd__o22ai_2 _17019_ (.A1(net601),
    .A2(_09764_),
    .B1(_09765_),
    .B2(net628),
    .Y(_09766_));
 sky130_fd_sc_hd__mux2i_1 _17020_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[433] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[497] ),
    .S(net358),
    .Y(_09767_));
 sky130_fd_sc_hd__mux2i_1 _17021_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[401] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[465] ),
    .S(net358),
    .Y(_09768_));
 sky130_fd_sc_hd__o22ai_2 _17022_ (.A1(net870),
    .A2(_09767_),
    .B1(_09768_),
    .B2(net892),
    .Y(_09769_));
 sky130_fd_sc_hd__mux2i_1 _17023_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[305] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[369] ),
    .S(net358),
    .Y(_09770_));
 sky130_fd_sc_hd__mux2i_1 _17024_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[273] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[337] ),
    .S(net358),
    .Y(_09771_));
 sky130_fd_sc_hd__o22ai_2 _17025_ (.A1(net759),
    .A2(_09770_),
    .B1(_09771_),
    .B2(net772),
    .Y(_09772_));
 sky130_fd_sc_hd__mux2i_2 _17026_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[817] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[881] ),
    .S(net358),
    .Y(_09773_));
 sky130_fd_sc_hd__mux2i_2 _17027_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[785] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[849] ),
    .S(net358),
    .Y(_09774_));
 sky130_fd_sc_hd__o22ai_4 _17028_ (.A1(net521),
    .A2(_09773_),
    .B1(_09774_),
    .B2(net508),
    .Y(_09775_));
 sky130_fd_sc_hd__nor4_4 _17029_ (.A(_09775_),
    .B(_09769_),
    .C(_09772_),
    .D(_09766_),
    .Y(_09776_));
 sky130_fd_sc_hd__mux2i_1 _17030_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[529] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[593] ),
    .S(net1093),
    .Y(_09777_));
 sky130_fd_sc_hd__mux2i_1 _17031_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[657] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[721] ),
    .S(net1093),
    .Y(_09778_));
 sky130_fd_sc_hd__a22oi_1 _17032_ (.A1(net325),
    .A2(_09777_),
    .B1(_09778_),
    .B2(net1119),
    .Y(_09779_));
 sky130_fd_sc_hd__mux2i_1 _17033_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[561] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[625] ),
    .S(net1093),
    .Y(_09780_));
 sky130_fd_sc_hd__mux2i_1 _17034_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[689] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[753] ),
    .S(net1093),
    .Y(_09781_));
 sky130_fd_sc_hd__a22oi_1 _17035_ (.A1(net328),
    .A2(_09780_),
    .B1(_09781_),
    .B2(net1153),
    .Y(_09782_));
 sky130_fd_sc_hd__nand3_2 _17036_ (.A(_08462_),
    .B(_09779_),
    .C(_09782_),
    .Y(_09783_));
 sky130_fd_sc_hd__nand3b_4 _17037_ (.A_N(_09763_),
    .B(_09783_),
    .C(net1304),
    .Y(_09784_));
 sky130_fd_sc_hd__o22a_1 _17038_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[49] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[17] ),
    .B2(_08503_),
    .X(_09785_));
 sky130_fd_sc_hd__o221ai_2 _17039_ (.A1(_08500_),
    .A2(net776),
    .B1(_09784_),
    .B2(_08504_),
    .C1(_09785_),
    .Y(_09786_));
 sky130_fd_sc_hd__o21ai_1 _17040_ (.A1(_09455_),
    .A2(_09458_),
    .B1(net396),
    .Y(_09787_));
 sky130_fd_sc_hd__nor2_2 _17041_ (.A(_08436_),
    .B(_09784_),
    .Y(_09788_));
 sky130_fd_sc_hd__a31oi_4 _17042_ (.A1(_08436_),
    .A2(_09457_),
    .A3(_09787_),
    .B1(_09788_),
    .Y(_09789_));
 sky130_fd_sc_hd__xor2_1 _17043_ (.A(net296),
    .B(_09789_),
    .X(_09790_));
 sky130_fd_sc_hd__nor2_1 _17044_ (.A(net312),
    .B(_09790_),
    .Y(_09791_));
 sky130_fd_sc_hd__a21oi_2 _17045_ (.A1(_08272_),
    .A2(_09786_),
    .B1(_09791_),
    .Y(_09792_));
 sky130_fd_sc_hd__xnor2_4 _17046_ (.A(_09792_),
    .B(_09758_),
    .Y(_09793_));
 sky130_fd_sc_hd__mux2i_1 _17047_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[208] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[240] ),
    .S(net434),
    .Y(_09794_));
 sky130_fd_sc_hd__mux2i_1 _17048_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[80] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[112] ),
    .S(net434),
    .Y(_09795_));
 sky130_fd_sc_hd__o22ai_1 _17049_ (.A1(_08815_),
    .A2(_09794_),
    .B1(_09795_),
    .B2(_08819_),
    .Y(_09796_));
 sky130_fd_sc_hd__mux2_1 _17050_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[144] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[176] ),
    .S(net434),
    .X(_09797_));
 sky130_fd_sc_hd__a32o_1 _17051_ (.A1(net434),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[48] ),
    .A3(net649),
    .B1(net1149),
    .B2(_09797_),
    .X(_09798_));
 sky130_fd_sc_hd__or3_2 _17052_ (.A(_08821_),
    .B(_09796_),
    .C(_09798_),
    .X(_09799_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_887 ();
 sky130_fd_sc_hd__mux2i_1 _17054_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[720] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[752] ),
    .S(net1556),
    .Y(_09801_));
 sky130_fd_sc_hd__mux2i_1 _17055_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[592] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[624] ),
    .S(net1556),
    .Y(_09802_));
 sky130_fd_sc_hd__a22oi_1 _17056_ (.A1(_08602_),
    .A2(_09801_),
    .B1(_09802_),
    .B2(net537),
    .Y(_09803_));
 sky130_fd_sc_hd__mux2i_1 _17057_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[656] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[688] ),
    .S(net428),
    .Y(_09804_));
 sky130_fd_sc_hd__mux2i_1 _17058_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[528] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[560] ),
    .S(net1556),
    .Y(_09805_));
 sky130_fd_sc_hd__a22oi_1 _17059_ (.A1(net621),
    .A2(_09804_),
    .B1(_09805_),
    .B2(net586),
    .Y(_09806_));
 sky130_fd_sc_hd__mux2i_1 _17060_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[464] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[496] ),
    .S(net912),
    .Y(_09807_));
 sky130_fd_sc_hd__mux2i_1 _17061_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[400] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[432] ),
    .S(net912),
    .Y(_09808_));
 sky130_fd_sc_hd__a22oi_1 _17062_ (.A1(_08593_),
    .A2(_09807_),
    .B1(_09808_),
    .B2(net1118),
    .Y(_09809_));
 sky130_fd_sc_hd__mux2i_1 _17063_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[272] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[304] ),
    .S(net1175),
    .Y(_09810_));
 sky130_fd_sc_hd__mux2i_1 _17064_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[336] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[368] ),
    .S(net1175),
    .Y(_09811_));
 sky130_fd_sc_hd__a22oi_1 _17065_ (.A1(_08597_),
    .A2(_09810_),
    .B1(_09811_),
    .B2(net876),
    .Y(_09812_));
 sky130_fd_sc_hd__and4_4 _17066_ (.A(_09803_),
    .B(_09806_),
    .C(_09809_),
    .D(_09812_),
    .X(_09813_));
 sky130_fd_sc_hd__mux2i_1 _17067_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[912] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[944] ),
    .S(net1074),
    .Y(_09814_));
 sky130_fd_sc_hd__mux2i_1 _17068_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[784] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[816] ),
    .S(net433),
    .Y(_09815_));
 sky130_fd_sc_hd__a22oi_1 _17069_ (.A1(net323),
    .A2(_09814_),
    .B1(_09815_),
    .B2(net1199),
    .Y(_09816_));
 sky130_fd_sc_hd__mux2i_1 _17070_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[976] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1008] ),
    .S(net432),
    .Y(_09817_));
 sky130_fd_sc_hd__mux2i_1 _17071_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[848] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[880] ),
    .S(net433),
    .Y(_09818_));
 sky130_fd_sc_hd__a22oi_1 _17072_ (.A1(_08803_),
    .A2(_09817_),
    .B1(_09818_),
    .B2(net614),
    .Y(_09819_));
 sky130_fd_sc_hd__a21o_2 _17073_ (.A1(_09816_),
    .A2(_09819_),
    .B1(_08809_),
    .X(_09820_));
 sky130_fd_sc_hd__nand3_4 _17074_ (.A(_09799_),
    .B(_09813_),
    .C(_09820_),
    .Y(_09821_));
 sky130_fd_sc_hd__nor2_1 _17075_ (.A(net310),
    .B(_09821_),
    .Y(_09822_));
 sky130_fd_sc_hd__a21oi_1 _17076_ (.A1(\cs_registers_i.pc_id_i[16] ),
    .A2(net310),
    .B1(_09822_),
    .Y(_09823_));
 sky130_fd_sc_hd__nand2_1 _17077_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[16] ),
    .B(_08368_),
    .Y(_09824_));
 sky130_fd_sc_hd__o21ai_4 _17078_ (.A1(net933),
    .A2(_09823_),
    .B1(_09824_),
    .Y(_09825_));
 sky130_fd_sc_hd__nand2_1 _17079_ (.A(net739),
    .B(_09825_),
    .Y(_09826_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_886 ();
 sky130_fd_sc_hd__nand3_1 _17081_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[48] ),
    .B(_08272_),
    .C(_08377_),
    .Y(_09828_));
 sky130_fd_sc_hd__nand2_2 _17082_ (.A(_09826_),
    .B(_09828_),
    .Y(_09829_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_885 ();
 sky130_fd_sc_hd__mux4_4 _17084_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[272] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[304] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[336] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[368] ),
    .S0(net373),
    .S1(net358),
    .X(_09831_));
 sky130_fd_sc_hd__mux2_1 _17085_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[48] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[112] ),
    .S(net1141),
    .X(_09832_));
 sky130_fd_sc_hd__a221o_1 _17086_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[80] ),
    .A2(net324),
    .B1(_09832_),
    .B2(net1133),
    .C1(net336),
    .X(_09833_));
 sky130_fd_sc_hd__o211ai_4 _17087_ (.A1(_08162_),
    .A2(_09831_),
    .B1(_09833_),
    .C1(_08491_),
    .Y(_09834_));
 sky130_fd_sc_hd__mux4_1 _17088_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[144] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[208] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[400] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[464] ),
    .S0(net363),
    .S1(net336),
    .X(_09835_));
 sky130_fd_sc_hd__nor2b_1 _17089_ (.A(net336),
    .B_N(net1133),
    .Y(_09836_));
 sky130_fd_sc_hd__mux2i_1 _17090_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[176] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[240] ),
    .S(net1141),
    .Y(_09837_));
 sky130_fd_sc_hd__a2bb2oi_1 _17091_ (.A1_N(net1133),
    .A2_N(_09835_),
    .B1(_09836_),
    .B2(_09837_),
    .Y(_09838_));
 sky130_fd_sc_hd__mux2i_1 _17092_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[432] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[496] ),
    .S(net1093),
    .Y(_09839_));
 sky130_fd_sc_hd__nand3_2 _17093_ (.A(net336),
    .B(net373),
    .C(_09839_),
    .Y(_09840_));
 sky130_fd_sc_hd__nand4_2 _17094_ (.A(_08161_),
    .B(net341),
    .C(_09838_),
    .D(_09840_),
    .Y(_09841_));
 sky130_fd_sc_hd__mux2i_1 _17095_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[560] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[624] ),
    .S(net357),
    .Y(_09842_));
 sky130_fd_sc_hd__mux2i_1 _17096_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[656] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[720] ),
    .S(net1093),
    .Y(_09843_));
 sky130_fd_sc_hd__a22oi_2 _17097_ (.A1(_09842_),
    .A2(net329),
    .B1(_09843_),
    .B2(net1119),
    .Y(_09844_));
 sky130_fd_sc_hd__mux2i_1 _17098_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[528] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[592] ),
    .S(net357),
    .Y(_09845_));
 sky130_fd_sc_hd__mux2i_1 _17099_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[688] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[752] ),
    .S(net1093),
    .Y(_09846_));
 sky130_fd_sc_hd__a22oi_2 _17100_ (.A1(net325),
    .A2(_09845_),
    .B1(_09846_),
    .B2(net1153),
    .Y(_09847_));
 sky130_fd_sc_hd__nand3_4 _17101_ (.A(_08462_),
    .B(_09844_),
    .C(_09847_),
    .Y(_09848_));
 sky130_fd_sc_hd__mux2i_1 _17102_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[816] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[880] ),
    .S(net361),
    .Y(_09849_));
 sky130_fd_sc_hd__mux2i_1 _17103_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[944] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1008] ),
    .S(net361),
    .Y(_09850_));
 sky130_fd_sc_hd__o22ai_1 _17104_ (.A1(net930),
    .A2(_09849_),
    .B1(_09850_),
    .B2(net1210),
    .Y(_09851_));
 sky130_fd_sc_hd__mux2i_1 _17105_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[784] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[848] ),
    .S(net361),
    .Y(_09852_));
 sky130_fd_sc_hd__mux2i_1 _17106_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[912] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[976] ),
    .S(net361),
    .Y(_09853_));
 sky130_fd_sc_hd__o22ai_1 _17107_ (.A1(net506),
    .A2(_09852_),
    .B1(_09853_),
    .B2(net935),
    .Y(_09854_));
 sky130_fd_sc_hd__nor2_2 _17108_ (.A(_09851_),
    .B(_09854_),
    .Y(_09855_));
 sky130_fd_sc_hd__and4_4 _17109_ (.A(_09834_),
    .B(_09841_),
    .C(_09848_),
    .D(_09855_),
    .X(_09856_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_884 ();
 sky130_fd_sc_hd__a211oi_1 _17111_ (.A1(net402),
    .A2(_09494_),
    .B1(_09496_),
    .C1(_08495_),
    .Y(_09858_));
 sky130_fd_sc_hd__a21oi_2 _17112_ (.A1(_08495_),
    .A2(_09856_),
    .B1(_09858_),
    .Y(_09859_));
 sky130_fd_sc_hd__xnor2_1 _17113_ (.A(net296),
    .B(_09859_),
    .Y(_09860_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_883 ();
 sky130_fd_sc_hd__o22ai_1 _17115_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[48] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[16] ),
    .B2(_08503_),
    .Y(_09862_));
 sky130_fd_sc_hd__a221oi_1 _17116_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(_09821_),
    .B1(_09856_),
    .B2(_08696_),
    .C1(_09862_),
    .Y(_09863_));
 sky130_fd_sc_hd__nand2_1 _17117_ (.A(net314),
    .B(_09863_),
    .Y(_09864_));
 sky130_fd_sc_hd__o21ai_2 _17118_ (.A1(net314),
    .A2(_09860_),
    .B1(_09864_),
    .Y(_09865_));
 sky130_fd_sc_hd__xor2_4 _17119_ (.A(_09829_),
    .B(_09865_),
    .X(_09866_));
 sky130_fd_sc_hd__nor2_1 _17120_ (.A(_09717_),
    .B(_09866_),
    .Y(_09867_));
 sky130_fd_sc_hd__inv_1 _17121_ (.A(_09865_),
    .Y(_09868_));
 sky130_fd_sc_hd__nor2_1 _17122_ (.A(_09682_),
    .B(_09716_),
    .Y(_09869_));
 sky130_fd_sc_hd__maj3_1 _17123_ (.A(_09829_),
    .B(_09868_),
    .C(_09869_),
    .X(_09870_));
 sky130_fd_sc_hd__a21oi_4 _17124_ (.A1(_09651_),
    .A2(_09867_),
    .B1(_09870_),
    .Y(_09871_));
 sky130_fd_sc_hd__xor2_4 _17125_ (.A(_09793_),
    .B(_09871_),
    .X(net158));
 sky130_fd_sc_hd__nand2_1 _17126_ (.A(_09682_),
    .B(_09716_),
    .Y(_09872_));
 sky130_fd_sc_hd__a21oi_2 _17127_ (.A1(_09651_),
    .A2(_09872_),
    .B1(_09869_),
    .Y(_09873_));
 sky130_fd_sc_hd__xor2_4 _17128_ (.A(_09866_),
    .B(_09873_),
    .X(net157));
 sky130_fd_sc_hd__mux4_1 _17129_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[914] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[946] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[978] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1010] ),
    .S0(net423),
    .S1(net1204),
    .X(_09874_));
 sky130_fd_sc_hd__nand2_1 _17130_ (.A(net393),
    .B(_09874_),
    .Y(_09875_));
 sky130_fd_sc_hd__mux4_1 _17131_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[786] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[818] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[850] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[882] ),
    .S0(net1016),
    .S1(net408),
    .X(_09876_));
 sky130_fd_sc_hd__nand2_1 _17132_ (.A(_08529_),
    .B(_09876_),
    .Y(_09877_));
 sky130_fd_sc_hd__and3_2 _17133_ (.A(_08618_),
    .B(_09875_),
    .C(_09877_),
    .X(_09878_));
 sky130_fd_sc_hd__mux2i_1 _17134_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[210] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[242] ),
    .S(net437),
    .Y(_09879_));
 sky130_fd_sc_hd__mux2i_1 _17135_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[146] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[178] ),
    .S(net437),
    .Y(_09880_));
 sky130_fd_sc_hd__a22oi_1 _17136_ (.A1(_08803_),
    .A2(_09879_),
    .B1(_09880_),
    .B2(net323),
    .Y(_09881_));
 sky130_fd_sc_hd__mux2_1 _17137_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[82] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[114] ),
    .S(net437),
    .X(_09882_));
 sky130_fd_sc_hd__a221o_1 _17138_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[50] ),
    .A2(net539),
    .B1(_09882_),
    .B2(net403),
    .C1(net397),
    .X(_09883_));
 sky130_fd_sc_hd__a21oi_2 _17139_ (.A1(_09881_),
    .A2(_09883_),
    .B1(_08821_),
    .Y(_09884_));
 sky130_fd_sc_hd__mux2_1 _17140_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[530] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[562] ),
    .S(net424),
    .X(_09885_));
 sky130_fd_sc_hd__mux2_1 _17141_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[594] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[626] ),
    .S(net424),
    .X(_09886_));
 sky130_fd_sc_hd__mux2_1 _17142_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[658] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[690] ),
    .S(net424),
    .X(_09887_));
 sky130_fd_sc_hd__a222oi_1 _17143_ (.A1(_08187_),
    .A2(_09885_),
    .B1(_09886_),
    .B2(_08807_),
    .C1(_09887_),
    .C2(net622),
    .Y(_09888_));
 sky130_fd_sc_hd__mux2_1 _17144_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[722] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[754] ),
    .S(net424),
    .X(_09889_));
 sky130_fd_sc_hd__a21oi_1 _17145_ (.A1(_08803_),
    .A2(_09889_),
    .B1(_09032_),
    .Y(_09890_));
 sky130_fd_sc_hd__mux4_1 _17146_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[402] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[434] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[466] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[498] ),
    .S0(net425),
    .S1(net408),
    .X(_09891_));
 sky130_fd_sc_hd__mux4_1 _17147_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[274] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[306] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[338] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[370] ),
    .S0(net425),
    .S1(net1204),
    .X(_09892_));
 sky130_fd_sc_hd__mux2_2 _17148_ (.A0(_09891_),
    .A1(_09892_),
    .S(_08529_),
    .X(_09893_));
 sky130_fd_sc_hd__o2bb2ai_2 _17149_ (.A1_N(_09888_),
    .A2_N(_09890_),
    .B1(_09893_),
    .B2(_09275_),
    .Y(_09894_));
 sky130_fd_sc_hd__nor3_4 _17150_ (.A(_09894_),
    .B(_09884_),
    .C(_09878_),
    .Y(_09895_));
 sky130_fd_sc_hd__mux2i_2 _17151_ (.A0(net961),
    .A1(\cs_registers_i.pc_id_i[18] ),
    .S(net310),
    .Y(_09896_));
 sky130_fd_sc_hd__nand2_1 _17152_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[18] ),
    .B(_08368_),
    .Y(_09897_));
 sky130_fd_sc_hd__o21ai_4 _17153_ (.A1(net1117),
    .A2(_09896_),
    .B1(_09897_),
    .Y(_09898_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_882 ();
 sky130_fd_sc_hd__and3_1 _17155_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[50] ),
    .B(_08272_),
    .C(_08377_),
    .X(_09900_));
 sky130_fd_sc_hd__a21oi_2 _17156_ (.A1(_08290_),
    .A2(_09898_),
    .B1(_09900_),
    .Y(_09901_));
 sky130_fd_sc_hd__mux2i_1 _17157_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[818] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[882] ),
    .S(net354),
    .Y(_09902_));
 sky130_fd_sc_hd__nor2b_1 _17158_ (.A(net354),
    .B_N(\gen_regfile_ff.register_file_i.rf_reg[946] ),
    .Y(_09903_));
 sky130_fd_sc_hd__a211oi_1 _17159_ (.A1(net354),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[1010] ),
    .B1(_08705_),
    .C1(_09903_),
    .Y(_09904_));
 sky130_fd_sc_hd__mux2i_1 _17160_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[914] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[978] ),
    .S(net354),
    .Y(_09905_));
 sky130_fd_sc_hd__mux2i_1 _17161_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[786] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[850] ),
    .S(net354),
    .Y(_09906_));
 sky130_fd_sc_hd__a22o_1 _17162_ (.A1(net326),
    .A2(_09905_),
    .B1(_09906_),
    .B2(net325),
    .X(_09907_));
 sky130_fd_sc_hd__a2111oi_2 _17163_ (.A1(net328),
    .A2(_09902_),
    .B1(_09904_),
    .C1(_08708_),
    .D1(_09907_),
    .Y(_09908_));
 sky130_fd_sc_hd__mux2i_1 _17164_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[690] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[754] ),
    .S(net353),
    .Y(_09909_));
 sky130_fd_sc_hd__mux2i_1 _17165_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[562] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[626] ),
    .S(net353),
    .Y(_09910_));
 sky130_fd_sc_hd__a22oi_1 _17166_ (.A1(_08152_),
    .A2(_09909_),
    .B1(_09910_),
    .B2(net328),
    .Y(_09911_));
 sky130_fd_sc_hd__mux2i_1 _17167_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[530] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[594] ),
    .S(net353),
    .Y(_09912_));
 sky130_fd_sc_hd__mux2i_1 _17168_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[658] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[722] ),
    .S(net353),
    .Y(_09913_));
 sky130_fd_sc_hd__a22oi_1 _17169_ (.A1(net325),
    .A2(_09912_),
    .B1(_09913_),
    .B2(net326),
    .Y(_09914_));
 sky130_fd_sc_hd__and3_1 _17170_ (.A(_08462_),
    .B(_09911_),
    .C(_09914_),
    .X(_09915_));
 sky130_fd_sc_hd__mux2i_1 _17171_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[274] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[338] ),
    .S(net349),
    .Y(_09916_));
 sky130_fd_sc_hd__mux2i_1 _17172_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[402] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[466] ),
    .S(net349),
    .Y(_09917_));
 sky130_fd_sc_hd__a22oi_1 _17173_ (.A1(net325),
    .A2(_09916_),
    .B1(_09917_),
    .B2(net327),
    .Y(_09918_));
 sky130_fd_sc_hd__mux2i_1 _17174_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[306] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[370] ),
    .S(net352),
    .Y(_09919_));
 sky130_fd_sc_hd__mux2i_1 _17175_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[434] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[498] ),
    .S(net349),
    .Y(_09920_));
 sky130_fd_sc_hd__a22oi_1 _17176_ (.A1(net329),
    .A2(_09919_),
    .B1(_09920_),
    .B2(_08152_),
    .Y(_09921_));
 sky130_fd_sc_hd__and3_1 _17177_ (.A(net703),
    .B(_09918_),
    .C(_09921_),
    .X(_09922_));
 sky130_fd_sc_hd__mux2_1 _17178_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[82] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[210] ),
    .S(net341),
    .X(_09923_));
 sky130_fd_sc_hd__a221oi_1 _17179_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[146] ),
    .A2(_08669_),
    .B1(_09923_),
    .B2(net364),
    .C1(net380),
    .Y(_09924_));
 sky130_fd_sc_hd__mux4_1 _17180_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[50] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[114] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[178] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[242] ),
    .S0(net364),
    .S1(net341),
    .X(_09925_));
 sky130_fd_sc_hd__o21ai_2 _17181_ (.A1(_08658_),
    .A2(_09925_),
    .B1(_08731_),
    .Y(_09926_));
 sky130_fd_sc_hd__nor2_2 _17182_ (.A(_09924_),
    .B(_09926_),
    .Y(_09927_));
 sky130_fd_sc_hd__nor4_4 _17183_ (.A(_09908_),
    .B(_09927_),
    .C(_09922_),
    .D(_09915_),
    .Y(_09928_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_880 ();
 sky130_fd_sc_hd__a211oi_1 _17186_ (.A1(net1140),
    .A2(_09494_),
    .B1(_09496_),
    .C1(_08495_),
    .Y(_09931_));
 sky130_fd_sc_hd__a21oi_2 _17187_ (.A1(_08495_),
    .A2(net305),
    .B1(_09931_),
    .Y(_09932_));
 sky130_fd_sc_hd__xnor2_1 _17188_ (.A(net296),
    .B(_09932_),
    .Y(_09933_));
 sky130_fd_sc_hd__o22ai_1 _17189_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[50] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[18] ),
    .B2(_08503_),
    .Y(_09934_));
 sky130_fd_sc_hd__a21oi_1 _17190_ (.A1(_08696_),
    .A2(net305),
    .B1(_09934_),
    .Y(_09935_));
 sky130_fd_sc_hd__o211ai_1 _17191_ (.A1(_08500_),
    .A2(net960),
    .B1(_09935_),
    .C1(net314),
    .Y(_09936_));
 sky130_fd_sc_hd__o21ai_2 _17192_ (.A1(net314),
    .A2(_09933_),
    .B1(_09936_),
    .Y(_09937_));
 sky130_fd_sc_hd__xnor2_2 _17193_ (.A(_09901_),
    .B(_09937_),
    .Y(_09938_));
 sky130_fd_sc_hd__or2_1 _17194_ (.A(_09938_),
    .B(_09793_),
    .X(_09939_));
 sky130_fd_sc_hd__nand2_1 _17195_ (.A(_09901_),
    .B(_09937_),
    .Y(_09940_));
 sky130_fd_sc_hd__o22ai_1 _17196_ (.A1(_09758_),
    .A2(_09792_),
    .B1(_09901_),
    .B2(_09937_),
    .Y(_09941_));
 sky130_fd_sc_hd__nand2_1 _17197_ (.A(_09940_),
    .B(_09941_),
    .Y(_09942_));
 sky130_fd_sc_hd__o21ai_2 _17198_ (.A1(_09871_),
    .A2(_09939_),
    .B1(_09942_),
    .Y(_09943_));
 sky130_fd_sc_hd__mux2_1 _17199_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[787] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[819] ),
    .S(net424),
    .X(_09944_));
 sky130_fd_sc_hd__nand2b_1 _17200_ (.A_N(\gen_regfile_ff.register_file_i.rf_reg[883] ),
    .B(net424),
    .Y(_09945_));
 sky130_fd_sc_hd__o221ai_2 _17201_ (.A1(net424),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[851] ),
    .B1(_09944_),
    .B2(net406),
    .C1(_09945_),
    .Y(_09946_));
 sky130_fd_sc_hd__mux2_1 _17202_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[915] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[947] ),
    .S(net424),
    .X(_09947_));
 sky130_fd_sc_hd__mux2_1 _17203_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[979] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1011] ),
    .S(net424),
    .X(_09948_));
 sky130_fd_sc_hd__o211ai_2 _17204_ (.A1(net406),
    .A2(_09947_),
    .B1(_09948_),
    .C1(net395),
    .Y(_09949_));
 sky130_fd_sc_hd__a221oi_2 _17205_ (.A1(net624),
    .A2(_09947_),
    .B1(_09944_),
    .B2(net649),
    .C1(_08809_),
    .Y(_09950_));
 sky130_fd_sc_hd__o211ai_4 _17206_ (.A1(net395),
    .A2(_09946_),
    .B1(_09949_),
    .C1(_09950_),
    .Y(_09951_));
 sky130_fd_sc_hd__mux4_1 _17207_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[83] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[115] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[211] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[243] ),
    .S0(net436),
    .S1(net396),
    .X(_09952_));
 sky130_fd_sc_hd__mux2_1 _17208_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[147] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[179] ),
    .S(net436),
    .X(_09953_));
 sky130_fd_sc_hd__a32o_1 _17209_ (.A1(net436),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[51] ),
    .A3(net1198),
    .B1(net323),
    .B2(_09953_),
    .X(_09954_));
 sky130_fd_sc_hd__a211o_2 _17210_ (.A1(net401),
    .A2(_09952_),
    .B1(_09954_),
    .C1(_08821_),
    .X(_09955_));
 sky130_fd_sc_hd__mux2i_1 _17211_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[275] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[307] ),
    .S(net938),
    .Y(_09956_));
 sky130_fd_sc_hd__mux2i_1 _17212_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[531] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[563] ),
    .S(net938),
    .Y(_09957_));
 sky130_fd_sc_hd__a22oi_1 _17213_ (.A1(net557),
    .A2(_09956_),
    .B1(_09957_),
    .B2(net863),
    .Y(_09958_));
 sky130_fd_sc_hd__mux2i_1 _17214_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[339] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[371] ),
    .S(net938),
    .Y(_09959_));
 sky130_fd_sc_hd__mux2i_1 _17215_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[403] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[435] ),
    .S(net938),
    .Y(_09960_));
 sky130_fd_sc_hd__a22oi_1 _17216_ (.A1(net713),
    .A2(_09959_),
    .B1(_09960_),
    .B2(net566),
    .Y(_09961_));
 sky130_fd_sc_hd__mux2i_1 _17217_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[659] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[691] ),
    .S(net733),
    .Y(_09962_));
 sky130_fd_sc_hd__mux2i_1 _17218_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[595] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[627] ),
    .S(net938),
    .Y(_09963_));
 sky130_fd_sc_hd__a22oi_1 _17219_ (.A1(net619),
    .A2(_09962_),
    .B1(_09963_),
    .B2(net716),
    .Y(_09964_));
 sky130_fd_sc_hd__mux2i_1 _17220_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[723] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[755] ),
    .S(net733),
    .Y(_09965_));
 sky130_fd_sc_hd__mux2i_1 _17221_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[467] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[499] ),
    .S(net938),
    .Y(_09966_));
 sky130_fd_sc_hd__a22oi_1 _17222_ (.A1(_08602_),
    .A2(_09965_),
    .B1(_09966_),
    .B2(_08593_),
    .Y(_09967_));
 sky130_fd_sc_hd__and4_4 _17223_ (.A(_09958_),
    .B(_09961_),
    .C(_09964_),
    .D(_09967_),
    .X(_09968_));
 sky130_fd_sc_hd__nand3_4 _17224_ (.A(_09951_),
    .B(_09955_),
    .C(_09968_),
    .Y(_09969_));
 sky130_fd_sc_hd__mux4_1 _17225_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[563] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[627] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[691] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[755] ),
    .S0(net349),
    .S1(net340),
    .X(_09970_));
 sky130_fd_sc_hd__mux2i_1 _17226_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[659] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[723] ),
    .S(net349),
    .Y(_09971_));
 sky130_fd_sc_hd__nand2_1 _17227_ (.A(net1013),
    .B(_09971_),
    .Y(_09972_));
 sky130_fd_sc_hd__mux2i_1 _17228_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[531] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[595] ),
    .S(net349),
    .Y(_09973_));
 sky130_fd_sc_hd__a21oi_1 _17229_ (.A1(net1045),
    .A2(_09973_),
    .B1(_08679_),
    .Y(_09974_));
 sky130_fd_sc_hd__o211a_1 _17230_ (.A1(_08658_),
    .A2(_09970_),
    .B1(_09972_),
    .C1(_09974_),
    .X(_09975_));
 sky130_fd_sc_hd__mux2i_2 _17231_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[915] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[979] ),
    .S(net359),
    .Y(_09976_));
 sky130_fd_sc_hd__nor2b_1 _17232_ (.A(net359),
    .B_N(\gen_regfile_ff.register_file_i.rf_reg[947] ),
    .Y(_09977_));
 sky130_fd_sc_hd__a211oi_2 _17233_ (.A1(net359),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[1011] ),
    .B1(_08705_),
    .C1(_09977_),
    .Y(_09978_));
 sky130_fd_sc_hd__mux2i_1 _17234_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[819] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[883] ),
    .S(net359),
    .Y(_09979_));
 sky130_fd_sc_hd__mux2i_1 _17235_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[787] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[851] ),
    .S(net359),
    .Y(_09980_));
 sky130_fd_sc_hd__a22o_1 _17236_ (.A1(net328),
    .A2(_09979_),
    .B1(_09980_),
    .B2(net325),
    .X(_09981_));
 sky130_fd_sc_hd__a2111oi_4 _17237_ (.A1(net1119),
    .A2(_09976_),
    .B1(_09978_),
    .C1(_09981_),
    .D1(_08708_),
    .Y(_09982_));
 sky130_fd_sc_hd__mux2_1 _17238_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[83] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[211] ),
    .S(net340),
    .X(_09983_));
 sky130_fd_sc_hd__a221oi_2 _17239_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[147] ),
    .A2(_08669_),
    .B1(_09983_),
    .B2(net1141),
    .C1(net983),
    .Y(_09984_));
 sky130_fd_sc_hd__mux4_1 _17240_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[51] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[115] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[179] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[243] ),
    .S0(net363),
    .S1(net340),
    .X(_09985_));
 sky130_fd_sc_hd__o21ai_1 _17241_ (.A1(_08658_),
    .A2(_09985_),
    .B1(_08731_),
    .Y(_09986_));
 sky130_fd_sc_hd__nor2_4 _17242_ (.A(_09984_),
    .B(_09986_),
    .Y(_09987_));
 sky130_fd_sc_hd__mux2i_1 _17243_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[275] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[339] ),
    .S(net351),
    .Y(_09988_));
 sky130_fd_sc_hd__mux2i_1 _17244_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[403] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[467] ),
    .S(net351),
    .Y(_09989_));
 sky130_fd_sc_hd__a22oi_1 _17245_ (.A1(net325),
    .A2(_09988_),
    .B1(_09989_),
    .B2(net1474),
    .Y(_09990_));
 sky130_fd_sc_hd__mux2i_1 _17246_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[307] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[371] ),
    .S(net350),
    .Y(_09991_));
 sky130_fd_sc_hd__mux2i_1 _17247_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[435] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[499] ),
    .S(net350),
    .Y(_09992_));
 sky130_fd_sc_hd__a22oi_1 _17248_ (.A1(net329),
    .A2(_09991_),
    .B1(_09992_),
    .B2(_08152_),
    .Y(_09993_));
 sky130_fd_sc_hd__and3_1 _17249_ (.A(net702),
    .B(_09990_),
    .C(_09993_),
    .X(_09994_));
 sky130_fd_sc_hd__nor4_4 _17250_ (.A(_09975_),
    .B(_09982_),
    .C(_09987_),
    .D(_09994_),
    .Y(_09995_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_878 ();
 sky130_fd_sc_hd__o22ai_1 _17253_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[51] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[19] ),
    .B2(_08503_),
    .Y(_09998_));
 sky130_fd_sc_hd__a221oi_1 _17254_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(_09969_),
    .B1(net304),
    .B2(_08696_),
    .C1(_09998_),
    .Y(_09999_));
 sky130_fd_sc_hd__a211oi_1 _17255_ (.A1(net385),
    .A2(_09494_),
    .B1(_09496_),
    .C1(_08495_),
    .Y(_10000_));
 sky130_fd_sc_hd__a21oi_2 _17256_ (.A1(_08495_),
    .A2(net304),
    .B1(_10000_),
    .Y(_10001_));
 sky130_fd_sc_hd__xnor2_1 _17257_ (.A(net296),
    .B(_10001_),
    .Y(_10002_));
 sky130_fd_sc_hd__nand2_1 _17258_ (.A(net1134),
    .B(_10002_),
    .Y(_10003_));
 sky130_fd_sc_hd__o21ai_2 _17259_ (.A1(_08290_),
    .A2(_09999_),
    .B1(_10003_),
    .Y(_10004_));
 sky130_fd_sc_hd__nor2_1 _17260_ (.A(net310),
    .B(_09969_),
    .Y(_10005_));
 sky130_fd_sc_hd__a21oi_1 _17261_ (.A1(\cs_registers_i.pc_id_i[19] ),
    .A2(net310),
    .B1(_10005_),
    .Y(_10006_));
 sky130_fd_sc_hd__nand2_1 _17262_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[19] ),
    .B(_08368_),
    .Y(_10007_));
 sky130_fd_sc_hd__o21ai_4 _17263_ (.A1(net933),
    .A2(_10006_),
    .B1(_10007_),
    .Y(_10008_));
 sky130_fd_sc_hd__nand2_1 _17264_ (.A(net739),
    .B(_10008_),
    .Y(_10009_));
 sky130_fd_sc_hd__nand3_1 _17265_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[51] ),
    .B(_08272_),
    .C(_08377_),
    .Y(_10010_));
 sky130_fd_sc_hd__nand2_2 _17266_ (.A(_10009_),
    .B(_10010_),
    .Y(_10011_));
 sky130_fd_sc_hd__xnor2_2 _17267_ (.A(_10004_),
    .B(_10011_),
    .Y(_10012_));
 sky130_fd_sc_hd__xnor2_4 _17268_ (.A(_10012_),
    .B(_09943_),
    .Y(net160));
 sky130_fd_sc_hd__maj3_2 _17269_ (.A(net1555),
    .B(_09792_),
    .C(_09758_),
    .X(_10013_));
 sky130_fd_sc_hd__xor2_4 _17270_ (.A(_09938_),
    .B(_10013_),
    .X(net159));
 sky130_fd_sc_hd__mux4_1 _17271_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[404] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[436] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[468] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[500] ),
    .S0(net379),
    .S1(net371),
    .X(_10014_));
 sky130_fd_sc_hd__mux4_1 _17272_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[148] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[180] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[212] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[244] ),
    .S0(net379),
    .S1(net371),
    .X(_10015_));
 sky130_fd_sc_hd__nand2b_1 _17273_ (.A_N(net337),
    .B(net339),
    .Y(_10016_));
 sky130_fd_sc_hd__o22ai_2 _17274_ (.A1(_09075_),
    .A2(_10014_),
    .B1(_10015_),
    .B2(_10016_),
    .Y(_10017_));
 sky130_fd_sc_hd__mux4_1 _17275_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[276] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[308] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[340] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[372] ),
    .S0(net379),
    .S1(net371),
    .X(_10018_));
 sky130_fd_sc_hd__nor3_1 _17276_ (.A(_08162_),
    .B(net339),
    .C(_10018_),
    .Y(_10019_));
 sky130_fd_sc_hd__inv_1 _17277_ (.A(\gen_regfile_ff.register_file_i.rf_reg[84] ),
    .Y(_10020_));
 sky130_fd_sc_hd__mux2i_2 _17278_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[52] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[116] ),
    .S(net356),
    .Y(_10021_));
 sky130_fd_sc_hd__nor2_1 _17279_ (.A(net337),
    .B(net342),
    .Y(_10022_));
 sky130_fd_sc_hd__o221ai_4 _17280_ (.A1(_10020_),
    .A2(_08142_),
    .B1(_10021_),
    .B2(_08658_),
    .C1(_10022_),
    .Y(_10023_));
 sky130_fd_sc_hd__nand4bb_4 _17281_ (.A_N(_10017_),
    .B_N(_10019_),
    .C(_10023_),
    .D(_08161_),
    .Y(_10024_));
 sky130_fd_sc_hd__mux2i_1 _17282_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[564] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[628] ),
    .S(net346),
    .Y(_10025_));
 sky130_fd_sc_hd__mux2i_1 _17283_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[660] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[724] ),
    .S(net346),
    .Y(_10026_));
 sky130_fd_sc_hd__a22oi_1 _17284_ (.A1(net889),
    .A2(_10025_),
    .B1(_10026_),
    .B2(net589),
    .Y(_10027_));
 sky130_fd_sc_hd__mux2i_1 _17285_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[532] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[596] ),
    .S(net346),
    .Y(_10028_));
 sky130_fd_sc_hd__mux2i_1 _17286_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[692] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[756] ),
    .S(net346),
    .Y(_10029_));
 sky130_fd_sc_hd__a22oi_1 _17287_ (.A1(net650),
    .A2(_10028_),
    .B1(_10029_),
    .B2(net1153),
    .Y(_10030_));
 sky130_fd_sc_hd__nand3_1 _17288_ (.A(net698),
    .B(_10027_),
    .C(_10030_),
    .Y(_10031_));
 sky130_fd_sc_hd__mux2i_1 _17289_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[788] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[852] ),
    .S(net346),
    .Y(_10032_));
 sky130_fd_sc_hd__nand2_1 _17290_ (.A(net650),
    .B(_10032_),
    .Y(_10033_));
 sky130_fd_sc_hd__mux2i_1 _17291_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[820] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[884] ),
    .S(net346),
    .Y(_10034_));
 sky130_fd_sc_hd__mux2i_1 _17292_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[916] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[980] ),
    .S(net346),
    .Y(_10035_));
 sky130_fd_sc_hd__a22oi_1 _17293_ (.A1(net890),
    .A2(_10034_),
    .B1(_10035_),
    .B2(net591),
    .Y(_10036_));
 sky130_fd_sc_hd__mux2i_1 _17294_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[948] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1012] ),
    .S(net346),
    .Y(_10037_));
 sky130_fd_sc_hd__a21oi_1 _17295_ (.A1(net1153),
    .A2(_10037_),
    .B1(_08708_),
    .Y(_10038_));
 sky130_fd_sc_hd__nand3_2 _17296_ (.A(_10033_),
    .B(_10036_),
    .C(_10038_),
    .Y(_10039_));
 sky130_fd_sc_hd__nand3_4 _17297_ (.A(_10024_),
    .B(_10031_),
    .C(_10039_),
    .Y(_10040_));
 sky130_fd_sc_hd__nand2_4 _17298_ (.A(net827),
    .B(_08449_),
    .Y(_10041_));
 sky130_fd_sc_hd__nand2_1 _17299_ (.A(net1133),
    .B(_09455_),
    .Y(_10042_));
 sky130_fd_sc_hd__a21oi_1 _17300_ (.A1(_10041_),
    .A2(_10042_),
    .B1(_08495_),
    .Y(_10043_));
 sky130_fd_sc_hd__a21oi_2 _17301_ (.A1(_08495_),
    .A2(_10040_),
    .B1(_10043_),
    .Y(_10044_));
 sky130_fd_sc_hd__xnor2_1 _17302_ (.A(net296),
    .B(_10044_),
    .Y(_10045_));
 sky130_fd_sc_hd__mux4_1 _17303_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[660] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[692] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[724] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[756] ),
    .S0(net420),
    .S1(net1009),
    .X(_10046_));
 sky130_fd_sc_hd__mux4_1 _17304_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[532] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[564] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[596] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[628] ),
    .S0(net420),
    .S1(net1009),
    .X(_10047_));
 sky130_fd_sc_hd__a22oi_2 _17305_ (.A1(net1247),
    .A2(_10046_),
    .B1(_10047_),
    .B2(_08342_),
    .Y(_10048_));
 sky130_fd_sc_hd__mux4_1 _17306_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[916] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[948] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[980] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1012] ),
    .S0(net418),
    .S1(net409),
    .X(_10049_));
 sky130_fd_sc_hd__mux4_1 _17307_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[788] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[820] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[852] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[884] ),
    .S0(net418),
    .S1(net409),
    .X(_10050_));
 sky130_fd_sc_hd__a22oi_2 _17308_ (.A1(_08324_),
    .A2(_10049_),
    .B1(_10050_),
    .B2(net330),
    .Y(_10051_));
 sky130_fd_sc_hd__nand3_2 _17309_ (.A(net386),
    .B(_10048_),
    .C(_10051_),
    .Y(_10052_));
 sky130_fd_sc_hd__mux4_1 _17310_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[148] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[180] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[212] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[244] ),
    .S0(net420),
    .S1(net412),
    .X(_10053_));
 sky130_fd_sc_hd__nor2_2 _17311_ (.A(_08529_),
    .B(_10053_),
    .Y(_10054_));
 sky130_fd_sc_hd__mux2_1 _17312_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[84] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[116] ),
    .S(net1147),
    .X(_10055_));
 sky130_fd_sc_hd__a221oi_4 _17313_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[52] ),
    .A2(_08321_),
    .B1(_10055_),
    .B2(net1072),
    .C1(net399),
    .Y(_10056_));
 sky130_fd_sc_hd__mux4_2 _17314_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[404] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[436] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[468] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[500] ),
    .S0(net420),
    .S1(net412),
    .X(_10057_));
 sky130_fd_sc_hd__mux4_1 _17315_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[276] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[308] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[340] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[372] ),
    .S0(net419),
    .S1(net1070),
    .X(_10058_));
 sky130_fd_sc_hd__a22oi_4 _17316_ (.A1(net565),
    .A2(_10057_),
    .B1(_10058_),
    .B2(net330),
    .Y(_10059_));
 sky130_fd_sc_hd__o311ai_4 _17317_ (.A1(net975),
    .A2(_10054_),
    .A3(_10056_),
    .B1(_10059_),
    .C1(_08512_),
    .Y(_10060_));
 sky130_fd_sc_hd__nand2_8 _17318_ (.A(_10052_),
    .B(_10060_),
    .Y(_10061_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_877 ();
 sky130_fd_sc_hd__o22ai_1 _17320_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[52] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[20] ),
    .B2(_08503_),
    .Y(_10063_));
 sky130_fd_sc_hd__nor2_1 _17321_ (.A(_08504_),
    .B(_10040_),
    .Y(_10064_));
 sky130_fd_sc_hd__a2111oi_1 _17322_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(_10061_),
    .B1(_10063_),
    .C1(_10064_),
    .D1(_08295_),
    .Y(_10065_));
 sky130_fd_sc_hd__a21oi_2 _17323_ (.A1(net1134),
    .A2(_10045_),
    .B1(_10065_),
    .Y(_10066_));
 sky130_fd_sc_hd__nor2_1 _17324_ (.A(net310),
    .B(_10061_),
    .Y(_10067_));
 sky130_fd_sc_hd__a21oi_1 _17325_ (.A1(\cs_registers_i.pc_id_i[20] ),
    .A2(net310),
    .B1(_10067_),
    .Y(_10068_));
 sky130_fd_sc_hd__nand2_1 _17326_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[20] ),
    .B(_08368_),
    .Y(_10069_));
 sky130_fd_sc_hd__o21ai_4 _17327_ (.A1(net933),
    .A2(_10068_),
    .B1(_10069_),
    .Y(_10070_));
 sky130_fd_sc_hd__nand2_1 _17328_ (.A(net739),
    .B(_10070_),
    .Y(_10071_));
 sky130_fd_sc_hd__nand3_1 _17329_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[52] ),
    .B(_08272_),
    .C(_08377_),
    .Y(_10072_));
 sky130_fd_sc_hd__nand2_1 _17330_ (.A(_10071_),
    .B(_10072_),
    .Y(_10073_));
 sky130_fd_sc_hd__xnor2_2 _17331_ (.A(_10066_),
    .B(_10073_),
    .Y(_10074_));
 sky130_fd_sc_hd__nor3_2 _17332_ (.A(_09939_),
    .B(_10012_),
    .C(_10074_),
    .Y(_10075_));
 sky130_fd_sc_hd__and2_0 _17333_ (.A(_09870_),
    .B(_10075_),
    .X(_10076_));
 sky130_fd_sc_hd__nand2_1 _17334_ (.A(_10004_),
    .B(_10011_),
    .Y(_10077_));
 sky130_fd_sc_hd__nor2_1 _17335_ (.A(_10004_),
    .B(_10011_),
    .Y(_10078_));
 sky130_fd_sc_hd__a21oi_1 _17336_ (.A1(_09942_),
    .A2(_10077_),
    .B1(_10078_),
    .Y(_10079_));
 sky130_fd_sc_hd__maj3_1 _17337_ (.A(_10066_),
    .B(_10073_),
    .C(_10079_),
    .X(_10080_));
 sky130_fd_sc_hd__a311o_4 _17338_ (.A1(_09651_),
    .A2(_09867_),
    .A3(_10075_),
    .B1(_10076_),
    .C1(_10080_),
    .X(_10081_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_874 ();
 sky130_fd_sc_hd__nand2_1 _17342_ (.A(net1141),
    .B(_09455_),
    .Y(_10085_));
 sky130_fd_sc_hd__mux4_2 _17343_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[149] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[181] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[213] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[245] ),
    .S0(net1029),
    .S1(net516),
    .X(_10086_));
 sky130_fd_sc_hd__mux2_1 _17344_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[53] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[117] ),
    .S(net1120),
    .X(_10087_));
 sky130_fd_sc_hd__a221o_1 _17345_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[85] ),
    .A2(net324),
    .B1(_10087_),
    .B2(net1476),
    .C1(net343),
    .X(_10088_));
 sky130_fd_sc_hd__o211ai_4 _17346_ (.A1(_08481_),
    .A2(_10086_),
    .B1(_10088_),
    .C1(_08731_),
    .Y(_10089_));
 sky130_fd_sc_hd__mux2i_1 _17347_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[309] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[373] ),
    .S(net347),
    .Y(_10090_));
 sky130_fd_sc_hd__mux2i_1 _17348_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[789] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[853] ),
    .S(net347),
    .Y(_10091_));
 sky130_fd_sc_hd__o22ai_2 _17349_ (.A1(net759),
    .A2(_10090_),
    .B1(_10091_),
    .B2(net508),
    .Y(_10092_));
 sky130_fd_sc_hd__mux2i_1 _17350_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[917] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[981] ),
    .S(net347),
    .Y(_10093_));
 sky130_fd_sc_hd__mux2i_1 _17351_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[821] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[885] ),
    .S(net347),
    .Y(_10094_));
 sky130_fd_sc_hd__o22ai_2 _17352_ (.A1(net601),
    .A2(_10093_),
    .B1(_10094_),
    .B2(net518),
    .Y(_10095_));
 sky130_fd_sc_hd__mux2i_1 _17353_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[949] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1013] ),
    .S(net347),
    .Y(_10096_));
 sky130_fd_sc_hd__mux2i_1 _17354_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[437] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[501] ),
    .S(net347),
    .Y(_10097_));
 sky130_fd_sc_hd__o22ai_2 _17355_ (.A1(net629),
    .A2(_10096_),
    .B1(_10097_),
    .B2(net870),
    .Y(_10098_));
 sky130_fd_sc_hd__mux2i_1 _17356_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[277] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[341] ),
    .S(net347),
    .Y(_10099_));
 sky130_fd_sc_hd__mux2i_1 _17357_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[405] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[469] ),
    .S(net347),
    .Y(_10100_));
 sky130_fd_sc_hd__o22ai_2 _17358_ (.A1(net772),
    .A2(_10099_),
    .B1(_10100_),
    .B2(net892),
    .Y(_10101_));
 sky130_fd_sc_hd__nor4_4 _17359_ (.A(_10092_),
    .B(_10101_),
    .C(_10098_),
    .D(_10095_),
    .Y(_10102_));
 sky130_fd_sc_hd__mux2i_1 _17360_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[661] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[725] ),
    .S(net347),
    .Y(_10103_));
 sky130_fd_sc_hd__mux2i_1 _17361_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[533] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[597] ),
    .S(net347),
    .Y(_10104_));
 sky130_fd_sc_hd__a22oi_2 _17362_ (.A1(net1013),
    .A2(_10103_),
    .B1(_10104_),
    .B2(net650),
    .Y(_10105_));
 sky130_fd_sc_hd__mux2i_1 _17363_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[565] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[629] ),
    .S(net347),
    .Y(_10106_));
 sky130_fd_sc_hd__mux2i_1 _17364_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[693] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[757] ),
    .S(net347),
    .Y(_10107_));
 sky130_fd_sc_hd__a22oi_2 _17365_ (.A1(net1201),
    .A2(_10106_),
    .B1(_10107_),
    .B2(net1153),
    .Y(_10108_));
 sky130_fd_sc_hd__nand3_4 _17366_ (.A(_08462_),
    .B(_10105_),
    .C(_10108_),
    .Y(_10109_));
 sky130_fd_sc_hd__nand3_4 _17367_ (.A(_10089_),
    .B(net1174),
    .C(_10109_),
    .Y(_10110_));
 sky130_fd_sc_hd__nor2_1 _17368_ (.A(_08436_),
    .B(_10110_),
    .Y(_10111_));
 sky130_fd_sc_hd__a31oi_4 _17369_ (.A1(_08436_),
    .A2(_10041_),
    .A3(_10085_),
    .B1(_10111_),
    .Y(_10112_));
 sky130_fd_sc_hd__xor2_1 _17370_ (.A(net296),
    .B(_10112_),
    .X(_10113_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_873 ();
 sky130_fd_sc_hd__mux4_2 _17372_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[661] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[693] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[725] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[757] ),
    .S0(net856),
    .S1(net405),
    .X(_10115_));
 sky130_fd_sc_hd__mux4_1 _17373_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[533] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[565] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[597] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[629] ),
    .S0(net856),
    .S1(net405),
    .X(_10116_));
 sky130_fd_sc_hd__a22oi_4 _17374_ (.A1(net610),
    .A2(_10115_),
    .B1(_10116_),
    .B2(_08342_),
    .Y(_10117_));
 sky130_fd_sc_hd__mux4_1 _17375_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[917] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[949] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[981] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1013] ),
    .S0(net1076),
    .S1(net405),
    .X(_10118_));
 sky130_fd_sc_hd__mux4_1 _17376_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[789] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[821] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[853] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[885] ),
    .S0(net856),
    .S1(net405),
    .X(_10119_));
 sky130_fd_sc_hd__a22oi_4 _17377_ (.A1(net565),
    .A2(_10118_),
    .B1(_10119_),
    .B2(net532),
    .Y(_10120_));
 sky130_fd_sc_hd__nand3_2 _17378_ (.A(net386),
    .B(_10117_),
    .C(_10120_),
    .Y(_10121_));
 sky130_fd_sc_hd__mux4_2 _17379_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[149] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[181] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[213] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[245] ),
    .S0(net752),
    .S1(net794),
    .X(_10122_));
 sky130_fd_sc_hd__nor2_2 _17380_ (.A(_08529_),
    .B(_10122_),
    .Y(_10123_));
 sky130_fd_sc_hd__mux2_1 _17381_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[85] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[117] ),
    .S(net1084),
    .X(_10124_));
 sky130_fd_sc_hd__a221oi_4 _17382_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[53] ),
    .A2(net544),
    .B1(_10124_),
    .B2(net413),
    .C1(net398),
    .Y(_10125_));
 sky130_fd_sc_hd__mux4_1 _17383_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[405] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[437] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[469] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[501] ),
    .S0(net1076),
    .S1(net405),
    .X(_10126_));
 sky130_fd_sc_hd__mux4_1 _17384_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[277] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[309] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[341] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[373] ),
    .S0(net1076),
    .S1(net405),
    .X(_10127_));
 sky130_fd_sc_hd__a22oi_4 _17385_ (.A1(_10126_),
    .A2(net565),
    .B1(_10127_),
    .B2(net532),
    .Y(_10128_));
 sky130_fd_sc_hd__o311ai_4 _17386_ (.A1(net1075),
    .A2(_10123_),
    .A3(_10125_),
    .B1(_10128_),
    .C1(_08512_),
    .Y(_10129_));
 sky130_fd_sc_hd__nand2_8 _17387_ (.A(_10121_),
    .B(_10129_),
    .Y(_10130_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_871 ();
 sky130_fd_sc_hd__o22ai_1 _17390_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[53] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[21] ),
    .B2(_08503_),
    .Y(_10133_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_870 ();
 sky130_fd_sc_hd__nor2_1 _17392_ (.A(_08504_),
    .B(_10110_),
    .Y(_10135_));
 sky130_fd_sc_hd__a2111oi_1 _17393_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(_10130_),
    .B1(_10133_),
    .C1(_10135_),
    .D1(net739),
    .Y(_10136_));
 sky130_fd_sc_hd__a21oi_2 _17394_ (.A1(net739),
    .A2(_10113_),
    .B1(_10136_),
    .Y(_10137_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_867 ();
 sky130_fd_sc_hd__nor2_1 _17398_ (.A(net310),
    .B(_10130_),
    .Y(_10141_));
 sky130_fd_sc_hd__a21oi_1 _17399_ (.A1(\cs_registers_i.pc_id_i[21] ),
    .A2(net310),
    .B1(_10141_),
    .Y(_10142_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_866 ();
 sky130_fd_sc_hd__nand2_1 _17401_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[21] ),
    .B(_08368_),
    .Y(_10144_));
 sky130_fd_sc_hd__o21ai_4 _17402_ (.A1(net933),
    .A2(_10142_),
    .B1(_10144_),
    .Y(_10145_));
 sky130_fd_sc_hd__nand2_1 _17403_ (.A(net739),
    .B(_10145_),
    .Y(_10146_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_865 ();
 sky130_fd_sc_hd__nand3_1 _17405_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[53] ),
    .B(_08272_),
    .C(_08377_),
    .Y(_10148_));
 sky130_fd_sc_hd__nand2_2 _17406_ (.A(_10146_),
    .B(_10148_),
    .Y(_10149_));
 sky130_fd_sc_hd__xnor2_2 _17407_ (.A(_10137_),
    .B(_10149_),
    .Y(_10150_));
 sky130_fd_sc_hd__xnor2_4 _17408_ (.A(_10150_),
    .B(_10081_),
    .Y(net162));
 sky130_fd_sc_hd__maj3_2 _17409_ (.A(_09943_),
    .B(_10004_),
    .C(_10011_),
    .X(_10151_));
 sky130_fd_sc_hd__xnor2_4 _17410_ (.A(_10151_),
    .B(_10074_),
    .Y(net161));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_864 ();
 sky130_fd_sc_hd__mux4_1 _17412_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[662] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[694] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[726] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[758] ),
    .S0(net418),
    .S1(net1233),
    .X(_10153_));
 sky130_fd_sc_hd__mux4_1 _17413_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[534] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[566] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[598] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[630] ),
    .S0(net418),
    .S1(net1233),
    .X(_10154_));
 sky130_fd_sc_hd__a22oi_4 _17414_ (.A1(net1247),
    .A2(_10153_),
    .B1(_10154_),
    .B2(_08342_),
    .Y(_10155_));
 sky130_fd_sc_hd__mux4_2 _17415_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[918] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[950] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[982] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1014] ),
    .S0(net419),
    .S1(net412),
    .X(_10156_));
 sky130_fd_sc_hd__mux4_1 _17416_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[790] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[822] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[854] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[886] ),
    .S0(net416),
    .S1(net1070),
    .X(_10157_));
 sky130_fd_sc_hd__a22oi_4 _17417_ (.A1(net1248),
    .A2(_10156_),
    .B1(_10157_),
    .B2(net330),
    .Y(_10158_));
 sky130_fd_sc_hd__nand3_2 _17418_ (.A(net386),
    .B(_10155_),
    .C(_10158_),
    .Y(_10159_));
 sky130_fd_sc_hd__mux4_2 _17419_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[150] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[182] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[214] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[246] ),
    .S0(net989),
    .S1(net794),
    .X(_10160_));
 sky130_fd_sc_hd__nor2_2 _17420_ (.A(_08529_),
    .B(_10160_),
    .Y(_10161_));
 sky130_fd_sc_hd__mux2_1 _17421_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[86] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[118] ),
    .S(net989),
    .X(_10162_));
 sky130_fd_sc_hd__a221oi_4 _17422_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[54] ),
    .A2(net543),
    .B1(_10162_),
    .B2(net413),
    .C1(net400),
    .Y(_10163_));
 sky130_fd_sc_hd__mux4_2 _17423_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[406] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[438] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[470] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[502] ),
    .S0(net419),
    .S1(net412),
    .X(_10164_));
 sky130_fd_sc_hd__mux4_1 _17424_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[278] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[310] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[342] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[374] ),
    .S0(net416),
    .S1(net1070),
    .X(_10165_));
 sky130_fd_sc_hd__a22oi_4 _17425_ (.A1(net565),
    .A2(_10164_),
    .B1(_10165_),
    .B2(net330),
    .Y(_10166_));
 sky130_fd_sc_hd__o311ai_4 _17426_ (.A1(net976),
    .A2(_10161_),
    .A3(_10163_),
    .B1(_10166_),
    .C1(_08512_),
    .Y(_10167_));
 sky130_fd_sc_hd__nand2_8 _17427_ (.A(_10159_),
    .B(_10167_),
    .Y(_10168_));
 sky130_fd_sc_hd__nor2_1 _17428_ (.A(net310),
    .B(_10168_),
    .Y(_10169_));
 sky130_fd_sc_hd__a21oi_1 _17429_ (.A1(\cs_registers_i.pc_id_i[22] ),
    .A2(net310),
    .B1(_10169_),
    .Y(_10170_));
 sky130_fd_sc_hd__nand2_1 _17430_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[22] ),
    .B(_08368_),
    .Y(_10171_));
 sky130_fd_sc_hd__o21ai_4 _17431_ (.A1(net933),
    .A2(_10170_),
    .B1(_10171_),
    .Y(_10172_));
 sky130_fd_sc_hd__nand2_1 _17432_ (.A(net739),
    .B(_10172_),
    .Y(_10173_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_863 ();
 sky130_fd_sc_hd__nand3_1 _17434_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[54] ),
    .B(_08272_),
    .C(_08377_),
    .Y(_10175_));
 sky130_fd_sc_hd__nand2_1 _17435_ (.A(_10173_),
    .B(_10175_),
    .Y(_10176_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_862 ();
 sky130_fd_sc_hd__mux4_1 _17437_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[150] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[182] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[214] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[246] ),
    .S0(net380),
    .S1(net1142),
    .X(_10178_));
 sky130_fd_sc_hd__mux2_1 _17438_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[54] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[118] ),
    .S(net1142),
    .X(_10179_));
 sky130_fd_sc_hd__a221o_1 _17439_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[86] ),
    .A2(_08484_),
    .B1(_10179_),
    .B2(net1476),
    .C1(net343),
    .X(_10180_));
 sky130_fd_sc_hd__o211ai_4 _17440_ (.A1(_08481_),
    .A2(_10178_),
    .B1(_10180_),
    .C1(_08731_),
    .Y(_10181_));
 sky130_fd_sc_hd__mux2i_1 _17441_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[662] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[726] ),
    .S(net346),
    .Y(_10182_));
 sky130_fd_sc_hd__mux2i_1 _17442_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[534] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[598] ),
    .S(net345),
    .Y(_10183_));
 sky130_fd_sc_hd__a22oi_1 _17443_ (.A1(net589),
    .A2(_10182_),
    .B1(_10183_),
    .B2(net650),
    .Y(_10184_));
 sky130_fd_sc_hd__mux2i_1 _17444_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[566] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[630] ),
    .S(net345),
    .Y(_10185_));
 sky130_fd_sc_hd__mux2i_1 _17445_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[694] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[758] ),
    .S(net346),
    .Y(_10186_));
 sky130_fd_sc_hd__a22oi_1 _17446_ (.A1(net889),
    .A2(_10185_),
    .B1(_10186_),
    .B2(net1153),
    .Y(_10187_));
 sky130_fd_sc_hd__nand3_2 _17447_ (.A(net698),
    .B(_10184_),
    .C(_10187_),
    .Y(_10188_));
 sky130_fd_sc_hd__mux2i_1 _17448_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[950] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1014] ),
    .S(net369),
    .Y(_10189_));
 sky130_fd_sc_hd__mux2i_1 _17449_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[310] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[374] ),
    .S(net370),
    .Y(_10190_));
 sky130_fd_sc_hd__o22ai_2 _17450_ (.A1(net634),
    .A2(_10189_),
    .B1(_10190_),
    .B2(net765),
    .Y(_10191_));
 sky130_fd_sc_hd__mux2i_1 _17451_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[438] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[502] ),
    .S(net369),
    .Y(_10192_));
 sky130_fd_sc_hd__mux2i_1 _17452_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[406] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[470] ),
    .S(net369),
    .Y(_10193_));
 sky130_fd_sc_hd__o22ai_2 _17453_ (.A1(net869),
    .A2(_10192_),
    .B1(_10193_),
    .B2(net897),
    .Y(_10194_));
 sky130_fd_sc_hd__mux2i_1 _17454_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[790] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[854] ),
    .S(net370),
    .Y(_10195_));
 sky130_fd_sc_hd__mux2i_1 _17455_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[822] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[886] ),
    .S(net370),
    .Y(_10196_));
 sky130_fd_sc_hd__o22ai_2 _17456_ (.A1(net501),
    .A2(_10195_),
    .B1(_10196_),
    .B2(net523),
    .Y(_10197_));
 sky130_fd_sc_hd__mux2i_1 _17457_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[278] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[342] ),
    .S(net370),
    .Y(_10198_));
 sky130_fd_sc_hd__mux2i_1 _17458_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[918] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[982] ),
    .S(net369),
    .Y(_10199_));
 sky130_fd_sc_hd__o22ai_2 _17459_ (.A1(net807),
    .A2(_10198_),
    .B1(_10199_),
    .B2(net606),
    .Y(_10200_));
 sky130_fd_sc_hd__nor4_4 _17460_ (.A(_10200_),
    .B(_10194_),
    .C(_10197_),
    .D(_10191_),
    .Y(_10201_));
 sky130_fd_sc_hd__nand3_4 _17461_ (.A(_10181_),
    .B(_10188_),
    .C(net1218),
    .Y(_10202_));
 sky130_fd_sc_hd__nand2_1 _17462_ (.A(net341),
    .B(_09455_),
    .Y(_10203_));
 sky130_fd_sc_hd__a21oi_1 _17463_ (.A1(_10041_),
    .A2(_10203_),
    .B1(_08495_),
    .Y(_10204_));
 sky130_fd_sc_hd__a21oi_2 _17464_ (.A1(_08495_),
    .A2(_10202_),
    .B1(_10204_),
    .Y(_10205_));
 sky130_fd_sc_hd__xnor2_1 _17465_ (.A(net296),
    .B(_10205_),
    .Y(_10206_));
 sky130_fd_sc_hd__nor2_1 _17466_ (.A(_08504_),
    .B(_10202_),
    .Y(_10207_));
 sky130_fd_sc_hd__o22ai_1 _17467_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[54] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[22] ),
    .B2(_08503_),
    .Y(_10208_));
 sky130_fd_sc_hd__a2111oi_1 _17468_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(_10168_),
    .B1(_10207_),
    .C1(_10208_),
    .D1(net739),
    .Y(_10209_));
 sky130_fd_sc_hd__a21oi_2 _17469_ (.A1(net739),
    .A2(_10206_),
    .B1(_10209_),
    .Y(_10210_));
 sky130_fd_sc_hd__nor2_1 _17470_ (.A(_10176_),
    .B(_10210_),
    .Y(_10211_));
 sky130_fd_sc_hd__nor2_1 _17471_ (.A(_10137_),
    .B(_10149_),
    .Y(_10212_));
 sky130_fd_sc_hd__nor2_1 _17472_ (.A(_10211_),
    .B(_10212_),
    .Y(_10213_));
 sky130_fd_sc_hd__a22oi_1 _17473_ (.A1(_10137_),
    .A2(_10149_),
    .B1(_10176_),
    .B2(_10210_),
    .Y(_10214_));
 sky130_fd_sc_hd__nor2_1 _17474_ (.A(_10211_),
    .B(_10214_),
    .Y(_10215_));
 sky130_fd_sc_hd__a21oi_4 _17475_ (.A1(_10081_),
    .A2(_10213_),
    .B1(_10215_),
    .Y(_10216_));
 sky130_fd_sc_hd__mux4_1 _17476_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[663] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[695] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[727] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[759] ),
    .S0(net417),
    .S1(net409),
    .X(_10217_));
 sky130_fd_sc_hd__mux4_1 _17477_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[535] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[567] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[599] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[631] ),
    .S0(net417),
    .S1(net409),
    .X(_10218_));
 sky130_fd_sc_hd__a22oi_4 _17478_ (.A1(net610),
    .A2(_10217_),
    .B1(_10218_),
    .B2(_08342_),
    .Y(_10219_));
 sky130_fd_sc_hd__mux4_1 _17479_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[919] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[951] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[983] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1015] ),
    .S0(net416),
    .S1(net404),
    .X(_10220_));
 sky130_fd_sc_hd__mux4_1 _17480_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[791] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[823] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[855] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[887] ),
    .S0(net416),
    .S1(net404),
    .X(_10221_));
 sky130_fd_sc_hd__a22oi_4 _17481_ (.A1(_10220_),
    .A2(net1248),
    .B1(_10221_),
    .B2(net531),
    .Y(_10222_));
 sky130_fd_sc_hd__nand3_2 _17482_ (.A(net386),
    .B(_10219_),
    .C(net1314),
    .Y(_10223_));
 sky130_fd_sc_hd__mux4_2 _17483_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[151] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[183] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[215] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[247] ),
    .S0(net752),
    .S1(net794),
    .X(_10224_));
 sky130_fd_sc_hd__nor2_2 _17484_ (.A(_08529_),
    .B(_10224_),
    .Y(_10225_));
 sky130_fd_sc_hd__mux2_1 _17485_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[87] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[119] ),
    .S(net1130),
    .X(_10226_));
 sky130_fd_sc_hd__a221oi_4 _17486_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[55] ),
    .A2(net544),
    .B1(_10226_),
    .B2(net413),
    .C1(net400),
    .Y(_10227_));
 sky130_fd_sc_hd__mux4_1 _17487_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[407] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[439] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[471] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[503] ),
    .S0(net416),
    .S1(net1113),
    .X(_10228_));
 sky130_fd_sc_hd__mux4_1 _17488_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[279] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[311] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[343] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[375] ),
    .S0(net416),
    .S1(net1070),
    .X(_10229_));
 sky130_fd_sc_hd__a22oi_4 _17489_ (.A1(_10228_),
    .A2(net1248),
    .B1(_10229_),
    .B2(net530),
    .Y(_10230_));
 sky130_fd_sc_hd__o311ai_4 _17490_ (.A1(net1075),
    .A2(_10225_),
    .A3(_10227_),
    .B1(_10230_),
    .C1(_08512_),
    .Y(_10231_));
 sky130_fd_sc_hd__nand2_8 _17491_ (.A(_10223_),
    .B(_10231_),
    .Y(_10232_));
 sky130_fd_sc_hd__inv_1 _17492_ (.A(_10232_),
    .Y(_10233_));
 sky130_fd_sc_hd__mux2i_1 _17493_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[535] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[599] ),
    .S(net344),
    .Y(_10234_));
 sky130_fd_sc_hd__nand2_1 _17494_ (.A(net650),
    .B(_10234_),
    .Y(_10235_));
 sky130_fd_sc_hd__mux2i_1 _17495_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[663] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[727] ),
    .S(net344),
    .Y(_10236_));
 sky130_fd_sc_hd__mux2i_1 _17496_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[567] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[631] ),
    .S(net344),
    .Y(_10237_));
 sky130_fd_sc_hd__a22oi_2 _17497_ (.A1(net1013),
    .A2(_10236_),
    .B1(_10237_),
    .B2(net1201),
    .Y(_10238_));
 sky130_fd_sc_hd__mux2i_1 _17498_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[695] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[759] ),
    .S(net344),
    .Y(_10239_));
 sky130_fd_sc_hd__a21oi_1 _17499_ (.A1(net1153),
    .A2(_10239_),
    .B1(_08679_),
    .Y(_10240_));
 sky130_fd_sc_hd__nand3_4 _17500_ (.A(_10235_),
    .B(_10238_),
    .C(_10240_),
    .Y(_10241_));
 sky130_fd_sc_hd__mux2i_1 _17501_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[951] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1015] ),
    .S(net368),
    .Y(_10242_));
 sky130_fd_sc_hd__mux2i_1 _17502_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[439] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[503] ),
    .S(net368),
    .Y(_10243_));
 sky130_fd_sc_hd__o22ai_2 _17503_ (.A1(net635),
    .A2(_10242_),
    .B1(_10243_),
    .B2(net867),
    .Y(_10244_));
 sky130_fd_sc_hd__mux2i_1 _17504_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[279] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[343] ),
    .S(net368),
    .Y(_10245_));
 sky130_fd_sc_hd__mux2i_1 _17505_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[311] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[375] ),
    .S(net368),
    .Y(_10246_));
 sky130_fd_sc_hd__o22ai_4 _17506_ (.A1(net771),
    .A2(_10245_),
    .B1(_10246_),
    .B2(net766),
    .Y(_10247_));
 sky130_fd_sc_hd__mux2i_1 _17507_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[919] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[983] ),
    .S(net368),
    .Y(_10248_));
 sky130_fd_sc_hd__mux2i_1 _17508_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[791] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[855] ),
    .S(net368),
    .Y(_10249_));
 sky130_fd_sc_hd__o22ai_2 _17509_ (.A1(net607),
    .A2(_10248_),
    .B1(_10249_),
    .B2(net505),
    .Y(_10250_));
 sky130_fd_sc_hd__mux2i_1 _17510_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[823] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[887] ),
    .S(net368),
    .Y(_10251_));
 sky130_fd_sc_hd__mux2i_2 _17511_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[407] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[471] ),
    .S(net368),
    .Y(_10252_));
 sky130_fd_sc_hd__o22ai_2 _17512_ (.A1(net526),
    .A2(_10251_),
    .B1(_10252_),
    .B2(net896),
    .Y(_10253_));
 sky130_fd_sc_hd__nor4_4 _17513_ (.A(_10250_),
    .B(_10247_),
    .C(_10244_),
    .D(_10253_),
    .Y(_10254_));
 sky130_fd_sc_hd__mux4_2 _17514_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[151] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[183] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[215] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[247] ),
    .S0(net1029),
    .S1(net515),
    .X(_10255_));
 sky130_fd_sc_hd__mux2_1 _17515_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[55] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[119] ),
    .S(net1120),
    .X(_10256_));
 sky130_fd_sc_hd__a221o_1 _17516_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[87] ),
    .A2(net324),
    .B1(_10256_),
    .B2(net1476),
    .C1(net343),
    .X(_10257_));
 sky130_fd_sc_hd__o211ai_4 _17517_ (.A1(_08481_),
    .A2(_10255_),
    .B1(_10257_),
    .C1(_08731_),
    .Y(_10258_));
 sky130_fd_sc_hd__nand3_4 _17518_ (.A(_10241_),
    .B(net743),
    .C(_10258_),
    .Y(_10259_));
 sky130_fd_sc_hd__nor2_1 _17519_ (.A(_08504_),
    .B(_10259_),
    .Y(_10260_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_861 ();
 sky130_fd_sc_hd__o22ai_1 _17521_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[55] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[23] ),
    .B2(_08503_),
    .Y(_10262_));
 sky130_fd_sc_hd__nor2_1 _17522_ (.A(_10260_),
    .B(_10262_),
    .Y(_10263_));
 sky130_fd_sc_hd__o21ai_2 _17523_ (.A1(_08500_),
    .A2(_10233_),
    .B1(_10263_),
    .Y(_10264_));
 sky130_fd_sc_hd__a221o_1 _17524_ (.A1(net827),
    .A2(_08449_),
    .B1(_09455_),
    .B2(net546),
    .C1(_08495_),
    .X(_10265_));
 sky130_fd_sc_hd__o21ai_4 _17525_ (.A1(_10259_),
    .A2(_08436_),
    .B1(_10265_),
    .Y(_10266_));
 sky130_fd_sc_hd__xnor2_2 _17526_ (.A(net297),
    .B(_10266_),
    .Y(_10267_));
 sky130_fd_sc_hd__nor2_1 _17527_ (.A(net313),
    .B(_10267_),
    .Y(_10268_));
 sky130_fd_sc_hd__a21oi_4 _17528_ (.A1(_08272_),
    .A2(_10264_),
    .B1(_10268_),
    .Y(_10269_));
 sky130_fd_sc_hd__nor2_1 _17529_ (.A(net310),
    .B(_10232_),
    .Y(_10270_));
 sky130_fd_sc_hd__a21oi_1 _17530_ (.A1(\cs_registers_i.pc_id_i[23] ),
    .A2(net310),
    .B1(_10270_),
    .Y(_10271_));
 sky130_fd_sc_hd__a2bb2oi_4 _17531_ (.A1_N(_10271_),
    .A2_N(net933),
    .B1(_08368_),
    .B2(\id_stage_i.controller_i.lsu_addr_last_i[23] ),
    .Y(_10272_));
 sky130_fd_sc_hd__nor2_1 _17532_ (.A(net313),
    .B(_10272_),
    .Y(_10273_));
 sky130_fd_sc_hd__a31oi_4 _17533_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[55] ),
    .A2(_08272_),
    .A3(_08377_),
    .B1(_10273_),
    .Y(_10274_));
 sky130_fd_sc_hd__xor2_4 _17534_ (.A(_10269_),
    .B(_10274_),
    .X(_10275_));
 sky130_fd_sc_hd__xnor2_4 _17535_ (.A(_10275_),
    .B(net656),
    .Y(net164));
 sky130_fd_sc_hd__maj3_2 _17536_ (.A(_10081_),
    .B(_10137_),
    .C(_10149_),
    .X(_10276_));
 sky130_fd_sc_hd__xnor2_2 _17537_ (.A(_10176_),
    .B(_10210_),
    .Y(_10277_));
 sky130_fd_sc_hd__xnor2_4 _17538_ (.A(_10276_),
    .B(_10277_),
    .Y(net163));
 sky130_fd_sc_hd__mux2_1 _17539_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[217] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[249] ),
    .S(net1084),
    .X(_10278_));
 sky130_fd_sc_hd__mux2_1 _17540_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[89] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[121] ),
    .S(net436),
    .X(_10279_));
 sky130_fd_sc_hd__o22ai_2 _17541_ (.A1(_08815_),
    .A2(_10278_),
    .B1(_10279_),
    .B2(_08819_),
    .Y(_10280_));
 sky130_fd_sc_hd__mux2_1 _17542_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[153] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[185] ),
    .S(net1084),
    .X(_10281_));
 sky130_fd_sc_hd__a221oi_2 _17543_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[57] ),
    .A2(_09530_),
    .B1(_10281_),
    .B2(net398),
    .C1(net402),
    .Y(_10282_));
 sky130_fd_sc_hd__o21ai_4 _17544_ (.A1(_10280_),
    .A2(_10282_),
    .B1(_08179_),
    .Y(_10283_));
 sky130_fd_sc_hd__mux2_1 _17545_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[793] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[825] ),
    .S(net799),
    .X(_10284_));
 sky130_fd_sc_hd__nand2b_1 _17546_ (.A_N(\gen_regfile_ff.register_file_i.rf_reg[889] ),
    .B(net799),
    .Y(_10285_));
 sky130_fd_sc_hd__o221ai_2 _17547_ (.A1(net799),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[857] ),
    .B1(_10284_),
    .B2(net1083),
    .C1(_10285_),
    .Y(_10286_));
 sky130_fd_sc_hd__mux2_1 _17548_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[921] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[953] ),
    .S(net799),
    .X(_10287_));
 sky130_fd_sc_hd__mux2_1 _17549_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[985] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1017] ),
    .S(net799),
    .X(_10288_));
 sky130_fd_sc_hd__o211ai_2 _17550_ (.A1(net1083),
    .A2(_10287_),
    .B1(_10288_),
    .C1(net393),
    .Y(_10289_));
 sky130_fd_sc_hd__a221oi_2 _17551_ (.A1(net623),
    .A2(_10287_),
    .B1(_10284_),
    .B2(net649),
    .C1(_08809_),
    .Y(_10290_));
 sky130_fd_sc_hd__o211ai_4 _17552_ (.A1(net393),
    .A2(_10286_),
    .B1(_10289_),
    .C1(_10290_),
    .Y(_10291_));
 sky130_fd_sc_hd__mux4_4 _17553_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[665] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[697] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[729] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[761] ),
    .S0(net856),
    .S1(net405),
    .X(_10292_));
 sky130_fd_sc_hd__mux4_4 _17554_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[537] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[569] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[601] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[633] ),
    .S0(net856),
    .S1(net405),
    .X(_10293_));
 sky130_fd_sc_hd__o22ai_1 _17555_ (.A1(_09279_),
    .A2(_10292_),
    .B1(_10293_),
    .B2(_09550_),
    .Y(_10294_));
 sky130_fd_sc_hd__mux4_1 _17556_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[345] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[377] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[473] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[505] ),
    .S0(net799),
    .S1(net393),
    .X(_10295_));
 sky130_fd_sc_hd__mux4_2 _17557_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[281] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[313] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[409] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[441] ),
    .S0(net799),
    .S1(net393),
    .X(_10296_));
 sky130_fd_sc_hd__o22ai_1 _17558_ (.A1(_09543_),
    .A2(_10295_),
    .B1(_10296_),
    .B2(_09546_),
    .Y(_10297_));
 sky130_fd_sc_hd__nor2_2 _17559_ (.A(_10294_),
    .B(_10297_),
    .Y(_10298_));
 sky130_fd_sc_hd__nand3_4 _17560_ (.A(_10283_),
    .B(_10291_),
    .C(_10298_),
    .Y(_10299_));
 sky130_fd_sc_hd__nor2_1 _17561_ (.A(net310),
    .B(_10299_),
    .Y(_10300_));
 sky130_fd_sc_hd__a21oi_1 _17562_ (.A1(\cs_registers_i.pc_id_i[25] ),
    .A2(net310),
    .B1(_10300_),
    .Y(_10301_));
 sky130_fd_sc_hd__nor2_1 _17563_ (.A(net933),
    .B(_10301_),
    .Y(_10302_));
 sky130_fd_sc_hd__a21oi_4 _17564_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[25] ),
    .A2(_08368_),
    .B1(_10302_),
    .Y(_10303_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_860 ();
 sky130_fd_sc_hd__a21oi_1 _17566_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[57] ),
    .A2(_08377_),
    .B1(net739),
    .Y(_10305_));
 sky130_fd_sc_hd__a21oi_4 _17567_ (.A1(net739),
    .A2(_10303_),
    .B1(_10305_),
    .Y(_10306_));
 sky130_fd_sc_hd__mux2_1 _17568_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[57] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[121] ),
    .S(net365),
    .X(_10307_));
 sky130_fd_sc_hd__a221oi_1 _17569_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[89] ),
    .A2(net324),
    .B1(_10307_),
    .B2(net983),
    .C1(net343),
    .Y(_10308_));
 sky130_fd_sc_hd__mux4_1 _17570_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[153] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[185] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[217] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[249] ),
    .S0(net375),
    .S1(net1077),
    .X(_10309_));
 sky130_fd_sc_hd__o21ai_0 _17571_ (.A1(_08481_),
    .A2(_10309_),
    .B1(_08731_),
    .Y(_10310_));
 sky130_fd_sc_hd__nor2_2 _17572_ (.A(_10308_),
    .B(_10310_),
    .Y(_10311_));
 sky130_fd_sc_hd__mux2i_1 _17573_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[569] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[633] ),
    .S(net349),
    .Y(_10312_));
 sky130_fd_sc_hd__mux2i_1 _17574_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[665] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[729] ),
    .S(net349),
    .Y(_10313_));
 sky130_fd_sc_hd__a22oi_2 _17575_ (.A1(net1201),
    .A2(_10312_),
    .B1(_10313_),
    .B2(net1013),
    .Y(_10314_));
 sky130_fd_sc_hd__mux2i_1 _17576_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[537] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[601] ),
    .S(net349),
    .Y(_10315_));
 sky130_fd_sc_hd__mux2i_1 _17577_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[697] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[761] ),
    .S(net349),
    .Y(_10316_));
 sky130_fd_sc_hd__a22oi_2 _17578_ (.A1(net650),
    .A2(_10315_),
    .B1(_10316_),
    .B2(net1153),
    .Y(_10317_));
 sky130_fd_sc_hd__nand3_4 _17579_ (.A(net698),
    .B(_10314_),
    .C(_10317_),
    .Y(_10318_));
 sky130_fd_sc_hd__mux2i_1 _17580_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[825] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[889] ),
    .S(net354),
    .Y(_10319_));
 sky130_fd_sc_hd__mux2i_1 _17581_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[313] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[377] ),
    .S(net1312),
    .Y(_10320_));
 sky130_fd_sc_hd__o22ai_2 _17582_ (.A1(net520),
    .A2(_10319_),
    .B1(_10320_),
    .B2(net761),
    .Y(_10321_));
 sky130_fd_sc_hd__mux2i_1 _17583_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[281] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[345] ),
    .S(net1312),
    .Y(_10322_));
 sky130_fd_sc_hd__mux2i_1 _17584_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[921] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[985] ),
    .S(net1312),
    .Y(_10323_));
 sky130_fd_sc_hd__o22ai_2 _17585_ (.A1(net772),
    .A2(_10322_),
    .B1(_10323_),
    .B2(net603),
    .Y(_10324_));
 sky130_fd_sc_hd__mux2i_1 _17586_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[953] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1017] ),
    .S(net354),
    .Y(_10325_));
 sky130_fd_sc_hd__mux2i_1 _17587_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[793] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[857] ),
    .S(net354),
    .Y(_10326_));
 sky130_fd_sc_hd__o22ai_2 _17588_ (.A1(net630),
    .A2(_10325_),
    .B1(_10326_),
    .B2(net509),
    .Y(_10327_));
 sky130_fd_sc_hd__mux2i_1 _17589_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[441] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[505] ),
    .S(net352),
    .Y(_10328_));
 sky130_fd_sc_hd__mux2i_1 _17590_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[409] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[473] ),
    .S(net352),
    .Y(_10329_));
 sky130_fd_sc_hd__o22ai_2 _17591_ (.A1(net872),
    .A2(_10328_),
    .B1(_10329_),
    .B2(net893),
    .Y(_10330_));
 sky130_fd_sc_hd__nor4_4 _17592_ (.A(_10330_),
    .B(_10324_),
    .C(_10321_),
    .D(_10327_),
    .Y(_10331_));
 sky130_fd_sc_hd__nand3b_4 _17593_ (.A_N(_10311_),
    .B(_10318_),
    .C(net937),
    .Y(_10332_));
 sky130_fd_sc_hd__nand2_1 _17594_ (.A(net582),
    .B(_09455_),
    .Y(_10333_));
 sky130_fd_sc_hd__a21oi_1 _17595_ (.A1(_10041_),
    .A2(_10333_),
    .B1(_08495_),
    .Y(_10334_));
 sky130_fd_sc_hd__a21oi_4 _17596_ (.A1(_08495_),
    .A2(_10332_),
    .B1(_10334_),
    .Y(_10335_));
 sky130_fd_sc_hd__xnor2_4 _17597_ (.A(net297),
    .B(_10335_),
    .Y(_10336_));
 sky130_fd_sc_hd__nor2_1 _17598_ (.A(_08504_),
    .B(_10332_),
    .Y(_10337_));
 sky130_fd_sc_hd__o22ai_1 _17599_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[57] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[25] ),
    .B2(_08503_),
    .Y(_10338_));
 sky130_fd_sc_hd__a2111oi_2 _17600_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(_10299_),
    .B1(_10337_),
    .C1(_10338_),
    .D1(net739),
    .Y(_10339_));
 sky130_fd_sc_hd__a21oi_4 _17601_ (.A1(net739),
    .A2(_10336_),
    .B1(_10339_),
    .Y(_10340_));
 sky130_fd_sc_hd__xnor2_2 _17602_ (.A(_10306_),
    .B(_10340_),
    .Y(_10341_));
 sky130_fd_sc_hd__clkinv_2 _17603_ (.A(_10341_),
    .Y(_10342_));
 sky130_fd_sc_hd__inv_2 _17604_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[56] ),
    .Y(_10343_));
 sky130_fd_sc_hd__mux2_1 _17605_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[216] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[248] ),
    .S(net1111),
    .X(_10344_));
 sky130_fd_sc_hd__mux2_1 _17606_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[88] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[120] ),
    .S(net1111),
    .X(_10345_));
 sky130_fd_sc_hd__o22ai_2 _17607_ (.A1(_08815_),
    .A2(_10344_),
    .B1(_10345_),
    .B2(_08819_),
    .Y(_10346_));
 sky130_fd_sc_hd__mux2_1 _17608_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[152] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[184] ),
    .S(net1111),
    .X(_10347_));
 sky130_fd_sc_hd__a221oi_2 _17609_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[56] ),
    .A2(_09530_),
    .B1(_10347_),
    .B2(net397),
    .C1(net403),
    .Y(_10348_));
 sky130_fd_sc_hd__o21ai_4 _17610_ (.A1(_10346_),
    .A2(_10348_),
    .B1(_08179_),
    .Y(_10349_));
 sky130_fd_sc_hd__mux2_1 _17611_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[792] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[824] ),
    .S(net1080),
    .X(_10350_));
 sky130_fd_sc_hd__nand2b_1 _17612_ (.A_N(\gen_regfile_ff.register_file_i.rf_reg[888] ),
    .B(net865),
    .Y(_10351_));
 sky130_fd_sc_hd__o221ai_2 _17613_ (.A1(net865),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[856] ),
    .B1(_10350_),
    .B2(net1009),
    .C1(_10351_),
    .Y(_10352_));
 sky130_fd_sc_hd__mux2_1 _17614_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[920] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[952] ),
    .S(net1080),
    .X(_10353_));
 sky130_fd_sc_hd__mux2_1 _17615_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[984] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1016] ),
    .S(net865),
    .X(_10354_));
 sky130_fd_sc_hd__o211ai_2 _17616_ (.A1(net1009),
    .A2(_10353_),
    .B1(_10354_),
    .C1(net394),
    .Y(_10355_));
 sky130_fd_sc_hd__a221oi_2 _17617_ (.A1(net1149),
    .A2(_10353_),
    .B1(_10350_),
    .B2(net649),
    .C1(_08809_),
    .Y(_10356_));
 sky130_fd_sc_hd__o211ai_4 _17618_ (.A1(net399),
    .A2(_10352_),
    .B1(_10355_),
    .C1(_10356_),
    .Y(_10357_));
 sky130_fd_sc_hd__mux4_1 _17619_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[664] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[696] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[728] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[760] ),
    .S0(net1080),
    .S1(net1083),
    .X(_10358_));
 sky130_fd_sc_hd__mux4_1 _17620_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[536] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[568] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[600] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[632] ),
    .S0(net1080),
    .S1(net1083),
    .X(_10359_));
 sky130_fd_sc_hd__o22ai_2 _17621_ (.A1(_09279_),
    .A2(_10358_),
    .B1(_10359_),
    .B2(_09550_),
    .Y(_10360_));
 sky130_fd_sc_hd__mux4_1 _17622_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[344] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[376] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[472] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[504] ),
    .S0(net989),
    .S1(net399),
    .X(_10361_));
 sky130_fd_sc_hd__mux4_1 _17623_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[280] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[312] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[408] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[440] ),
    .S0(net963),
    .S1(net399),
    .X(_10362_));
 sky130_fd_sc_hd__o22ai_2 _17624_ (.A1(_09543_),
    .A2(_10361_),
    .B1(_10362_),
    .B2(_09546_),
    .Y(_10363_));
 sky130_fd_sc_hd__nor2_2 _17625_ (.A(_10360_),
    .B(_10363_),
    .Y(_10364_));
 sky130_fd_sc_hd__nand3_4 _17626_ (.A(_10349_),
    .B(_10357_),
    .C(_10364_),
    .Y(_10365_));
 sky130_fd_sc_hd__nand2_1 _17627_ (.A(\cs_registers_i.pc_id_i[24] ),
    .B(net310),
    .Y(_10366_));
 sky130_fd_sc_hd__o21ai_0 _17628_ (.A1(net310),
    .A2(_10365_),
    .B1(_10366_),
    .Y(_10367_));
 sky130_fd_sc_hd__a22o_4 _17629_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[24] ),
    .A2(_08368_),
    .B1(_08372_),
    .B2(_10367_),
    .X(_10368_));
 sky130_fd_sc_hd__nand2_1 _17630_ (.A(net739),
    .B(_10368_),
    .Y(_10369_));
 sky130_fd_sc_hd__o31ai_4 _17631_ (.A1(_10343_),
    .A2(_08290_),
    .A3(_08503_),
    .B1(_10369_),
    .Y(_10370_));
 sky130_fd_sc_hd__mux2i_2 _17632_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[184] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[248] ),
    .S(net364),
    .Y(_10371_));
 sky130_fd_sc_hd__mux2i_2 _17633_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[152] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[216] ),
    .S(net364),
    .Y(_10372_));
 sky130_fd_sc_hd__mux2_1 _17634_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[56] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[120] ),
    .S(net364),
    .X(_10373_));
 sky130_fd_sc_hd__a221oi_2 _17635_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[88] ),
    .A2(net324),
    .B1(_10373_),
    .B2(net1476),
    .C1(net343),
    .Y(_10374_));
 sky130_fd_sc_hd__a221oi_4 _17636_ (.A1(_08152_),
    .A2(_10371_),
    .B1(_10372_),
    .B2(net592),
    .C1(_10374_),
    .Y(_10375_));
 sky130_fd_sc_hd__mux4_1 _17637_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[536] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[600] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[664] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[728] ),
    .S0(net354),
    .S1(net342),
    .X(_10376_));
 sky130_fd_sc_hd__nand2_1 _17638_ (.A(_08658_),
    .B(_10376_),
    .Y(_10377_));
 sky130_fd_sc_hd__mux4_1 _17639_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[568] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[632] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[696] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[760] ),
    .S0(net354),
    .S1(net342),
    .X(_10378_));
 sky130_fd_sc_hd__nand2_1 _17640_ (.A(net1220),
    .B(_10378_),
    .Y(_10379_));
 sky130_fd_sc_hd__nand3_2 _17641_ (.A(net698),
    .B(_10377_),
    .C(_10379_),
    .Y(_10380_));
 sky130_fd_sc_hd__nand2b_1 _17642_ (.A_N(net333),
    .B(net335),
    .Y(_10381_));
 sky130_fd_sc_hd__mux4_1 _17643_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[280] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[312] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[344] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[376] ),
    .S0(net378),
    .S1(net356),
    .X(_10382_));
 sky130_fd_sc_hd__nor3_1 _17644_ (.A(net342),
    .B(_10381_),
    .C(_10382_),
    .Y(_10383_));
 sky130_fd_sc_hd__mux4_1 _17645_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[408] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[440] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[472] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[504] ),
    .S0(net1310),
    .S1(net356),
    .X(_10384_));
 sky130_fd_sc_hd__nor3_1 _17646_ (.A(_08481_),
    .B(_10381_),
    .C(_10384_),
    .Y(_10385_));
 sky130_fd_sc_hd__mux4_1 _17647_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[792] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[856] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[920] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[984] ),
    .S0(net356),
    .S1(net342),
    .X(_10386_));
 sky130_fd_sc_hd__nand3b_1 _17648_ (.A_N(net1310),
    .B(net335),
    .C(net333),
    .Y(_10387_));
 sky130_fd_sc_hd__nand3_1 _17649_ (.A(net333),
    .B(net335),
    .C(net1309),
    .Y(_10388_));
 sky130_fd_sc_hd__mux4_1 _17650_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[824] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[888] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[952] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1016] ),
    .S0(net355),
    .S1(net342),
    .X(_10389_));
 sky130_fd_sc_hd__o22ai_2 _17651_ (.A1(_10386_),
    .A2(_10387_),
    .B1(_10388_),
    .B2(_10389_),
    .Y(_10390_));
 sky130_fd_sc_hd__nor3_2 _17652_ (.A(_10383_),
    .B(_10385_),
    .C(_10390_),
    .Y(_10391_));
 sky130_fd_sc_hd__o211ai_4 _17653_ (.A1(_10375_),
    .A2(_08163_),
    .B1(_10380_),
    .C1(_10391_),
    .Y(_10392_));
 sky130_fd_sc_hd__o22ai_1 _17654_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[56] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[24] ),
    .B2(_08503_),
    .Y(_10393_));
 sky130_fd_sc_hd__a221oi_2 _17655_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(_10365_),
    .B1(net1212),
    .B2(_08696_),
    .C1(_10393_),
    .Y(_10394_));
 sky130_fd_sc_hd__a221oi_1 _17656_ (.A1(net828),
    .A2(_08449_),
    .B1(_09455_),
    .B2(net756),
    .C1(_08495_),
    .Y(_10395_));
 sky130_fd_sc_hd__a21oi_2 _17657_ (.A1(_08495_),
    .A2(net1212),
    .B1(_10395_),
    .Y(_10396_));
 sky130_fd_sc_hd__xnor2_1 _17658_ (.A(net297),
    .B(_10396_),
    .Y(_10397_));
 sky130_fd_sc_hd__nand2_1 _17659_ (.A(net739),
    .B(_10397_),
    .Y(_10398_));
 sky130_fd_sc_hd__o21ai_2 _17660_ (.A1(_08290_),
    .A2(_10394_),
    .B1(_10398_),
    .Y(_10399_));
 sky130_fd_sc_hd__nor2_1 _17661_ (.A(_10370_),
    .B(_10399_),
    .Y(_10400_));
 sky130_fd_sc_hd__and2_1 _17662_ (.A(_10269_),
    .B(_10274_),
    .X(_10401_));
 sky130_fd_sc_hd__nor2_8 _17663_ (.A(_10401_),
    .B(net656),
    .Y(_10402_));
 sky130_fd_sc_hd__nor2_1 _17664_ (.A(_10269_),
    .B(_10274_),
    .Y(_10403_));
 sky130_fd_sc_hd__nor2_4 _17665_ (.A(_10402_),
    .B(_10403_),
    .Y(_10404_));
 sky130_fd_sc_hd__nand2_1 _17666_ (.A(_10370_),
    .B(_10399_),
    .Y(_10405_));
 sky130_fd_sc_hd__o21ai_4 _17667_ (.A1(_10400_),
    .A2(_10404_),
    .B1(_10405_),
    .Y(_10406_));
 sky130_fd_sc_hd__xnor2_4 _17668_ (.A(_10342_),
    .B(_10406_),
    .Y(_10407_));
 sky130_fd_sc_hd__inv_2 _17669_ (.A(_10407_),
    .Y(net166));
 sky130_fd_sc_hd__inv_1 _17670_ (.A(_10403_),
    .Y(_10408_));
 sky130_fd_sc_hd__a21oi_4 _17671_ (.A1(net656),
    .A2(_10408_),
    .B1(_10401_),
    .Y(_10409_));
 sky130_fd_sc_hd__xnor2_2 _17672_ (.A(_10370_),
    .B(_10399_),
    .Y(_10410_));
 sky130_fd_sc_hd__xnor2_4 _17673_ (.A(_10409_),
    .B(_10410_),
    .Y(net165));
 sky130_fd_sc_hd__inv_1 _17674_ (.A(_10410_),
    .Y(_10411_));
 sky130_fd_sc_hd__mux2_1 _17675_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[58] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[122] ),
    .S(net366),
    .X(_10412_));
 sky130_fd_sc_hd__a221oi_1 _17676_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[90] ),
    .A2(net324),
    .B1(_10412_),
    .B2(net380),
    .C1(net342),
    .Y(_10413_));
 sky130_fd_sc_hd__mux4_1 _17677_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[154] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[186] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[218] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[250] ),
    .S0(net1029),
    .S1(net1120),
    .X(_10414_));
 sky130_fd_sc_hd__o21ai_0 _17678_ (.A1(_08481_),
    .A2(_10414_),
    .B1(_08731_),
    .Y(_10415_));
 sky130_fd_sc_hd__or2_2 _17679_ (.A(_10413_),
    .B(_10415_),
    .X(_10416_));
 sky130_fd_sc_hd__mux2i_1 _17680_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[570] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[634] ),
    .S(net348),
    .Y(_10417_));
 sky130_fd_sc_hd__mux2i_1 _17681_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[538] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[602] ),
    .S(net348),
    .Y(_10418_));
 sky130_fd_sc_hd__a22oi_2 _17682_ (.A1(net1201),
    .A2(_10417_),
    .B1(_10418_),
    .B2(net650),
    .Y(_10419_));
 sky130_fd_sc_hd__mux2i_1 _17683_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[698] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[762] ),
    .S(net348),
    .Y(_10420_));
 sky130_fd_sc_hd__mux2i_1 _17684_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[666] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[730] ),
    .S(net348),
    .Y(_10421_));
 sky130_fd_sc_hd__a22oi_2 _17685_ (.A1(net1153),
    .A2(_10420_),
    .B1(_10421_),
    .B2(net1013),
    .Y(_10422_));
 sky130_fd_sc_hd__nand3_4 _17686_ (.A(net698),
    .B(_10419_),
    .C(_10422_),
    .Y(_10423_));
 sky130_fd_sc_hd__mux2i_1 _17687_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[410] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[474] ),
    .S(net348),
    .Y(_10424_));
 sky130_fd_sc_hd__mux2i_1 _17688_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[442] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[506] ),
    .S(net348),
    .Y(_10425_));
 sky130_fd_sc_hd__o22ai_2 _17689_ (.A1(net892),
    .A2(_10424_),
    .B1(_10425_),
    .B2(net871),
    .Y(_10426_));
 sky130_fd_sc_hd__mux2i_1 _17690_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[282] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[346] ),
    .S(net348),
    .Y(_10427_));
 sky130_fd_sc_hd__mux2i_1 _17691_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[314] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[378] ),
    .S(net348),
    .Y(_10428_));
 sky130_fd_sc_hd__o22ai_2 _17692_ (.A1(net772),
    .A2(_10427_),
    .B1(_10428_),
    .B2(net760),
    .Y(_10429_));
 sky130_fd_sc_hd__mux2i_1 _17693_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[794] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[858] ),
    .S(net348),
    .Y(_10430_));
 sky130_fd_sc_hd__mux2i_1 _17694_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[826] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[890] ),
    .S(net348),
    .Y(_10431_));
 sky130_fd_sc_hd__o22ai_2 _17695_ (.A1(net508),
    .A2(_10430_),
    .B1(_10431_),
    .B2(net519),
    .Y(_10432_));
 sky130_fd_sc_hd__mux2i_1 _17696_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[922] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[986] ),
    .S(net348),
    .Y(_10433_));
 sky130_fd_sc_hd__mux2i_1 _17697_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[954] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1018] ),
    .S(net348),
    .Y(_10434_));
 sky130_fd_sc_hd__o22ai_2 _17698_ (.A1(net602),
    .A2(_10433_),
    .B1(_10434_),
    .B2(net629),
    .Y(_10435_));
 sky130_fd_sc_hd__nor4_4 _17699_ (.A(_10426_),
    .B(_10429_),
    .C(_10435_),
    .D(_10432_),
    .Y(_10436_));
 sky130_fd_sc_hd__nand3_4 _17700_ (.A(_10416_),
    .B(_10423_),
    .C(net884),
    .Y(_10437_));
 sky130_fd_sc_hd__nand2_1 _17701_ (.A(net667),
    .B(_09455_),
    .Y(_10438_));
 sky130_fd_sc_hd__a21oi_1 _17702_ (.A1(_10041_),
    .A2(_10438_),
    .B1(_08495_),
    .Y(_10439_));
 sky130_fd_sc_hd__a21oi_2 _17703_ (.A1(_08495_),
    .A2(_10437_),
    .B1(_10439_),
    .Y(_10440_));
 sky130_fd_sc_hd__xnor2_1 _17704_ (.A(net297),
    .B(_10440_),
    .Y(_10441_));
 sky130_fd_sc_hd__mux4_1 _17705_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[666] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[698] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[730] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[762] ),
    .S0(net1135),
    .S1(net1233),
    .X(_10442_));
 sky130_fd_sc_hd__mux4_1 _17706_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[538] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[570] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[602] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[634] ),
    .S0(net1135),
    .S1(net1233),
    .X(_10443_));
 sky130_fd_sc_hd__a22oi_4 _17707_ (.A1(net611),
    .A2(_10442_),
    .B1(_10443_),
    .B2(_08342_),
    .Y(_10444_));
 sky130_fd_sc_hd__mux4_1 _17708_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[922] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[954] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[986] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1018] ),
    .S0(net1135),
    .S1(net1233),
    .X(_10445_));
 sky130_fd_sc_hd__mux4_1 _17709_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[794] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[826] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[858] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[890] ),
    .S0(net1135),
    .S1(net1233),
    .X(_10446_));
 sky130_fd_sc_hd__a22oi_4 _17710_ (.A1(net1248),
    .A2(_10445_),
    .B1(_10446_),
    .B2(net532),
    .Y(_10447_));
 sky130_fd_sc_hd__nand3_2 _17711_ (.A(net386),
    .B(_10444_),
    .C(_10447_),
    .Y(_10448_));
 sky130_fd_sc_hd__mux4_2 _17712_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[154] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[186] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[218] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[250] ),
    .S0(net853),
    .S1(net794),
    .X(_10449_));
 sky130_fd_sc_hd__nor2_2 _17713_ (.A(_08529_),
    .B(_10449_),
    .Y(_10450_));
 sky130_fd_sc_hd__mux2_1 _17714_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[90] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[122] ),
    .S(net1084),
    .X(_10451_));
 sky130_fd_sc_hd__a221oi_4 _17715_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[58] ),
    .A2(net539),
    .B1(_10451_),
    .B2(net413),
    .C1(net400),
    .Y(_10452_));
 sky130_fd_sc_hd__mux4_1 _17716_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[410] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[442] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[474] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[506] ),
    .S0(net1135),
    .S1(net1233),
    .X(_10453_));
 sky130_fd_sc_hd__mux4_1 _17717_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[282] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[314] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[346] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[378] ),
    .S0(net1135),
    .S1(net1233),
    .X(_10454_));
 sky130_fd_sc_hd__a22oi_4 _17718_ (.A1(net1248),
    .A2(_10453_),
    .B1(_10454_),
    .B2(net532),
    .Y(_10455_));
 sky130_fd_sc_hd__o311ai_4 _17719_ (.A1(net1075),
    .A2(_10450_),
    .A3(_10452_),
    .B1(_10455_),
    .C1(_08512_),
    .Y(_10456_));
 sky130_fd_sc_hd__nand2_8 _17720_ (.A(_10448_),
    .B(_10456_),
    .Y(_10457_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_858 ();
 sky130_fd_sc_hd__o22ai_1 _17723_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[58] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[26] ),
    .B2(_08503_),
    .Y(_10460_));
 sky130_fd_sc_hd__nor2_1 _17724_ (.A(_08504_),
    .B(_10437_),
    .Y(_10461_));
 sky130_fd_sc_hd__a2111oi_0 _17725_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(_10457_),
    .B1(_10460_),
    .C1(_10461_),
    .D1(net739),
    .Y(_10462_));
 sky130_fd_sc_hd__a21o_2 _17726_ (.A1(net739),
    .A2(_10441_),
    .B1(_10462_),
    .X(_10463_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_857 ();
 sky130_fd_sc_hd__nor2_1 _17728_ (.A(net310),
    .B(_10457_),
    .Y(_10465_));
 sky130_fd_sc_hd__a21oi_1 _17729_ (.A1(\cs_registers_i.pc_id_i[26] ),
    .A2(net310),
    .B1(_10465_),
    .Y(_10466_));
 sky130_fd_sc_hd__nand2_1 _17730_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[26] ),
    .B(_08368_),
    .Y(_10467_));
 sky130_fd_sc_hd__o21ai_4 _17731_ (.A1(net933),
    .A2(_10466_),
    .B1(_10467_),
    .Y(_10468_));
 sky130_fd_sc_hd__and3_1 _17732_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[58] ),
    .B(_08272_),
    .C(_08377_),
    .X(_10469_));
 sky130_fd_sc_hd__a21oi_2 _17733_ (.A1(_08290_),
    .A2(_10468_),
    .B1(_10469_),
    .Y(_10470_));
 sky130_fd_sc_hd__xor2_4 _17734_ (.A(_10463_),
    .B(_10470_),
    .X(_10471_));
 sky130_fd_sc_hd__nand4_4 _17735_ (.A(_10275_),
    .B(_10342_),
    .C(_10411_),
    .D(_10471_),
    .Y(_10472_));
 sky130_fd_sc_hd__nand2_1 _17736_ (.A(_10463_),
    .B(_10470_),
    .Y(_10473_));
 sky130_fd_sc_hd__maj3_1 _17737_ (.A(_10370_),
    .B(_10399_),
    .C(_10403_),
    .X(_10474_));
 sky130_fd_sc_hd__maj3_1 _17738_ (.A(_10306_),
    .B(_10340_),
    .C(_10474_),
    .X(_10475_));
 sky130_fd_sc_hd__nor2_1 _17739_ (.A(_10463_),
    .B(_10470_),
    .Y(_10476_));
 sky130_fd_sc_hd__a21oi_4 _17740_ (.A1(_10475_),
    .A2(_10473_),
    .B1(_10476_),
    .Y(_10477_));
 sky130_fd_sc_hd__o21ai_4 _17741_ (.A1(_10472_),
    .A2(_10216_),
    .B1(_10477_),
    .Y(_10478_));
 sky130_fd_sc_hd__mux4_2 _17742_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[923] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[955] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[987] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1019] ),
    .S0(net856),
    .S1(net405),
    .X(_10479_));
 sky130_fd_sc_hd__mux4_1 _17743_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[795] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[827] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[859] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[891] ),
    .S0(net856),
    .S1(net405),
    .X(_10480_));
 sky130_fd_sc_hd__mux4_1 _17744_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[667] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[699] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[731] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[763] ),
    .S0(net1284),
    .S1(net405),
    .X(_10481_));
 sky130_fd_sc_hd__mux4_1 _17745_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[539] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[571] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[603] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[635] ),
    .S0(net1076),
    .S1(net405),
    .X(_10482_));
 sky130_fd_sc_hd__a22o_4 _17746_ (.A1(net610),
    .A2(_10481_),
    .B1(_10482_),
    .B2(_08342_),
    .X(_10483_));
 sky130_fd_sc_hd__a221oi_4 _17747_ (.A1(net1248),
    .A2(_10479_),
    .B1(_10480_),
    .B2(net534),
    .C1(_10483_),
    .Y(_10484_));
 sky130_fd_sc_hd__mux4_2 _17748_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[155] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[187] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[219] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[251] ),
    .S0(net854),
    .S1(net794),
    .X(_10485_));
 sky130_fd_sc_hd__nor2_1 _17749_ (.A(_08529_),
    .B(_10485_),
    .Y(_10486_));
 sky130_fd_sc_hd__mux2_1 _17750_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[91] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[123] ),
    .S(net1084),
    .X(_10487_));
 sky130_fd_sc_hd__a221oi_1 _17751_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[59] ),
    .A2(net539),
    .B1(_10487_),
    .B2(net413),
    .C1(net400),
    .Y(_10488_));
 sky130_fd_sc_hd__mux4_2 _17752_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[411] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[443] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[475] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[507] ),
    .S0(net1284),
    .S1(net405),
    .X(_10489_));
 sky130_fd_sc_hd__mux4_1 _17753_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[283] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[315] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[347] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[379] ),
    .S0(net1284),
    .S1(net405),
    .X(_10490_));
 sky130_fd_sc_hd__a22oi_4 _17754_ (.A1(net565),
    .A2(_10489_),
    .B1(_10490_),
    .B2(net533),
    .Y(_10491_));
 sky130_fd_sc_hd__o31a_1 _17755_ (.A1(net390),
    .A2(_10486_),
    .A3(_10488_),
    .B1(_10491_),
    .X(_10492_));
 sky130_fd_sc_hd__mux2_8 _17756_ (.A0(_10484_),
    .A1(_10492_),
    .S(_08512_),
    .X(_10493_));
 sky130_fd_sc_hd__nor2_1 _17757_ (.A(net310),
    .B(_10493_),
    .Y(_10494_));
 sky130_fd_sc_hd__a21oi_1 _17758_ (.A1(\cs_registers_i.pc_id_i[27] ),
    .A2(net310),
    .B1(_10494_),
    .Y(_10495_));
 sky130_fd_sc_hd__nand2_1 _17759_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[27] ),
    .B(_08368_),
    .Y(_10496_));
 sky130_fd_sc_hd__o21ai_4 _17760_ (.A1(net933),
    .A2(_10495_),
    .B1(_10496_),
    .Y(_10497_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_856 ();
 sky130_fd_sc_hd__and3_1 _17762_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[59] ),
    .B(_08272_),
    .C(_08377_),
    .X(_10499_));
 sky130_fd_sc_hd__a21oi_2 _17763_ (.A1(_08290_),
    .A2(_10497_),
    .B1(_10499_),
    .Y(_10500_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_855 ();
 sky130_fd_sc_hd__nand2_1 _17765_ (.A(net805),
    .B(_09455_),
    .Y(_10502_));
 sky130_fd_sc_hd__mux2i_1 _17766_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[667] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[731] ),
    .S(net347),
    .Y(_10503_));
 sky130_fd_sc_hd__mux2i_1 _17767_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[571] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[635] ),
    .S(net347),
    .Y(_10504_));
 sky130_fd_sc_hd__a22oi_1 _17768_ (.A1(net1474),
    .A2(_10503_),
    .B1(_10504_),
    .B2(net329),
    .Y(_10505_));
 sky130_fd_sc_hd__mux2i_1 _17769_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[539] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[603] ),
    .S(net347),
    .Y(_10506_));
 sky130_fd_sc_hd__mux2i_1 _17770_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[699] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[763] ),
    .S(net347),
    .Y(_10507_));
 sky130_fd_sc_hd__a22oi_1 _17771_ (.A1(net1043),
    .A2(_10506_),
    .B1(_10507_),
    .B2(_08152_),
    .Y(_10508_));
 sky130_fd_sc_hd__and3_2 _17772_ (.A(net698),
    .B(_10505_),
    .C(_10508_),
    .X(_10509_));
 sky130_fd_sc_hd__mux2_1 _17773_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[59] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[123] ),
    .S(net366),
    .X(_10510_));
 sky130_fd_sc_hd__a221oi_2 _17774_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[91] ),
    .A2(net324),
    .B1(_10510_),
    .B2(net1476),
    .C1(net342),
    .Y(_10511_));
 sky130_fd_sc_hd__mux4_1 _17775_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[155] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[187] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[219] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[251] ),
    .S0(net381),
    .S1(net514),
    .X(_10512_));
 sky130_fd_sc_hd__o21ai_2 _17776_ (.A1(_08481_),
    .A2(_10512_),
    .B1(_08731_),
    .Y(_10513_));
 sky130_fd_sc_hd__nor2_4 _17777_ (.A(_10511_),
    .B(_10513_),
    .Y(_10514_));
 sky130_fd_sc_hd__mux4_1 _17778_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[411] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[443] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[475] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[507] ),
    .S0(net1309),
    .S1(net348),
    .X(_10515_));
 sky130_fd_sc_hd__mux4_1 _17779_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[923] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[955] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[987] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1019] ),
    .S0(net1309),
    .S1(net348),
    .X(_10516_));
 sky130_fd_sc_hd__a32oi_1 _17780_ (.A1(net338),
    .A2(net700),
    .A3(_10515_),
    .B1(_10516_),
    .B2(_08688_),
    .Y(_10517_));
 sky130_fd_sc_hd__mux4_1 _17781_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[283] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[315] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[347] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[379] ),
    .S0(net1309),
    .S1(net348),
    .X(_10518_));
 sky130_fd_sc_hd__mux4_1 _17782_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[795] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[827] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[859] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[891] ),
    .S0(net1309),
    .S1(net347),
    .X(_10519_));
 sky130_fd_sc_hd__a32oi_1 _17783_ (.A1(_08481_),
    .A2(net700),
    .A3(_10518_),
    .B1(_10519_),
    .B2(_08687_),
    .Y(_10520_));
 sky130_fd_sc_hd__nand2_1 _17784_ (.A(_10517_),
    .B(_10520_),
    .Y(_10521_));
 sky130_fd_sc_hd__or3_4 _17785_ (.A(_10509_),
    .B(_10514_),
    .C(_10521_),
    .X(_10522_));
 sky130_fd_sc_hd__nor2_1 _17786_ (.A(_08436_),
    .B(_10522_),
    .Y(_10523_));
 sky130_fd_sc_hd__a31oi_2 _17787_ (.A1(_08436_),
    .A2(_10041_),
    .A3(_10502_),
    .B1(_10523_),
    .Y(_10524_));
 sky130_fd_sc_hd__xnor2_1 _17788_ (.A(net296),
    .B(_10524_),
    .Y(_10525_));
 sky130_fd_sc_hd__o22ai_1 _17789_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[59] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[27] ),
    .B2(_08503_),
    .Y(_10526_));
 sky130_fd_sc_hd__a21oi_1 _17790_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(_10493_),
    .B1(_10526_),
    .Y(_10527_));
 sky130_fd_sc_hd__o211ai_1 _17791_ (.A1(_08504_),
    .A2(_10522_),
    .B1(_10527_),
    .C1(net314),
    .Y(_10528_));
 sky130_fd_sc_hd__o21ai_2 _17792_ (.A1(net314),
    .A2(_10525_),
    .B1(_10528_),
    .Y(_10529_));
 sky130_fd_sc_hd__xnor2_2 _17793_ (.A(_10500_),
    .B(_10529_),
    .Y(_10530_));
 sky130_fd_sc_hd__xnor2_4 _17794_ (.A(_10530_),
    .B(net1071),
    .Y(net168));
 sky130_fd_sc_hd__nand2_1 _17795_ (.A(_10306_),
    .B(_10340_),
    .Y(_10531_));
 sky130_fd_sc_hd__nand2_1 _17796_ (.A(_10405_),
    .B(_10531_),
    .Y(_10532_));
 sky130_fd_sc_hd__nand2_1 _17797_ (.A(_10400_),
    .B(_10531_),
    .Y(_10533_));
 sky130_fd_sc_hd__o221ai_4 _17798_ (.A1(_10306_),
    .A2(_10340_),
    .B1(_10532_),
    .B2(_10409_),
    .C1(_10533_),
    .Y(_10534_));
 sky130_fd_sc_hd__xor2_4 _17799_ (.A(_10471_),
    .B(_10534_),
    .X(_10535_));
 sky130_fd_sc_hd__inv_8 _17800_ (.A(net1041),
    .Y(net167));
 sky130_fd_sc_hd__mux2_1 _17801_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[221] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[253] ),
    .S(net1129),
    .X(_10536_));
 sky130_fd_sc_hd__mux2_1 _17802_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[93] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[125] ),
    .S(net434),
    .X(_10537_));
 sky130_fd_sc_hd__o22ai_2 _17803_ (.A1(_08815_),
    .A2(_10536_),
    .B1(_10537_),
    .B2(_08819_),
    .Y(_10538_));
 sky130_fd_sc_hd__mux2_1 _17804_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[157] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[189] ),
    .S(net1129),
    .X(_10539_));
 sky130_fd_sc_hd__a221oi_2 _17805_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[61] ),
    .A2(_09530_),
    .B1(_10539_),
    .B2(net398),
    .C1(net401),
    .Y(_10540_));
 sky130_fd_sc_hd__o21ai_4 _17806_ (.A1(_10538_),
    .A2(_10540_),
    .B1(_08179_),
    .Y(_10541_));
 sky130_fd_sc_hd__mux2_1 _17807_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[541] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[573] ),
    .S(net436),
    .X(_10542_));
 sky130_fd_sc_hd__nand2b_1 _17808_ (.A_N(\gen_regfile_ff.register_file_i.rf_reg[637] ),
    .B(net436),
    .Y(_10543_));
 sky130_fd_sc_hd__o221ai_4 _17809_ (.A1(net436),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[605] ),
    .B1(_10542_),
    .B2(net401),
    .C1(_10543_),
    .Y(_10544_));
 sky130_fd_sc_hd__mux2_1 _17810_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[669] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[701] ),
    .S(net436),
    .X(_10545_));
 sky130_fd_sc_hd__mux2_1 _17811_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[733] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[765] ),
    .S(net436),
    .X(_10546_));
 sky130_fd_sc_hd__o211ai_2 _17812_ (.A1(net401),
    .A2(_10545_),
    .B1(_10546_),
    .C1(net396),
    .Y(_10547_));
 sky130_fd_sc_hd__a221oi_2 _17813_ (.A1(net1149),
    .A2(_10545_),
    .B1(_10542_),
    .B2(net649),
    .C1(_09032_),
    .Y(_10548_));
 sky130_fd_sc_hd__o211ai_4 _17814_ (.A1(net396),
    .A2(_10544_),
    .B1(_10547_),
    .C1(_10548_),
    .Y(_10549_));
 sky130_fd_sc_hd__mux4_1 _17815_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[925] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[957] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[989] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1021] ),
    .S0(net962),
    .S1(net406),
    .X(_10550_));
 sky130_fd_sc_hd__mux4_1 _17816_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[797] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[829] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[861] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[893] ),
    .S0(net962),
    .S1(net406),
    .X(_10551_));
 sky130_fd_sc_hd__o22ai_1 _17817_ (.A1(_09265_),
    .A2(_10550_),
    .B1(_10551_),
    .B2(_09264_),
    .Y(_10552_));
 sky130_fd_sc_hd__mux4_1 _17818_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[349] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[381] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[477] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[509] ),
    .S0(net962),
    .S1(net395),
    .X(_10553_));
 sky130_fd_sc_hd__mux4_1 _17819_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[285] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[317] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[413] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[445] ),
    .S0(net962),
    .S1(net395),
    .X(_10554_));
 sky130_fd_sc_hd__o22ai_2 _17820_ (.A1(_09543_),
    .A2(_10553_),
    .B1(_10554_),
    .B2(_09546_),
    .Y(_10555_));
 sky130_fd_sc_hd__nor2_2 _17821_ (.A(_10552_),
    .B(_10555_),
    .Y(_10556_));
 sky130_fd_sc_hd__nand3_4 _17822_ (.A(_10541_),
    .B(_10549_),
    .C(_10556_),
    .Y(_10557_));
 sky130_fd_sc_hd__nor2_1 _17823_ (.A(net310),
    .B(_10557_),
    .Y(_10558_));
 sky130_fd_sc_hd__a21oi_1 _17824_ (.A1(\cs_registers_i.pc_id_i[29] ),
    .A2(net310),
    .B1(_10558_),
    .Y(_10559_));
 sky130_fd_sc_hd__nand2_1 _17825_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[29] ),
    .B(_08368_),
    .Y(_10560_));
 sky130_fd_sc_hd__o21ai_4 _17826_ (.A1(net933),
    .A2(_10559_),
    .B1(_10560_),
    .Y(_10561_));
 sky130_fd_sc_hd__nand2_1 _17827_ (.A(net739),
    .B(_10561_),
    .Y(_10562_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_854 ();
 sky130_fd_sc_hd__nand3_1 _17829_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[61] ),
    .B(_08272_),
    .C(_08377_),
    .Y(_10564_));
 sky130_fd_sc_hd__nand2_1 _17830_ (.A(_10562_),
    .B(_10564_),
    .Y(_10565_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_853 ();
 sky130_fd_sc_hd__nand2_1 _17832_ (.A(net675),
    .B(_09455_),
    .Y(_10567_));
 sky130_fd_sc_hd__mux2i_1 _17833_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[285] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[349] ),
    .S(net359),
    .Y(_10568_));
 sky130_fd_sc_hd__mux2i_1 _17834_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[317] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[381] ),
    .S(net359),
    .Y(_10569_));
 sky130_fd_sc_hd__a22oi_1 _17835_ (.A1(net325),
    .A2(_10568_),
    .B1(_10569_),
    .B2(net328),
    .Y(_10570_));
 sky130_fd_sc_hd__mux2i_1 _17836_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[413] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[477] ),
    .S(net359),
    .Y(_10571_));
 sky130_fd_sc_hd__mux2i_1 _17837_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[445] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[509] ),
    .S(net359),
    .Y(_10572_));
 sky130_fd_sc_hd__a22oi_1 _17838_ (.A1(net1119),
    .A2(_10571_),
    .B1(_10572_),
    .B2(net1153),
    .Y(_10573_));
 sky130_fd_sc_hd__nand3_2 _17839_ (.A(net701),
    .B(_10570_),
    .C(_10573_),
    .Y(_10574_));
 sky130_fd_sc_hd__mux2i_1 _17840_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[573] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[637] ),
    .S(net1030),
    .Y(_10575_));
 sky130_fd_sc_hd__mux2i_1 _17841_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[669] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[733] ),
    .S(net1030),
    .Y(_10576_));
 sky130_fd_sc_hd__a22oi_1 _17842_ (.A1(net328),
    .A2(_10575_),
    .B1(_10576_),
    .B2(net592),
    .Y(_10577_));
 sky130_fd_sc_hd__mux2i_1 _17843_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[541] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[605] ),
    .S(net1030),
    .Y(_10578_));
 sky130_fd_sc_hd__mux2i_1 _17844_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[701] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[765] ),
    .S(net1030),
    .Y(_10579_));
 sky130_fd_sc_hd__a22oi_1 _17845_ (.A1(net325),
    .A2(_10578_),
    .B1(_10579_),
    .B2(net1153),
    .Y(_10580_));
 sky130_fd_sc_hd__nand3_1 _17846_ (.A(net698),
    .B(_10577_),
    .C(_10580_),
    .Y(_10581_));
 sky130_fd_sc_hd__mux2_1 _17847_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[61] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[125] ),
    .S(net363),
    .X(_10582_));
 sky130_fd_sc_hd__a221oi_2 _17848_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[93] ),
    .A2(net324),
    .B1(_10582_),
    .B2(net983),
    .C1(net341),
    .Y(_10583_));
 sky130_fd_sc_hd__mux4_1 _17849_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[157] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[189] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[221] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[253] ),
    .S0(net375),
    .S1(net1077),
    .X(_10584_));
 sky130_fd_sc_hd__o21ai_2 _17850_ (.A1(_08481_),
    .A2(_10584_),
    .B1(_08731_),
    .Y(_10585_));
 sky130_fd_sc_hd__mux4_1 _17851_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[925] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[957] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[989] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1021] ),
    .S0(net373),
    .S1(net359),
    .X(_10586_));
 sky130_fd_sc_hd__mux4_1 _17852_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[797] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[829] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[861] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[893] ),
    .S0(net373),
    .S1(net359),
    .X(_10587_));
 sky130_fd_sc_hd__a22oi_1 _17853_ (.A1(_08688_),
    .A2(_10586_),
    .B1(_10587_),
    .B2(_08687_),
    .Y(_10588_));
 sky130_fd_sc_hd__o21a_1 _17854_ (.A1(_10583_),
    .A2(_10585_),
    .B1(_10588_),
    .X(_10589_));
 sky130_fd_sc_hd__nand3_4 _17855_ (.A(_10574_),
    .B(_10581_),
    .C(_10589_),
    .Y(_10590_));
 sky130_fd_sc_hd__nor2_1 _17856_ (.A(_08436_),
    .B(_10590_),
    .Y(_10591_));
 sky130_fd_sc_hd__a31oi_2 _17857_ (.A1(_08436_),
    .A2(_10041_),
    .A3(_10567_),
    .B1(_10591_),
    .Y(_10592_));
 sky130_fd_sc_hd__xor2_1 _17858_ (.A(net296),
    .B(_10592_),
    .X(_10593_));
 sky130_fd_sc_hd__o22ai_1 _17859_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[61] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[29] ),
    .B2(_08503_),
    .Y(_10594_));
 sky130_fd_sc_hd__nor2_1 _17860_ (.A(_08504_),
    .B(_10590_),
    .Y(_10595_));
 sky130_fd_sc_hd__a2111oi_1 _17861_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(_10557_),
    .B1(_10594_),
    .C1(_10595_),
    .D1(net739),
    .Y(_10596_));
 sky130_fd_sc_hd__a21oi_2 _17862_ (.A1(net739),
    .A2(_10593_),
    .B1(_10596_),
    .Y(_10597_));
 sky130_fd_sc_hd__xnor2_2 _17863_ (.A(_10565_),
    .B(_10597_),
    .Y(_10598_));
 sky130_fd_sc_hd__mux2_1 _17864_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[60] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[124] ),
    .S(net1120),
    .X(_10599_));
 sky130_fd_sc_hd__a22oi_2 _17865_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[92] ),
    .A2(net324),
    .B1(_10599_),
    .B2(net983),
    .Y(_10600_));
 sky130_fd_sc_hd__mux4_1 _17866_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[156] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[188] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[220] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[252] ),
    .S0(net983),
    .S1(net1120),
    .X(_10601_));
 sky130_fd_sc_hd__nand2_1 _17867_ (.A(net343),
    .B(_10601_),
    .Y(_10602_));
 sky130_fd_sc_hd__o211ai_4 _17868_ (.A1(net343),
    .A2(_10600_),
    .B1(_10602_),
    .C1(_08731_),
    .Y(_10603_));
 sky130_fd_sc_hd__mux4_1 _17869_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[540] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[604] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[668] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[732] ),
    .S0(net354),
    .S1(net342),
    .X(_10604_));
 sky130_fd_sc_hd__nor3_1 _17870_ (.A(net1220),
    .B(_08679_),
    .C(_10604_),
    .Y(_10605_));
 sky130_fd_sc_hd__and2_0 _17871_ (.A(\gen_regfile_ff.register_file_i.rf_reg[924] ),
    .B(\gen_regfile_ff.register_file_i.rf_reg[956] ),
    .X(_10606_));
 sky130_fd_sc_hd__and4_1 _17872_ (.A(net356),
    .B(net342),
    .C(\gen_regfile_ff.register_file_i.rf_reg[988] ),
    .D(\gen_regfile_ff.register_file_i.rf_reg[1020] ),
    .X(_10607_));
 sky130_fd_sc_hd__mux4_1 _17873_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[796] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[860] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[924] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[988] ),
    .S0(net356),
    .S1(net342),
    .X(_10608_));
 sky130_fd_sc_hd__a2111oi_1 _17874_ (.A1(_08669_),
    .A2(_10606_),
    .B1(_10607_),
    .C1(_10608_),
    .D1(_10387_),
    .Y(_10609_));
 sky130_fd_sc_hd__mux4_1 _17875_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[572] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[636] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[700] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[764] ),
    .S0(net354),
    .S1(net342),
    .X(_10610_));
 sky130_fd_sc_hd__nor3_1 _17876_ (.A(_08658_),
    .B(_08679_),
    .C(_10610_),
    .Y(_10611_));
 sky130_fd_sc_hd__mux4_1 _17877_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[284] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[316] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[348] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[380] ),
    .S0(net1220),
    .S1(net356),
    .X(_10612_));
 sky130_fd_sc_hd__nor3_1 _17878_ (.A(net342),
    .B(_10381_),
    .C(_10612_),
    .Y(_10613_));
 sky130_fd_sc_hd__nor4_2 _17879_ (.A(_10605_),
    .B(_10609_),
    .C(_10611_),
    .D(_10613_),
    .Y(_10614_));
 sky130_fd_sc_hd__mux4_1 _17880_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[828] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[892] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[956] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1020] ),
    .S0(net356),
    .S1(net342),
    .X(_10615_));
 sky130_fd_sc_hd__nor3_1 _17881_ (.A(_08161_),
    .B(_08658_),
    .C(_10615_),
    .Y(_10616_));
 sky130_fd_sc_hd__mux4_1 _17882_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[412] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[444] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[476] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[508] ),
    .S0(net1220),
    .S1(net356),
    .X(_10617_));
 sky130_fd_sc_hd__nor3_1 _17883_ (.A(net333),
    .B(_08481_),
    .C(_10617_),
    .Y(_10618_));
 sky130_fd_sc_hd__o21ai_2 _17884_ (.A1(_10616_),
    .A2(_10618_),
    .B1(net335),
    .Y(_10619_));
 sky130_fd_sc_hd__nand3_4 _17885_ (.A(_10603_),
    .B(_10614_),
    .C(_10619_),
    .Y(_10620_));
 sky130_fd_sc_hd__a221oi_4 _17886_ (.A1(net829),
    .A2(_08449_),
    .B1(_09455_),
    .B2(net815),
    .C1(_08495_),
    .Y(_10621_));
 sky130_fd_sc_hd__a21oi_2 _17887_ (.A1(_08495_),
    .A2(_10620_),
    .B1(_10621_),
    .Y(_10622_));
 sky130_fd_sc_hd__xor2_1 _17888_ (.A(net296),
    .B(_10622_),
    .X(_10623_));
 sky130_fd_sc_hd__mux2_1 _17889_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[156] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[188] ),
    .S(net753),
    .X(_10624_));
 sky130_fd_sc_hd__a22oi_2 _17890_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[60] ),
    .A2(_09530_),
    .B1(_10624_),
    .B2(net398),
    .Y(_10625_));
 sky130_fd_sc_hd__mux4_1 _17891_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[92] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[124] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[220] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[252] ),
    .S0(net753),
    .S1(net398),
    .X(_10626_));
 sky130_fd_sc_hd__nand2_1 _17892_ (.A(net403),
    .B(_10626_),
    .Y(_10627_));
 sky130_fd_sc_hd__o211ai_4 _17893_ (.A1(net403),
    .A2(_10625_),
    .B1(_10627_),
    .C1(_08179_),
    .Y(_10628_));
 sky130_fd_sc_hd__mux2_1 _17894_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[924] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[956] ),
    .S(net1080),
    .X(_10629_));
 sky130_fd_sc_hd__nand2b_1 _17895_ (.A_N(\gen_regfile_ff.register_file_i.rf_reg[1020] ),
    .B(net865),
    .Y(_10630_));
 sky130_fd_sc_hd__o221ai_2 _17896_ (.A1(net865),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[988] ),
    .B1(_10629_),
    .B2(net1009),
    .C1(_10630_),
    .Y(_10631_));
 sky130_fd_sc_hd__mux2_1 _17897_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[796] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[828] ),
    .S(net865),
    .X(_10632_));
 sky130_fd_sc_hd__mux2_1 _17898_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[860] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[892] ),
    .S(net865),
    .X(_10633_));
 sky130_fd_sc_hd__o211ai_2 _17899_ (.A1(net1009),
    .A2(_10632_),
    .B1(_10633_),
    .C1(_08529_),
    .Y(_10634_));
 sky130_fd_sc_hd__a221oi_2 _17900_ (.A1(net1149),
    .A2(_10629_),
    .B1(_10632_),
    .B2(net649),
    .C1(_08809_),
    .Y(_10635_));
 sky130_fd_sc_hd__o211ai_4 _17901_ (.A1(_08529_),
    .A2(_10631_),
    .B1(_10634_),
    .C1(_10635_),
    .Y(_10636_));
 sky130_fd_sc_hd__mux4_1 _17902_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[348] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[380] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[476] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[508] ),
    .S0(net963),
    .S1(net399),
    .X(_10637_));
 sky130_fd_sc_hd__mux4_1 _17903_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[284] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[316] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[412] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[444] ),
    .S0(net963),
    .S1(net399),
    .X(_10638_));
 sky130_fd_sc_hd__o22ai_2 _17904_ (.A1(_09543_),
    .A2(_10637_),
    .B1(_10638_),
    .B2(_09546_),
    .Y(_10639_));
 sky130_fd_sc_hd__mux4_1 _17905_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[668] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[700] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[732] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[764] ),
    .S0(net865),
    .S1(net1083),
    .X(_10640_));
 sky130_fd_sc_hd__mux4_1 _17906_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[540] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[572] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[604] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[636] ),
    .S0(net865),
    .S1(net1083),
    .X(_10641_));
 sky130_fd_sc_hd__o22ai_2 _17907_ (.A1(_09279_),
    .A2(_10640_),
    .B1(_10641_),
    .B2(_09550_),
    .Y(_10642_));
 sky130_fd_sc_hd__nor2_2 _17908_ (.A(_10639_),
    .B(_10642_),
    .Y(_10643_));
 sky130_fd_sc_hd__nand3_4 _17909_ (.A(_10628_),
    .B(_10636_),
    .C(_10643_),
    .Y(_10644_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_852 ();
 sky130_fd_sc_hd__o22ai_1 _17911_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[60] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[28] ),
    .B2(_08503_),
    .Y(_10646_));
 sky130_fd_sc_hd__a21oi_1 _17912_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(_10644_),
    .B1(_10646_),
    .Y(_10647_));
 sky130_fd_sc_hd__nor2_1 _17913_ (.A(_08504_),
    .B(_10620_),
    .Y(_10648_));
 sky130_fd_sc_hd__a21oi_1 _17914_ (.A1(_08504_),
    .A2(_10647_),
    .B1(_10648_),
    .Y(_10649_));
 sky130_fd_sc_hd__nor2_1 _17915_ (.A(net739),
    .B(_10649_),
    .Y(_10650_));
 sky130_fd_sc_hd__a21oi_2 _17916_ (.A1(net739),
    .A2(_10623_),
    .B1(_10650_),
    .Y(_10651_));
 sky130_fd_sc_hd__nor2_1 _17917_ (.A(net310),
    .B(_10644_),
    .Y(_10652_));
 sky130_fd_sc_hd__a21oi_1 _17918_ (.A1(\cs_registers_i.pc_id_i[28] ),
    .A2(net310),
    .B1(_10652_),
    .Y(_10653_));
 sky130_fd_sc_hd__nand2_1 _17919_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[28] ),
    .B(_08368_),
    .Y(_10654_));
 sky130_fd_sc_hd__o21ai_4 _17920_ (.A1(net933),
    .A2(_10653_),
    .B1(_10654_),
    .Y(_10655_));
 sky130_fd_sc_hd__nand2_1 _17921_ (.A(net739),
    .B(_10655_),
    .Y(_10656_));
 sky130_fd_sc_hd__nand3_1 _17922_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[60] ),
    .B(_08272_),
    .C(_08377_),
    .Y(_10657_));
 sky130_fd_sc_hd__nand2_1 _17923_ (.A(_10656_),
    .B(_10657_),
    .Y(_10658_));
 sky130_fd_sc_hd__xnor2_2 _17924_ (.A(_10651_),
    .B(_10658_),
    .Y(_10659_));
 sky130_fd_sc_hd__or2_0 _17925_ (.A(_10530_),
    .B(_10659_),
    .X(_10660_));
 sky130_fd_sc_hd__inv_1 _17926_ (.A(_10660_),
    .Y(_10661_));
 sky130_fd_sc_hd__nor2_1 _17927_ (.A(_10500_),
    .B(_10529_),
    .Y(_10662_));
 sky130_fd_sc_hd__maj3_1 _17928_ (.A(_10651_),
    .B(_10658_),
    .C(_10662_),
    .X(_10663_));
 sky130_fd_sc_hd__a21oi_4 _17929_ (.A1(_10478_),
    .A2(_10661_),
    .B1(_10663_),
    .Y(_10664_));
 sky130_fd_sc_hd__xnor2_4 _17930_ (.A(_10598_),
    .B(_10664_),
    .Y(_10665_));
 sky130_fd_sc_hd__inv_4 _17931_ (.A(net850),
    .Y(net170));
 sky130_fd_sc_hd__nand2_1 _17932_ (.A(_10500_),
    .B(_10529_),
    .Y(_10666_));
 sky130_fd_sc_hd__o21ai_4 _17933_ (.A1(_10662_),
    .A2(net1071),
    .B1(_10666_),
    .Y(_10667_));
 sky130_fd_sc_hd__xor2_4 _17934_ (.A(_10659_),
    .B(_10667_),
    .X(net169));
 sky130_fd_sc_hd__mux4_1 _17935_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[159] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[191] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[223] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[255] ),
    .S0(net1129),
    .S1(net402),
    .X(_10668_));
 sky130_fd_sc_hd__nand2_1 _17936_ (.A(net396),
    .B(_10668_),
    .Y(_10669_));
 sky130_fd_sc_hd__mux2i_1 _17937_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[95] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[127] ),
    .S(net1129),
    .Y(_10670_));
 sky130_fd_sc_hd__a21oi_1 _17938_ (.A1(net1129),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[63] ),
    .B1(net402),
    .Y(_10671_));
 sky130_fd_sc_hd__a211o_1 _17939_ (.A1(net402),
    .A2(_10670_),
    .B1(_10671_),
    .C1(net396),
    .X(_10672_));
 sky130_fd_sc_hd__mux4_1 _17940_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[927] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[959] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[991] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1023] ),
    .S0(net912),
    .S1(net401),
    .X(_10673_));
 sky130_fd_sc_hd__mux4_1 _17941_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[799] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[831] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[863] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[895] ),
    .S0(net912),
    .S1(net401),
    .X(_10674_));
 sky130_fd_sc_hd__o22ai_4 _17942_ (.A1(_09265_),
    .A2(_10673_),
    .B1(_10674_),
    .B2(_09264_),
    .Y(_10675_));
 sky130_fd_sc_hd__a31oi_4 _17943_ (.A1(_08179_),
    .A2(_10669_),
    .A3(_10672_),
    .B1(_10675_),
    .Y(_10676_));
 sky130_fd_sc_hd__mux2i_1 _17944_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[287] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[319] ),
    .S(net1074),
    .Y(_10677_));
 sky130_fd_sc_hd__mux2i_1 _17945_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[415] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[447] ),
    .S(net1074),
    .Y(_10678_));
 sky130_fd_sc_hd__a22oi_1 _17946_ (.A1(net649),
    .A2(_10677_),
    .B1(_10678_),
    .B2(net625),
    .Y(_10679_));
 sky130_fd_sc_hd__mux2i_1 _17947_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[479] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[511] ),
    .S(net1074),
    .Y(_10680_));
 sky130_fd_sc_hd__mux2i_1 _17948_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[351] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[383] ),
    .S(net1074),
    .Y(_10681_));
 sky130_fd_sc_hd__a22oi_1 _17949_ (.A1(_08803_),
    .A2(_10680_),
    .B1(_10681_),
    .B2(net614),
    .Y(_10682_));
 sky130_fd_sc_hd__a21o_2 _17950_ (.A1(_10679_),
    .A2(_10682_),
    .B1(_09275_),
    .X(_10683_));
 sky130_fd_sc_hd__mux2i_1 _17951_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[543] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[575] ),
    .S(net1074),
    .Y(_10684_));
 sky130_fd_sc_hd__mux2i_1 _17952_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[735] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[767] ),
    .S(net1074),
    .Y(_10685_));
 sky130_fd_sc_hd__a22oi_1 _17953_ (.A1(net649),
    .A2(_10684_),
    .B1(_10685_),
    .B2(_08803_),
    .Y(_10686_));
 sky130_fd_sc_hd__mux2i_1 _17954_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[671] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[703] ),
    .S(net1074),
    .Y(_10687_));
 sky130_fd_sc_hd__mux2i_1 _17955_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[607] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[639] ),
    .S(net1074),
    .Y(_10688_));
 sky130_fd_sc_hd__a22oi_1 _17956_ (.A1(net1149),
    .A2(_10687_),
    .B1(_10688_),
    .B2(net617),
    .Y(_10689_));
 sky130_fd_sc_hd__a21o_2 _17957_ (.A1(_10686_),
    .A2(_10689_),
    .B1(_09032_),
    .X(_10690_));
 sky130_fd_sc_hd__and3_4 _17958_ (.A(_10676_),
    .B(_10683_),
    .C(_10690_),
    .X(_10691_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_851 ();
 sky130_fd_sc_hd__mux2i_2 _17960_ (.A0(_10691_),
    .A1(\cs_registers_i.pc_id_i[31] ),
    .S(net310),
    .Y(_10693_));
 sky130_fd_sc_hd__nand2_1 _17961_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[31] ),
    .B(_08368_),
    .Y(_10694_));
 sky130_fd_sc_hd__o21ai_4 _17962_ (.A1(net933),
    .A2(_10693_),
    .B1(_10694_),
    .Y(_10695_));
 sky130_fd_sc_hd__mux2_1 _17963_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[63] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[127] ),
    .S(net1077),
    .X(_10696_));
 sky130_fd_sc_hd__a221oi_2 _17964_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[95] ),
    .A2(net324),
    .B1(_10696_),
    .B2(net1133),
    .C1(net341),
    .Y(_10697_));
 sky130_fd_sc_hd__mux4_1 _17965_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[159] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[191] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[223] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[255] ),
    .S0(net374),
    .S1(net1141),
    .X(_10698_));
 sky130_fd_sc_hd__nor2_1 _17966_ (.A(_08481_),
    .B(_10698_),
    .Y(_10699_));
 sky130_fd_sc_hd__or3_4 _17967_ (.A(_08163_),
    .B(_10697_),
    .C(_10699_),
    .X(_10700_));
 sky130_fd_sc_hd__mux2i_1 _17968_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[575] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[639] ),
    .S(net361),
    .Y(_10701_));
 sky130_fd_sc_hd__mux2i_1 _17969_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[671] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[735] ),
    .S(net361),
    .Y(_10702_));
 sky130_fd_sc_hd__a22oi_2 _17970_ (.A1(net328),
    .A2(_10701_),
    .B1(_10702_),
    .B2(net1119),
    .Y(_10703_));
 sky130_fd_sc_hd__mux2i_1 _17971_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[543] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[607] ),
    .S(net361),
    .Y(_10704_));
 sky130_fd_sc_hd__mux2i_1 _17972_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[703] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[767] ),
    .S(net361),
    .Y(_10705_));
 sky130_fd_sc_hd__a22oi_2 _17973_ (.A1(net325),
    .A2(_10704_),
    .B1(_10705_),
    .B2(net1153),
    .Y(_10706_));
 sky130_fd_sc_hd__nand3_4 _17974_ (.A(net698),
    .B(_10703_),
    .C(_10706_),
    .Y(_10707_));
 sky130_fd_sc_hd__mux2i_1 _17975_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[415] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[479] ),
    .S(net362),
    .Y(_10708_));
 sky130_fd_sc_hd__mux2i_1 _17976_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[447] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[511] ),
    .S(net362),
    .Y(_10709_));
 sky130_fd_sc_hd__o22ai_2 _17977_ (.A1(net894),
    .A2(_10708_),
    .B1(_10709_),
    .B2(net873),
    .Y(_10710_));
 sky130_fd_sc_hd__mux2i_1 _17978_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[287] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[351] ),
    .S(net1030),
    .Y(_10711_));
 sky130_fd_sc_hd__mux2i_1 _17979_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[319] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[383] ),
    .S(net1030),
    .Y(_10712_));
 sky130_fd_sc_hd__o22ai_2 _17980_ (.A1(net773),
    .A2(_10711_),
    .B1(_10712_),
    .B2(net763),
    .Y(_10713_));
 sky130_fd_sc_hd__mux2i_2 _17981_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[799] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[863] ),
    .S(net360),
    .Y(_10714_));
 sky130_fd_sc_hd__mux2i_2 _17982_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[831] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[895] ),
    .S(net360),
    .Y(_10715_));
 sky130_fd_sc_hd__o22ai_4 _17983_ (.A1(net506),
    .A2(_10714_),
    .B1(_10715_),
    .B2(net930),
    .Y(_10716_));
 sky130_fd_sc_hd__mux2i_2 _17984_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[927] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[991] ),
    .S(net1030),
    .Y(_10717_));
 sky130_fd_sc_hd__mux2i_2 _17985_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[959] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1023] ),
    .S(net1030),
    .Y(_10718_));
 sky130_fd_sc_hd__o22ai_4 _17986_ (.A1(net934),
    .A2(_10717_),
    .B1(_10718_),
    .B2(net1210),
    .Y(_10719_));
 sky130_fd_sc_hd__nor4_4 _17987_ (.A(_10710_),
    .B(_10713_),
    .C(_10716_),
    .D(_10719_),
    .Y(_10720_));
 sky130_fd_sc_hd__nand3_4 _17988_ (.A(_10700_),
    .B(_10707_),
    .C(_10720_),
    .Y(_10721_));
 sky130_fd_sc_hd__o21ai_0 _17989_ (.A1(_08640_),
    .A2(_08646_),
    .B1(net826),
    .Y(_10722_));
 sky130_fd_sc_hd__nor2_1 _17990_ (.A(_08495_),
    .B(_10722_),
    .Y(_10723_));
 sky130_fd_sc_hd__a21oi_4 _17991_ (.A1(_08495_),
    .A2(_10721_),
    .B1(_10723_),
    .Y(_10724_));
 sky130_fd_sc_hd__xor2_2 _17992_ (.A(net297),
    .B(_10724_),
    .X(_10725_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_850 ();
 sky130_fd_sc_hd__clkinv_2 _17994_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[63] ),
    .Y(_10727_));
 sky130_fd_sc_hd__inv_1 _17995_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[31] ),
    .Y(_10728_));
 sky130_fd_sc_hd__a221oi_2 _17996_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .A2(_10727_),
    .B1(_10728_),
    .B2(_08377_),
    .C1(net739),
    .Y(_10729_));
 sky130_fd_sc_hd__o221ai_4 _17997_ (.A1(_08500_),
    .A2(_10691_),
    .B1(_10721_),
    .B2(_08504_),
    .C1(_10729_),
    .Y(_10730_));
 sky130_fd_sc_hd__nand2_1 _17998_ (.A(_10725_),
    .B(_10730_),
    .Y(_10731_));
 sky130_fd_sc_hd__xor2_1 _17999_ (.A(_10695_),
    .B(_10731_),
    .X(_10732_));
 sky130_fd_sc_hd__nand2_1 _18000_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[63] ),
    .B(_08377_),
    .Y(_10733_));
 sky130_fd_sc_hd__xnor2_1 _18001_ (.A(_10730_),
    .B(_10733_),
    .Y(_10734_));
 sky130_fd_sc_hd__nand2_1 _18002_ (.A(net313),
    .B(_10734_),
    .Y(_10735_));
 sky130_fd_sc_hd__o21ai_2 _18003_ (.A1(net313),
    .A2(_10732_),
    .B1(_10735_),
    .Y(_10736_));
 sky130_fd_sc_hd__mux2_1 _18004_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[62] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[126] ),
    .S(net1077),
    .X(_10737_));
 sky130_fd_sc_hd__a221oi_1 _18005_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[94] ),
    .A2(net324),
    .B1(_10737_),
    .B2(net983),
    .C1(net341),
    .Y(_10738_));
 sky130_fd_sc_hd__mux4_1 _18006_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[158] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[190] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[222] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[254] ),
    .S0(net1154),
    .S1(net1077),
    .X(_10739_));
 sky130_fd_sc_hd__o21ai_0 _18007_ (.A1(_08481_),
    .A2(_10739_),
    .B1(_08731_),
    .Y(_10740_));
 sky130_fd_sc_hd__nor2_2 _18008_ (.A(_10738_),
    .B(_10740_),
    .Y(_10741_));
 sky130_fd_sc_hd__mux2i_1 _18009_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[830] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[894] ),
    .S(net1312),
    .Y(_10742_));
 sky130_fd_sc_hd__mux2i_1 _18010_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[286] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[350] ),
    .S(net1312),
    .Y(_10743_));
 sky130_fd_sc_hd__o22ai_1 _18011_ (.A1(net518),
    .A2(_10742_),
    .B1(_10743_),
    .B2(net772),
    .Y(_10744_));
 sky130_fd_sc_hd__mux2i_1 _18012_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[798] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[862] ),
    .S(net1312),
    .Y(_10745_));
 sky130_fd_sc_hd__mux2i_1 _18013_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[926] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[990] ),
    .S(net1312),
    .Y(_10746_));
 sky130_fd_sc_hd__o22ai_1 _18014_ (.A1(net508),
    .A2(_10745_),
    .B1(_10746_),
    .B2(net604),
    .Y(_10747_));
 sky130_fd_sc_hd__mux2i_1 _18015_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[446] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[510] ),
    .S(net349),
    .Y(_10748_));
 sky130_fd_sc_hd__mux2i_1 _18016_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[958] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1022] ),
    .S(net1312),
    .Y(_10749_));
 sky130_fd_sc_hd__o22ai_1 _18017_ (.A1(net870),
    .A2(_10748_),
    .B1(_10749_),
    .B2(net631),
    .Y(_10750_));
 sky130_fd_sc_hd__mux2i_1 _18018_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[414] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[478] ),
    .S(net349),
    .Y(_10751_));
 sky130_fd_sc_hd__mux2i_1 _18019_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[318] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[382] ),
    .S(net1312),
    .Y(_10752_));
 sky130_fd_sc_hd__o22ai_1 _18020_ (.A1(net892),
    .A2(_10751_),
    .B1(_10752_),
    .B2(net762),
    .Y(_10753_));
 sky130_fd_sc_hd__or4_4 _18021_ (.A(_10744_),
    .B(_10747_),
    .C(_10750_),
    .D(_10753_),
    .X(_10754_));
 sky130_fd_sc_hd__mux2i_1 _18022_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[670] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[734] ),
    .S(net988),
    .Y(_10755_));
 sky130_fd_sc_hd__mux2i_1 _18023_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[542] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[606] ),
    .S(net988),
    .Y(_10756_));
 sky130_fd_sc_hd__a22oi_1 _18024_ (.A1(net593),
    .A2(_10755_),
    .B1(_10756_),
    .B2(net325),
    .Y(_10757_));
 sky130_fd_sc_hd__mux2i_1 _18025_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[574] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[638] ),
    .S(net988),
    .Y(_10758_));
 sky130_fd_sc_hd__mux2i_1 _18026_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[702] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[766] ),
    .S(net988),
    .Y(_10759_));
 sky130_fd_sc_hd__a22oi_1 _18027_ (.A1(net328),
    .A2(_10758_),
    .B1(_10759_),
    .B2(net1153),
    .Y(_10760_));
 sky130_fd_sc_hd__and3_1 _18028_ (.A(net698),
    .B(_10757_),
    .C(_10760_),
    .X(_10761_));
 sky130_fd_sc_hd__nor3_4 _18029_ (.A(_10741_),
    .B(_10761_),
    .C(_10754_),
    .Y(_10762_));
 sky130_fd_sc_hd__a221oi_2 _18030_ (.A1(net830),
    .A2(_08449_),
    .B1(_09455_),
    .B2(net921),
    .C1(_08495_),
    .Y(_10763_));
 sky130_fd_sc_hd__a21oi_2 _18031_ (.A1(_08495_),
    .A2(net1164),
    .B1(_10763_),
    .Y(_10764_));
 sky130_fd_sc_hd__xnor2_1 _18032_ (.A(net296),
    .B(_10764_),
    .Y(_10765_));
 sky130_fd_sc_hd__mux2_1 _18033_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[734] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[766] ),
    .S(net1111),
    .X(_10766_));
 sky130_fd_sc_hd__mux2_1 _18034_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[670] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[702] ),
    .S(net1111),
    .X(_10767_));
 sky130_fd_sc_hd__o22ai_1 _18035_ (.A1(_08815_),
    .A2(_10766_),
    .B1(_10767_),
    .B2(_08811_),
    .Y(_10768_));
 sky130_fd_sc_hd__mux2i_1 _18036_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[606] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[638] ),
    .S(net1123),
    .Y(_10769_));
 sky130_fd_sc_hd__mux2i_1 _18037_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[542] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[574] ),
    .S(net962),
    .Y(_10770_));
 sky130_fd_sc_hd__a22oi_1 _18038_ (.A1(net613),
    .A2(_10769_),
    .B1(_10770_),
    .B2(net649),
    .Y(_10771_));
 sky130_fd_sc_hd__nand2b_1 _18039_ (.A_N(_10768_),
    .B(_10771_),
    .Y(_10772_));
 sky130_fd_sc_hd__mux4_1 _18040_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[926] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[958] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[990] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[1022] ),
    .S0(net1012),
    .S1(net1083),
    .X(_10773_));
 sky130_fd_sc_hd__mux4_1 _18041_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[798] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[830] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[862] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[894] ),
    .S0(net1012),
    .S1(net1078),
    .X(_10774_));
 sky130_fd_sc_hd__mux2_2 _18042_ (.A0(_10773_),
    .A1(_10774_),
    .S(_08529_),
    .X(_10775_));
 sky130_fd_sc_hd__nand2_1 _18043_ (.A(net1140),
    .B(_10775_),
    .Y(_10776_));
 sky130_fd_sc_hd__o21ai_1 _18044_ (.A1(net1140),
    .A2(_10772_),
    .B1(_10776_),
    .Y(_10777_));
 sky130_fd_sc_hd__mux2_1 _18045_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[222] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[254] ),
    .S(net436),
    .X(_10778_));
 sky130_fd_sc_hd__mux2_1 _18046_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[158] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[190] ),
    .S(net436),
    .X(_10779_));
 sky130_fd_sc_hd__o22ai_2 _18047_ (.A1(_08815_),
    .A2(_10778_),
    .B1(_10779_),
    .B2(_08811_),
    .Y(_10780_));
 sky130_fd_sc_hd__mux2_1 _18048_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[94] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[126] ),
    .S(net436),
    .X(_10781_));
 sky130_fd_sc_hd__a221oi_2 _18049_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[62] ),
    .A2(net541),
    .B1(_10781_),
    .B2(net403),
    .C1(net397),
    .Y(_10782_));
 sky130_fd_sc_hd__o21ai_0 _18050_ (.A1(_10780_),
    .A2(_10782_),
    .B1(_08309_),
    .Y(_10783_));
 sky130_fd_sc_hd__mux4_1 _18051_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[414] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[446] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[478] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[510] ),
    .S0(net423),
    .S1(net1204),
    .X(_10784_));
 sky130_fd_sc_hd__mux4_1 _18052_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[286] ),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[318] ),
    .A2(\gen_regfile_ff.register_file_i.rf_reg[350] ),
    .A3(\gen_regfile_ff.register_file_i.rf_reg[382] ),
    .S0(net1012),
    .S1(net1204),
    .X(_10785_));
 sky130_fd_sc_hd__mux2i_4 _18053_ (.A0(_10784_),
    .A1(_10785_),
    .S(_08529_),
    .Y(_10786_));
 sky130_fd_sc_hd__nand2_1 _18054_ (.A(net1140),
    .B(_10786_),
    .Y(_10787_));
 sky130_fd_sc_hd__and3_1 _18055_ (.A(_08512_),
    .B(_10783_),
    .C(_10787_),
    .X(_10788_));
 sky130_fd_sc_hd__a21oi_4 _18056_ (.A1(net383),
    .A2(_10777_),
    .B1(_10788_),
    .Y(_10789_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_849 ();
 sky130_fd_sc_hd__o22ai_1 _18058_ (.A1(_08502_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[62] ),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[30] ),
    .B2(_08503_),
    .Y(_10791_));
 sky130_fd_sc_hd__or3_4 _18059_ (.A(_10741_),
    .B(_10754_),
    .C(_10761_),
    .X(_10792_));
 sky130_fd_sc_hd__nor2_1 _18060_ (.A(_08504_),
    .B(_10792_),
    .Y(_10793_));
 sky130_fd_sc_hd__a2111o_1 _18061_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .A2(_10789_),
    .B1(_10791_),
    .C1(_10793_),
    .D1(net739),
    .X(_10794_));
 sky130_fd_sc_hd__o21ai_2 _18062_ (.A1(net313),
    .A2(_10765_),
    .B1(_10794_),
    .Y(_10795_));
 sky130_fd_sc_hd__nor2_1 _18063_ (.A(net310),
    .B(_10789_),
    .Y(_10796_));
 sky130_fd_sc_hd__a21oi_1 _18064_ (.A1(\cs_registers_i.pc_id_i[30] ),
    .A2(net310),
    .B1(_10796_),
    .Y(_10797_));
 sky130_fd_sc_hd__nand2_1 _18065_ (.A(\id_stage_i.controller_i.lsu_addr_last_i[30] ),
    .B(_08368_),
    .Y(_10798_));
 sky130_fd_sc_hd__o21ai_4 _18066_ (.A1(net933),
    .A2(_10797_),
    .B1(_10798_),
    .Y(_10799_));
 sky130_fd_sc_hd__and3_1 _18067_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[62] ),
    .B(_08272_),
    .C(_08377_),
    .X(_10800_));
 sky130_fd_sc_hd__a21oi_1 _18068_ (.A1(_08290_),
    .A2(_10799_),
    .B1(_10800_),
    .Y(_10801_));
 sky130_fd_sc_hd__or2_0 _18069_ (.A(_10565_),
    .B(_10597_),
    .X(_10802_));
 sky130_fd_sc_hd__a21oi_1 _18070_ (.A1(_10565_),
    .A2(_10597_),
    .B1(_10663_),
    .Y(_10803_));
 sky130_fd_sc_hd__o21ai_1 _18071_ (.A1(_10477_),
    .A2(_10660_),
    .B1(_10803_),
    .Y(_10804_));
 sky130_fd_sc_hd__nor4_4 _18072_ (.A(_10660_),
    .B(_10472_),
    .C(_10598_),
    .D(_10216_),
    .Y(_10805_));
 sky130_fd_sc_hd__a21oi_4 _18073_ (.A1(_10802_),
    .A2(_10804_),
    .B1(_10805_),
    .Y(_10806_));
 sky130_fd_sc_hd__maj3_2 _18074_ (.A(_10806_),
    .B(_10801_),
    .C(_10795_),
    .X(_10807_));
 sky130_fd_sc_hd__xnor2_4 _18075_ (.A(_10736_),
    .B(_10807_),
    .Y(net173));
 sky130_fd_sc_hd__xnor2_2 _18076_ (.A(_10795_),
    .B(_10801_),
    .Y(_10808_));
 sky130_fd_sc_hd__xnor2_4 _18077_ (.A(net779),
    .B(_10808_),
    .Y(_10809_));
 sky130_fd_sc_hd__clkinv_4 _18078_ (.A(_10809_),
    .Y(net172));
 sky130_fd_sc_hd__inv_8 _18079_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .Y(_10810_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_845 ();
 sky130_fd_sc_hd__nand3_4 _18084_ (.A(net442),
    .B(_08269_),
    .C(_08272_),
    .Y(_10815_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_841 ();
 sky130_fd_sc_hd__nor2b_1 _18089_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .B_N(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_10820_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_839 ();
 sky130_fd_sc_hd__nor2_1 _18092_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .Y(_10823_));
 sky130_fd_sc_hd__nand2_1 _18093_ (.A(_10820_),
    .B(_10823_),
    .Y(_10824_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_838 ();
 sky130_fd_sc_hd__nand2_1 _18095_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .B(_10815_),
    .Y(_10826_));
 sky130_fd_sc_hd__o41ai_1 _18096_ (.A1(_10810_),
    .A2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .A3(_10815_),
    .A4(_10824_),
    .B1(_10826_),
    .Y(_00002_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_830 ();
 sky130_fd_sc_hd__mux2i_1 _18105_ (.A0(net107),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_10835_));
 sky130_fd_sc_hd__mux2_1 _18106_ (.A0(net104),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_10836_));
 sky130_fd_sc_hd__nand2_1 _18107_ (.A(\cs_registers_i.pc_if_i[1] ),
    .B(_10836_),
    .Y(_10837_));
 sky130_fd_sc_hd__o21a_4 _18108_ (.A1(\cs_registers_i.pc_if_i[1] ),
    .A2(_10835_),
    .B1(_10837_),
    .X(_10838_));
 sky130_fd_sc_hd__clkinv_8 _18109_ (.A(_10838_),
    .Y(_10839_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_828 ();
 sky130_fd_sc_hd__mux2i_1 _18112_ (.A0(net96),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_10841_));
 sky130_fd_sc_hd__mux2_1 _18113_ (.A0(net103),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_10842_));
 sky130_fd_sc_hd__nand2_1 _18114_ (.A(net451),
    .B(_10842_),
    .Y(_10843_));
 sky130_fd_sc_hd__o21a_4 _18115_ (.A1(net451),
    .A2(_10841_),
    .B1(_10843_),
    .X(_10844_));
 sky130_fd_sc_hd__inv_6 _18116_ (.A(_10844_),
    .Y(\if_stage_i.compressed_decoder_i.instr_i[0] ));
 sky130_fd_sc_hd__nor2_2 _18117_ (.A(net25),
    .B(\load_store_unit_i.lsu_err_q ),
    .Y(_10845_));
 sky130_fd_sc_hd__nor2b_2 _18118_ (.A(\load_store_unit_i.ls_fsm_cs[0] ),
    .B_N(net59),
    .Y(_10846_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_827 ();
 sky130_fd_sc_hd__nor2_1 _18120_ (.A(\load_store_unit_i.ls_fsm_cs[2] ),
    .B(\load_store_unit_i.ls_fsm_cs[1] ),
    .Y(_10848_));
 sky130_fd_sc_hd__nand2_4 _18121_ (.A(_10846_),
    .B(_10848_),
    .Y(_10849_));
 sky130_fd_sc_hd__nor3_1 _18122_ (.A(\load_store_unit_i.data_we_q ),
    .B(_10845_),
    .C(_10849_),
    .Y(\id_stage_i.controller_i.load_err_d ));
 sky130_fd_sc_hd__nor2_2 _18123_ (.A(_10845_),
    .B(_10849_),
    .Y(_10850_));
 sky130_fd_sc_hd__and2_0 _18124_ (.A(\load_store_unit_i.data_we_q ),
    .B(_10850_),
    .X(\id_stage_i.controller_i.store_err_d ));
 sky130_fd_sc_hd__and3_2 _18125_ (.A(_08208_),
    .B(_08253_),
    .C(_08267_),
    .X(_10851_));
 sky130_fd_sc_hd__a22o_4 _18126_ (.A1(net920),
    .A2(_08450_),
    .B1(_09413_),
    .B2(_08495_),
    .X(_10852_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_826 ();
 sky130_fd_sc_hd__nand2_8 _18128_ (.A(_10851_),
    .B(_08632_),
    .Y(_10854_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_825 ();
 sky130_fd_sc_hd__nor2_4 _18130_ (.A(net1136),
    .B(_10854_),
    .Y(_10856_));
 sky130_fd_sc_hd__nand2_1 _18131_ (.A(net682),
    .B(_08190_),
    .Y(_10857_));
 sky130_fd_sc_hd__a211oi_4 _18132_ (.A1(_08416_),
    .A2(_10857_),
    .B1(_10854_),
    .C1(_08109_),
    .Y(_10858_));
 sky130_fd_sc_hd__inv_1 _18133_ (.A(\cs_registers_i.priv_lvl_q[1] ),
    .Y(_10859_));
 sky130_fd_sc_hd__nor2_1 _18134_ (.A(\cs_registers_i.priv_lvl_q[0] ),
    .B(net1143),
    .Y(_10860_));
 sky130_fd_sc_hd__o21ai_0 _18135_ (.A1(_10859_),
    .A2(_09261_),
    .B1(_10860_),
    .Y(_10861_));
 sky130_fd_sc_hd__nand2_1 _18136_ (.A(_10859_),
    .B(_09261_),
    .Y(_10862_));
 sky130_fd_sc_hd__a21oi_1 _18137_ (.A1(_10861_),
    .A2(_10862_),
    .B1(_10854_),
    .Y(_10863_));
 sky130_fd_sc_hd__a31o_1 _18138_ (.A1(_10852_),
    .A2(_10856_),
    .A3(_10858_),
    .B1(_10863_),
    .X(_10864_));
 sky130_fd_sc_hd__and4_4 _18139_ (.A(_09063_),
    .B(_09068_),
    .C(_09077_),
    .D(_09084_),
    .X(_10865_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_824 ();
 sky130_fd_sc_hd__nand2_1 _18141_ (.A(net583),
    .B(_08450_),
    .Y(_10867_));
 sky130_fd_sc_hd__o21ai_4 _18142_ (.A1(_08436_),
    .A2(_10865_),
    .B1(_10867_),
    .Y(_10868_));
 sky130_fd_sc_hd__nor2_8 _18143_ (.A(_08268_),
    .B(_08581_),
    .Y(_10869_));
 sky130_fd_sc_hd__nor2b_1 _18144_ (.A(net818),
    .B_N(net926),
    .Y(_10870_));
 sky130_fd_sc_hd__and3_1 _18145_ (.A(_10868_),
    .B(_10869_),
    .C(_10870_),
    .X(_10871_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_823 ();
 sky130_fd_sc_hd__nand4_1 _18147_ (.A(net814),
    .B(net674),
    .C(_08436_),
    .D(_08449_),
    .Y(_10873_));
 sky130_fd_sc_hd__nand2_1 _18148_ (.A(_09221_),
    .B(_09260_),
    .Y(_10874_));
 sky130_fd_sc_hd__nand2_4 _18149_ (.A(_10873_),
    .B(_10874_),
    .Y(_10875_));
 sky130_fd_sc_hd__nand2_4 _18150_ (.A(_10869_),
    .B(_10875_),
    .Y(_10876_));
 sky130_fd_sc_hd__nor3b_2 _18151_ (.A(_10876_),
    .B(net1145),
    .C_N(net1136),
    .Y(_10877_));
 sky130_fd_sc_hd__nand2b_4 _18152_ (.A_N(net1131),
    .B(net709),
    .Y(_10878_));
 sky130_fd_sc_hd__nand2_1 _18153_ (.A(_10869_),
    .B(_10878_),
    .Y(_10879_));
 sky130_fd_sc_hd__nor3_4 _18154_ (.A(_10852_),
    .B(_10856_),
    .C(_10876_),
    .Y(_10880_));
 sky130_fd_sc_hd__a31oi_1 _18155_ (.A1(\cs_registers_i.debug_mode_i ),
    .A2(_10877_),
    .A3(_10879_),
    .B1(_10880_),
    .Y(_10881_));
 sky130_fd_sc_hd__nand2_1 _18156_ (.A(_10880_),
    .B(_10879_),
    .Y(_10882_));
 sky130_fd_sc_hd__o21ai_2 _18157_ (.A1(net974),
    .A2(_10881_),
    .B1(_10882_),
    .Y(_10883_));
 sky130_fd_sc_hd__a21oi_2 _18158_ (.A1(net817),
    .A2(net925),
    .B1(_10854_),
    .Y(_10884_));
 sky130_fd_sc_hd__a21oi_1 _18159_ (.A1(net782),
    .A2(_08745_),
    .B1(_10854_),
    .Y(_10885_));
 sky130_fd_sc_hd__or2_2 _18160_ (.A(_10884_),
    .B(_10885_),
    .X(_10886_));
 sky130_fd_sc_hd__nor4_4 _18161_ (.A(_10852_),
    .B(_10856_),
    .C(_10876_),
    .D(_10886_),
    .Y(_10887_));
 sky130_fd_sc_hd__nor2_2 _18162_ (.A(net926),
    .B(_10885_),
    .Y(_10888_));
 sky130_fd_sc_hd__nand3_4 _18163_ (.A(net819),
    .B(_10880_),
    .C(_10888_),
    .Y(_10889_));
 sky130_fd_sc_hd__inv_1 _18164_ (.A(_10889_),
    .Y(_10890_));
 sky130_fd_sc_hd__nor2_2 _18165_ (.A(net639),
    .B(net723),
    .Y(_10891_));
 sky130_fd_sc_hd__nor3_4 _18166_ (.A(net1131),
    .B(net709),
    .C(_10854_),
    .Y(_10892_));
 sky130_fd_sc_hd__nand2_8 _18167_ (.A(_10891_),
    .B(_10892_),
    .Y(_10893_));
 sky130_fd_sc_hd__or2_2 _18168_ (.A(net636),
    .B(net728),
    .X(_10894_));
 sky130_fd_sc_hd__nor2_4 _18169_ (.A(_10894_),
    .B(_10878_),
    .Y(_10895_));
 sky130_fd_sc_hd__nor2_8 _18170_ (.A(_10854_),
    .B(_10895_),
    .Y(_10896_));
 sky130_fd_sc_hd__nand2_1 _18171_ (.A(_10893_),
    .B(_10896_),
    .Y(_10897_));
 sky130_fd_sc_hd__o21ai_1 _18172_ (.A1(_10887_),
    .A2(_10890_),
    .B1(_10897_),
    .Y(_10898_));
 sky130_fd_sc_hd__nor2_8 _18173_ (.A(_10854_),
    .B(_10878_),
    .Y(_10899_));
 sky130_fd_sc_hd__nand2_1 _18174_ (.A(_10894_),
    .B(_10899_),
    .Y(_10900_));
 sky130_fd_sc_hd__nor3_1 _18175_ (.A(_08898_),
    .B(_08639_),
    .C(_08900_),
    .Y(_10901_));
 sky130_fd_sc_hd__a21oi_4 _18176_ (.A1(net1085),
    .A2(_08495_),
    .B1(_10901_),
    .Y(_10902_));
 sky130_fd_sc_hd__nor2_4 _18177_ (.A(_10902_),
    .B(net724),
    .Y(_10903_));
 sky130_fd_sc_hd__nor2_1 _18178_ (.A(net783),
    .B(_10884_),
    .Y(_10904_));
 sky130_fd_sc_hd__nand2_2 _18179_ (.A(_10880_),
    .B(_10904_),
    .Y(_10905_));
 sky130_fd_sc_hd__nand2_4 _18180_ (.A(net964),
    .B(_10895_),
    .Y(_10906_));
 sky130_fd_sc_hd__nor2_8 _18181_ (.A(_10905_),
    .B(_10906_),
    .Y(_10907_));
 sky130_fd_sc_hd__a31oi_4 _18182_ (.A1(_10887_),
    .A2(_10903_),
    .A3(_10899_),
    .B1(_10907_),
    .Y(_10908_));
 sky130_fd_sc_hd__o21ai_1 _18183_ (.A1(_10889_),
    .A2(_10900_),
    .B1(_10908_),
    .Y(_10909_));
 sky130_fd_sc_hd__a21oi_1 _18184_ (.A1(net640),
    .A2(net723),
    .B1(_10878_),
    .Y(_10910_));
 sky130_fd_sc_hd__o21ai_0 _18185_ (.A1(_10854_),
    .A2(_10910_),
    .B1(_08745_),
    .Y(_10911_));
 sky130_fd_sc_hd__and3_1 _18186_ (.A(_10880_),
    .B(_10904_),
    .C(_10911_),
    .X(_10912_));
 sky130_fd_sc_hd__nand3_1 _18187_ (.A(net783),
    .B(_10852_),
    .C(_10869_),
    .Y(_10913_));
 sky130_fd_sc_hd__nor4_4 _18188_ (.A(net1136),
    .B(_10854_),
    .C(_10876_),
    .D(_10884_),
    .Y(_10914_));
 sky130_fd_sc_hd__nor4b_4 _18189_ (.A(_08745_),
    .B(_10893_),
    .C(_10913_),
    .D_N(_10914_),
    .Y(_10915_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_822 ();
 sky130_fd_sc_hd__nor2_1 _18191_ (.A(net820),
    .B(net723),
    .Y(_10917_));
 sky130_fd_sc_hd__and3_4 _18192_ (.A(_10892_),
    .B(_10887_),
    .C(_10903_),
    .X(_10918_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_821 ();
 sky130_fd_sc_hd__a41o_1 _18194_ (.A1(_10888_),
    .A2(_10899_),
    .A3(_10917_),
    .A4(_10877_),
    .B1(_10918_),
    .X(_10920_));
 sky130_fd_sc_hd__nor4_1 _18195_ (.A(_10909_),
    .B(_10912_),
    .C(_10915_),
    .D(_10920_),
    .Y(_10921_));
 sky130_fd_sc_hd__nand2_1 _18196_ (.A(_10898_),
    .B(_10921_),
    .Y(_10922_));
 sky130_fd_sc_hd__nand2_1 _18197_ (.A(_08745_),
    .B(_10903_),
    .Y(_10923_));
 sky130_fd_sc_hd__o21ai_1 _18198_ (.A1(_10878_),
    .A2(_10923_),
    .B1(net783),
    .Y(_10924_));
 sky130_fd_sc_hd__a21oi_4 _18199_ (.A1(_10869_),
    .A2(_10924_),
    .B1(_10852_),
    .Y(_10925_));
 sky130_fd_sc_hd__nand2_8 _18200_ (.A(_10914_),
    .B(_10925_),
    .Y(_10926_));
 sky130_fd_sc_hd__and3_4 _18201_ (.A(_10856_),
    .B(_10875_),
    .C(_10870_),
    .X(_10927_));
 sky130_fd_sc_hd__nand2_8 _18202_ (.A(_10925_),
    .B(_10927_),
    .Y(_10928_));
 sky130_fd_sc_hd__nand2_8 _18203_ (.A(_10926_),
    .B(_10928_),
    .Y(_10929_));
 sky130_fd_sc_hd__a211oi_4 _18204_ (.A1(_10871_),
    .A2(_10883_),
    .B1(_10922_),
    .C1(_10929_),
    .Y(_10930_));
 sky130_fd_sc_hd__o21ai_4 _18205_ (.A1(_10864_),
    .A2(_10930_),
    .B1(_10869_),
    .Y(_10931_));
 sky130_fd_sc_hd__nand2_1 _18206_ (.A(_10851_),
    .B(_10931_),
    .Y(_10932_));
 sky130_fd_sc_hd__nand2_1 _18207_ (.A(\id_stage_i.controller_i.instr_valid_i ),
    .B(_10932_),
    .Y(_10933_));
 sky130_fd_sc_hd__and3_2 _18208_ (.A(\id_stage_i.controller_i.instr_valid_i ),
    .B(_08206_),
    .C(net486),
    .X(_10934_));
 sky130_fd_sc_hd__nand4_4 _18209_ (.A(_08111_),
    .B(_08117_),
    .C(_08143_),
    .D(_10934_),
    .Y(_10935_));
 sky130_fd_sc_hd__nand3_1 _18210_ (.A(\cs_registers_i.csr_mstatus_tw_o ),
    .B(_08158_),
    .C(_10934_),
    .Y(_10936_));
 sky130_fd_sc_hd__and2_1 _18211_ (.A(\cs_registers_i.priv_lvl_q[0] ),
    .B(\cs_registers_i.priv_lvl_q[1] ),
    .X(_10937_));
 sky130_fd_sc_hd__a21oi_1 _18212_ (.A1(_10935_),
    .A2(_10936_),
    .B1(_10937_),
    .Y(_10938_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_820 ();
 sky130_fd_sc_hd__nor4_2 _18214_ (.A(net663),
    .B(net822),
    .C(_08121_),
    .D(_08123_),
    .Y(_10940_));
 sky130_fd_sc_hd__nand3_4 _18215_ (.A(_10940_),
    .B(_08143_),
    .C(_10934_),
    .Y(_10941_));
 sky130_fd_sc_hd__nor2_1 _18216_ (.A(\cs_registers_i.debug_mode_i ),
    .B(_10941_),
    .Y(_10942_));
 sky130_fd_sc_hd__nor2_1 _18217_ (.A(_10938_),
    .B(_10942_),
    .Y(_10943_));
 sky130_fd_sc_hd__nor2b_2 _18218_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .B_N(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .Y(_10944_));
 sky130_fd_sc_hd__nand2_8 _18219_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .B(_10944_),
    .Y(_10945_));
 sky130_fd_sc_hd__nor2_8 _18220_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .B(_10945_),
    .Y(_10946_));
 sky130_fd_sc_hd__a21oi_1 _18221_ (.A1(_10933_),
    .A2(_10943_),
    .B1(_10946_),
    .Y(\id_stage_i.controller_i.illegal_insn_d ));
 sky130_fd_sc_hd__a31o_2 _18222_ (.A1(_08164_),
    .A2(_08206_),
    .A3(net487),
    .B1(\id_stage_i.controller_i.instr_fetch_err_i ),
    .X(_10947_));
 sky130_fd_sc_hd__o21ai_0 _18223_ (.A1(_10932_),
    .A2(_10947_),
    .B1(\id_stage_i.controller_i.instr_valid_i ),
    .Y(_10948_));
 sky130_fd_sc_hd__a21oi_2 _18224_ (.A1(_10943_),
    .A2(_10948_),
    .B1(_10946_),
    .Y(\id_stage_i.controller_i.exc_req_d ));
 sky130_fd_sc_hd__nor3_1 _18225_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .B(_10815_),
    .C(_10824_),
    .Y(_10949_));
 sky130_fd_sc_hd__nand2_2 _18226_ (.A(net442),
    .B(_08272_),
    .Y(_10950_));
 sky130_fd_sc_hd__nor3_4 _18227_ (.A(_08109_),
    .B(_08268_),
    .C(_10950_),
    .Y(_10951_));
 sky130_fd_sc_hd__nand2_8 _18228_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .B(_10951_),
    .Y(_10952_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_818 ();
 sky130_fd_sc_hd__o21ai_0 _18231_ (.A1(_10810_),
    .A2(_10949_),
    .B1(_10952_),
    .Y(_00005_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_817 ();
 sky130_fd_sc_hd__inv_1 _18233_ (.A(_10400_),
    .Y(_10956_));
 sky130_fd_sc_hd__a311oi_1 _18234_ (.A1(_10341_),
    .A2(_10956_),
    .A3(_10402_),
    .B1(net992),
    .C1(net164),
    .Y(_10957_));
 sky130_fd_sc_hd__nor2_1 _18235_ (.A(net1560),
    .B(net1581),
    .Y(_10958_));
 sky130_fd_sc_hd__nand2_4 _18236_ (.A(net1278),
    .B(net881),
    .Y(_10959_));
 sky130_fd_sc_hd__xnor2_4 _18237_ (.A(_10959_),
    .B(_09118_),
    .Y(net176));
 sky130_fd_sc_hd__xor2_4 _18238_ (.A(_09295_),
    .B(_09296_),
    .X(net175));
 sky130_fd_sc_hd__nand2_1 _18239_ (.A(_08638_),
    .B(_08700_),
    .Y(_10960_));
 sky130_fd_sc_hd__nand2_1 _18240_ (.A(_08701_),
    .B(_10960_),
    .Y(_10961_));
 sky130_fd_sc_hd__xnor2_4 _18241_ (.A(_10961_),
    .B(_09294_),
    .Y(net174));
 sky130_fd_sc_hd__nand2_1 _18242_ (.A(_10341_),
    .B(_10474_),
    .Y(_10962_));
 sky130_fd_sc_hd__and3_1 _18243_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[32] ),
    .B(_08377_),
    .C(_08953_),
    .X(_10963_));
 sky130_fd_sc_hd__nor2_1 _18244_ (.A(_08956_),
    .B(_10963_),
    .Y(_10964_));
 sky130_fd_sc_hd__nand2_1 _18245_ (.A(_10902_),
    .B(_08953_),
    .Y(_10965_));
 sky130_fd_sc_hd__xnor2_1 _18246_ (.A(_08897_),
    .B(_10965_),
    .Y(_10966_));
 sky130_fd_sc_hd__nor2_2 _18247_ (.A(net1106),
    .B(_10966_),
    .Y(_10967_));
 sky130_fd_sc_hd__a21oi_4 _18248_ (.A1(net1107),
    .A2(_10964_),
    .B1(_10967_),
    .Y(_10968_));
 sky130_fd_sc_hd__xnor2_4 _18249_ (.A(net1110),
    .B(_09046_),
    .Y(_10969_));
 sky130_fd_sc_hd__xnor2_4 _18250_ (.A(_09039_),
    .B(_10969_),
    .Y(_10970_));
 sky130_fd_sc_hd__nor2_8 _18251_ (.A(_10968_),
    .B(_10970_),
    .Y(_10971_));
 sky130_fd_sc_hd__nor2_1 _18252_ (.A(_10341_),
    .B(_10403_),
    .Y(_10972_));
 sky130_fd_sc_hd__xor2_2 _18253_ (.A(_08844_),
    .B(_08852_),
    .X(_10973_));
 sky130_fd_sc_hd__xnor2_4 _18254_ (.A(_10973_),
    .B(_09047_),
    .Y(_10974_));
 sky130_fd_sc_hd__clkinv_8 _18255_ (.A(_10974_),
    .Y(net171));
 sky130_fd_sc_hd__a31oi_1 _18256_ (.A1(_10405_),
    .A2(_10401_),
    .A3(_10972_),
    .B1(net171),
    .Y(_10975_));
 sky130_fd_sc_hd__o2111ai_1 _18257_ (.A1(_10341_),
    .A2(_10956_),
    .B1(_10962_),
    .C1(_10971_),
    .D1(_10975_),
    .Y(_10976_));
 sky130_fd_sc_hd__or4_1 _18258_ (.A(net176),
    .B(net175),
    .C(net174),
    .D(_10976_),
    .X(_10977_));
 sky130_fd_sc_hd__or4_1 _18259_ (.A(net177),
    .B(net180),
    .C(net179),
    .D(_10977_),
    .X(_10978_));
 sky130_fd_sc_hd__nor4_2 _18260_ (.A(net152),
    .B(net1578),
    .C(net1583),
    .D(_10978_),
    .Y(_10979_));
 sky130_fd_sc_hd__nor4_1 _18261_ (.A(net178),
    .B(net154),
    .C(net153),
    .D(net721),
    .Y(_10980_));
 sky130_fd_sc_hd__nand3_1 _18262_ (.A(_10958_),
    .B(_10979_),
    .C(_10980_),
    .Y(_10981_));
 sky130_fd_sc_hd__or2_0 _18263_ (.A(net1241),
    .B(net1255),
    .X(_10982_));
 sky130_fd_sc_hd__a31o_1 _18264_ (.A1(net657),
    .A2(_10405_),
    .A3(_10972_),
    .B1(net1260),
    .X(_10983_));
 sky130_fd_sc_hd__nor4_2 _18265_ (.A(net689),
    .B(_10981_),
    .C(_10982_),
    .D(_10983_),
    .Y(_10984_));
 sky130_fd_sc_hd__nor2_1 _18266_ (.A(net165),
    .B(net687),
    .Y(_10985_));
 sky130_fd_sc_hd__nand4_1 _18267_ (.A(_10809_),
    .B(_10957_),
    .C(_10985_),
    .D(_10984_),
    .Y(_10986_));
 sky130_fd_sc_hd__nand2_1 _18268_ (.A(_10535_),
    .B(net851),
    .Y(_10987_));
 sky130_fd_sc_hd__nor4_4 _18269_ (.A(net493),
    .B(net482),
    .C(_10986_),
    .D(_10987_),
    .Y(_10988_));
 sky130_fd_sc_hd__nand2_1 _18270_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .B(_10951_),
    .Y(_10989_));
 sky130_fd_sc_hd__o22ai_1 _18271_ (.A1(_08500_),
    .A2(_10951_),
    .B1(_10988_),
    .B2(_10989_),
    .Y(_00004_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_815 ();
 sky130_fd_sc_hd__a21oi_1 _18274_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .A2(_10988_),
    .B1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .Y(_10992_));
 sky130_fd_sc_hd__nand2_1 _18275_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_valid ),
    .B(_10815_),
    .Y(_10993_));
 sky130_fd_sc_hd__o21ai_0 _18276_ (.A1(_10815_),
    .A2(_10992_),
    .B1(_10993_),
    .Y(_00003_));
 sky130_fd_sc_hd__inv_6 _18277_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .Y(_10994_));
 sky130_fd_sc_hd__nor3_4 _18278_ (.A(\id_stage_i.controller_i.store_err_q ),
    .B(\id_stage_i.controller_i.exc_req_q ),
    .C(\id_stage_i.controller_i.load_err_q ),
    .Y(_10995_));
 sky130_fd_sc_hd__nand3_4 _18279_ (.A(_10935_),
    .B(_10941_),
    .C(_10995_),
    .Y(_10996_));
 sky130_fd_sc_hd__nor2_1 _18280_ (.A(\cs_registers_i.priv_lvl_q[0] ),
    .B(\cs_registers_i.priv_lvl_q[1] ),
    .Y(_10997_));
 sky130_fd_sc_hd__a22o_1 _18281_ (.A1(\cs_registers_i.dcsr_q[15] ),
    .A2(_10937_),
    .B1(_10997_),
    .B2(\cs_registers_i.dcsr_q[12] ),
    .X(_10998_));
 sky130_fd_sc_hd__nor2_1 _18282_ (.A(\cs_registers_i.debug_mode_i ),
    .B(_10998_),
    .Y(_10999_));
 sky130_fd_sc_hd__and3_1 _18283_ (.A(\id_stage_i.controller_i.instr_valid_i ),
    .B(_08206_),
    .C(net485),
    .X(_11000_));
 sky130_fd_sc_hd__nor2_1 _18284_ (.A(\id_stage_i.controller_i.instr_fetch_err_i ),
    .B(\id_stage_i.controller_i.illegal_insn_q ),
    .Y(_11001_));
 sky130_fd_sc_hd__nand4_4 _18285_ (.A(net382),
    .B(_08164_),
    .C(_11000_),
    .D(_11001_),
    .Y(_11002_));
 sky130_fd_sc_hd__nor3_2 _18286_ (.A(_10995_),
    .B(_10999_),
    .C(_11002_),
    .Y(_11003_));
 sky130_fd_sc_hd__nor3_2 _18287_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .B(_10945_),
    .C(_11003_),
    .Y(_11004_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_814 ();
 sky130_fd_sc_hd__or3_4 _18289_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .B(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .C(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .X(_11006_));
 sky130_fd_sc_hd__nor2_1 _18290_ (.A(\cs_registers_i.dcsr_q[2] ),
    .B(net60),
    .Y(_11007_));
 sky130_fd_sc_hd__nor2_2 _18291_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .B(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .Y(_11008_));
 sky130_fd_sc_hd__nand2_8 _18292_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .B(_11008_),
    .Y(_11009_));
 sky130_fd_sc_hd__a21o_1 _18293_ (.A1(_08104_),
    .A2(_11007_),
    .B1(_11009_),
    .X(_11010_));
 sky130_fd_sc_hd__nand2_1 _18294_ (.A(_11006_),
    .B(_11010_),
    .Y(_11011_));
 sky130_fd_sc_hd__and2_2 _18295_ (.A(\cs_registers_i.mie_q[14] ),
    .B(net135),
    .X(_11012_));
 sky130_fd_sc_hd__a22oi_4 _18296_ (.A1(\cs_registers_i.mie_q[4] ),
    .A2(net139),
    .B1(\cs_registers_i.mie_q[5] ),
    .B2(net140),
    .Y(_11013_));
 sky130_fd_sc_hd__and2_0 _18297_ (.A(\cs_registers_i.mie_q[6] ),
    .B(net141),
    .X(_11014_));
 sky130_fd_sc_hd__a21oi_2 _18298_ (.A1(\cs_registers_i.mie_q[7] ),
    .A2(net142),
    .B1(_11014_),
    .Y(_11015_));
 sky130_fd_sc_hd__a22oi_4 _18299_ (.A1(\cs_registers_i.mie_q[2] ),
    .A2(net137),
    .B1(\cs_registers_i.mie_q[3] ),
    .B2(net138),
    .Y(_11016_));
 sky130_fd_sc_hd__a22oi_2 _18300_ (.A1(\cs_registers_i.mie_q[0] ),
    .A2(net130),
    .B1(\cs_registers_i.mie_q[1] ),
    .B2(net136),
    .Y(_11017_));
 sky130_fd_sc_hd__nand4_4 _18301_ (.A(_11013_),
    .B(_11015_),
    .C(_11016_),
    .D(_11017_),
    .Y(_11018_));
 sky130_fd_sc_hd__nand2_1 _18302_ (.A(\cs_registers_i.mie_q[13] ),
    .B(net134),
    .Y(_11019_));
 sky130_fd_sc_hd__nand2_1 _18303_ (.A(\cs_registers_i.mie_q[12] ),
    .B(net133),
    .Y(_11020_));
 sky130_fd_sc_hd__and2_2 _18304_ (.A(_11019_),
    .B(_11020_),
    .X(_11021_));
 sky130_fd_sc_hd__and2_0 _18305_ (.A(\cs_registers_i.mie_q[11] ),
    .B(net132),
    .X(_11022_));
 sky130_fd_sc_hd__a21o_1 _18306_ (.A1(\cs_registers_i.mie_q[10] ),
    .A2(net131),
    .B1(_11022_),
    .X(_11023_));
 sky130_fd_sc_hd__a221oi_4 _18307_ (.A1(\cs_registers_i.mie_q[8] ),
    .A2(net143),
    .B1(\cs_registers_i.mie_q[9] ),
    .B2(net144),
    .C1(_11023_),
    .Y(_11024_));
 sky130_fd_sc_hd__nand2_1 _18308_ (.A(_11021_),
    .B(_11024_),
    .Y(_11025_));
 sky130_fd_sc_hd__nor3_2 _18309_ (.A(_11012_),
    .B(_11018_),
    .C(_11025_),
    .Y(_11026_));
 sky130_fd_sc_hd__nand2_1 _18310_ (.A(net129),
    .B(\cs_registers_i.mie_q[15] ),
    .Y(_11027_));
 sky130_fd_sc_hd__nand2_1 _18311_ (.A(\cs_registers_i.mie_q[17] ),
    .B(net146),
    .Y(_11028_));
 sky130_fd_sc_hd__nand3_2 _18312_ (.A(_11026_),
    .B(_11027_),
    .C(_11028_),
    .Y(_11029_));
 sky130_fd_sc_hd__a211oi_4 _18313_ (.A1(\cs_registers_i.mie_q[16] ),
    .A2(net147),
    .B1(_11029_),
    .C1(net145),
    .Y(_11030_));
 sky130_fd_sc_hd__nand2b_1 _18314_ (.A_N(\cs_registers_i.debug_mode_i ),
    .B(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .Y(_11031_));
 sky130_fd_sc_hd__clkinv_2 _18315_ (.A(\cs_registers_i.nmi_mode_i ),
    .Y(_11032_));
 sky130_fd_sc_hd__o21ai_4 _18316_ (.A1(net145),
    .A2(\cs_registers_i.csr_mstatus_mie_o ),
    .B1(_11032_),
    .Y(_11033_));
 sky130_fd_sc_hd__nor4_4 _18317_ (.A(_10945_),
    .B(_11030_),
    .C(_11031_),
    .D(_11033_),
    .Y(_11034_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_813 ();
 sky130_fd_sc_hd__nor2_4 _18319_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .B(_08106_),
    .Y(_11036_));
 sky130_fd_sc_hd__nand2_8 _18320_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .B(_11036_),
    .Y(_11037_));
 sky130_fd_sc_hd__a21oi_1 _18321_ (.A1(_08443_),
    .A2(_08440_),
    .B1(\id_stage_i.id_fsm_q ),
    .Y(_11038_));
 sky130_fd_sc_hd__a21oi_2 _18322_ (.A1(_08269_),
    .A2(_11038_),
    .B1(\id_stage_i.branch_set ),
    .Y(_11039_));
 sky130_fd_sc_hd__and2_4 _18323_ (.A(\id_stage_i.controller_i.instr_valid_i ),
    .B(\id_stage_i.controller_i.instr_fetch_err_i ),
    .X(_11040_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_812 ();
 sky130_fd_sc_hd__nor3_4 _18325_ (.A(_11037_),
    .B(_11039_),
    .C(_11040_),
    .Y(_11042_));
 sky130_fd_sc_hd__a2111o_4 _18326_ (.A1(_10996_),
    .A2(_11004_),
    .B1(_11042_),
    .C1(_11034_),
    .D1(_11011_),
    .X(_11043_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_807 ();
 sky130_fd_sc_hd__nor2_1 _18332_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q ),
    .B(net1026),
    .Y(_11049_));
 sky130_fd_sc_hd__nor2_1 _18333_ (.A(_10994_),
    .B(_11049_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ));
 sky130_fd_sc_hd__mux2i_1 _18334_ (.A0(net100),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_11050_));
 sky130_fd_sc_hd__mux2_1 _18335_ (.A0(net117),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_11051_));
 sky130_fd_sc_hd__nand2_1 _18336_ (.A(net451),
    .B(_11051_),
    .Y(_11052_));
 sky130_fd_sc_hd__o21a_4 _18337_ (.A1(net451),
    .A2(_11050_),
    .B1(_11052_),
    .X(_11053_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_806 ();
 sky130_fd_sc_hd__inv_8 _18339_ (.A(_11053_),
    .Y(_11055_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_805 ();
 sky130_fd_sc_hd__mux2i_1 _18341_ (.A0(net101),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_11056_));
 sky130_fd_sc_hd__mux2_1 _18342_ (.A0(net119),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_11057_));
 sky130_fd_sc_hd__nand2_1 _18343_ (.A(net451),
    .B(_11057_),
    .Y(_11058_));
 sky130_fd_sc_hd__o21a_4 _18344_ (.A1(net451),
    .A2(_11056_),
    .B1(_11058_),
    .X(_11059_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_804 ();
 sky130_fd_sc_hd__inv_12 _18346_ (.A(_11059_),
    .Y(_11061_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_801 ();
 sky130_fd_sc_hd__mux2i_1 _18350_ (.A0(net102),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_11064_));
 sky130_fd_sc_hd__mux2_1 _18351_ (.A0(net120),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_11065_));
 sky130_fd_sc_hd__nand2_1 _18352_ (.A(net451),
    .B(_11065_),
    .Y(_11066_));
 sky130_fd_sc_hd__o21a_4 _18353_ (.A1(net451),
    .A2(_11064_),
    .B1(_11066_),
    .X(_11067_));
 sky130_fd_sc_hd__inv_8 _18354_ (.A(_11067_),
    .Y(_11068_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_799 ();
 sky130_fd_sc_hd__mux2i_1 _18357_ (.A0(net97),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_11070_));
 sky130_fd_sc_hd__mux2_1 _18358_ (.A0(net114),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_11071_));
 sky130_fd_sc_hd__nand2_1 _18359_ (.A(net450),
    .B(_11071_),
    .Y(_11072_));
 sky130_fd_sc_hd__o21a_2 _18360_ (.A1(net450),
    .A2(_11070_),
    .B1(_11072_),
    .X(_11073_));
 sky130_fd_sc_hd__inv_6 _18361_ (.A(_11073_),
    .Y(_11074_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_798 ();
 sky130_fd_sc_hd__mux2i_2 _18363_ (.A0(net98),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_11075_));
 sky130_fd_sc_hd__mux2_1 _18364_ (.A0(net115),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_11076_));
 sky130_fd_sc_hd__nand2_1 _18365_ (.A(net450),
    .B(_11076_),
    .Y(_11077_));
 sky130_fd_sc_hd__o21ai_4 _18366_ (.A1(net450),
    .A2(_11075_),
    .B1(_11077_),
    .Y(_11078_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_797 ();
 sky130_fd_sc_hd__mux2i_2 _18368_ (.A0(net123),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_11079_));
 sky130_fd_sc_hd__mux2_1 _18369_ (.A0(net109),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_11080_));
 sky130_fd_sc_hd__nand2_1 _18370_ (.A(net449),
    .B(_11080_),
    .Y(_11081_));
 sky130_fd_sc_hd__o21ai_4 _18371_ (.A1(net449),
    .A2(_11079_),
    .B1(_11081_),
    .Y(_11082_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_796 ();
 sky130_fd_sc_hd__mux2i_1 _18373_ (.A0(net124),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_11083_));
 sky130_fd_sc_hd__mux2_1 _18374_ (.A0(net110),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_11084_));
 sky130_fd_sc_hd__nand2_1 _18375_ (.A(net449),
    .B(_11084_),
    .Y(_11085_));
 sky130_fd_sc_hd__o21a_4 _18376_ (.A1(net449),
    .A2(_11083_),
    .B1(_11085_),
    .X(_11086_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_795 ();
 sky130_fd_sc_hd__inv_2 _18378_ (.A(_11086_),
    .Y(\if_stage_i.compressed_decoder_i.instr_i[6] ));
 sky130_fd_sc_hd__mux2i_2 _18379_ (.A0(net118),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_11088_));
 sky130_fd_sc_hd__mux2_1 _18380_ (.A0(net105),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_11089_));
 sky130_fd_sc_hd__nand2_1 _18381_ (.A(net449),
    .B(_11089_),
    .Y(_11090_));
 sky130_fd_sc_hd__o21ai_4 _18382_ (.A1(net449),
    .A2(_11088_),
    .B1(_11090_),
    .Y(_11091_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_794 ();
 sky130_fd_sc_hd__mux2i_2 _18384_ (.A0(net121),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_11092_));
 sky130_fd_sc_hd__mux2_1 _18385_ (.A0(net106),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_11093_));
 sky130_fd_sc_hd__nand2_1 _18386_ (.A(net450),
    .B(_11093_),
    .Y(_11094_));
 sky130_fd_sc_hd__o21ai_4 _18387_ (.A1(net450),
    .A2(_11092_),
    .B1(_11094_),
    .Y(_11095_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_793 ();
 sky130_fd_sc_hd__mux2i_1 _18389_ (.A0(net122),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_11096_));
 sky130_fd_sc_hd__mux2_1 _18390_ (.A0(net108),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_11097_));
 sky130_fd_sc_hd__nand2_1 _18391_ (.A(net449),
    .B(_11097_),
    .Y(_11098_));
 sky130_fd_sc_hd__o21a_2 _18392_ (.A1(net449),
    .A2(_11096_),
    .B1(_11098_),
    .X(_11099_));
 sky130_fd_sc_hd__inv_4 _18393_ (.A(_11099_),
    .Y(\if_stage_i.compressed_decoder_i.instr_i[4] ));
 sky130_fd_sc_hd__mux2i_2 _18394_ (.A0(net125),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_11100_));
 sky130_fd_sc_hd__mux2_1 _18395_ (.A0(net111),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_11101_));
 sky130_fd_sc_hd__nand2_1 _18396_ (.A(net449),
    .B(_11101_),
    .Y(_11102_));
 sky130_fd_sc_hd__o21ai_4 _18397_ (.A1(net449),
    .A2(_11100_),
    .B1(_11102_),
    .Y(_11103_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_792 ();
 sky130_fd_sc_hd__mux2i_2 _18399_ (.A0(net126),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_11104_));
 sky130_fd_sc_hd__mux2_1 _18400_ (.A0(net112),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_11105_));
 sky130_fd_sc_hd__nand2_1 _18401_ (.A(net450),
    .B(_11105_),
    .Y(_11106_));
 sky130_fd_sc_hd__o21ai_4 _18402_ (.A1(net450),
    .A2(_11104_),
    .B1(_11106_),
    .Y(_11107_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_791 ();
 sky130_fd_sc_hd__mux2i_2 _18404_ (.A0(net127),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_11108_));
 sky130_fd_sc_hd__mux2_1 _18405_ (.A0(net113),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_11109_));
 sky130_fd_sc_hd__nand2_1 _18406_ (.A(net450),
    .B(_11109_),
    .Y(_11110_));
 sky130_fd_sc_hd__o21ai_4 _18407_ (.A1(net450),
    .A2(_11108_),
    .B1(_11110_),
    .Y(\if_stage_i.compressed_decoder_i.instr_i[9] ));
 sky130_fd_sc_hd__mux2i_1 _18408_ (.A0(net99),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_11111_));
 sky130_fd_sc_hd__mux2_1 _18409_ (.A0(net116),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_11112_));
 sky130_fd_sc_hd__nand2_1 _18410_ (.A(net451),
    .B(_11112_),
    .Y(_11113_));
 sky130_fd_sc_hd__o21a_4 _18411_ (.A1(net451),
    .A2(_11111_),
    .B1(_11113_),
    .X(_11114_));
 sky130_fd_sc_hd__inv_6 _18412_ (.A(_11114_),
    .Y(_11115_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_788 ();
 sky130_fd_sc_hd__mux2_1 _18416_ (.A0(net96),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[0] ));
 sky130_fd_sc_hd__mux2_1 _18417_ (.A0(net107),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[1] ));
 sky130_fd_sc_hd__mux2i_4 _18418_ (.A0(net118),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Y(_11118_));
 sky130_fd_sc_hd__inv_1 _18419_ (.A(_11118_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[2] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_787 ();
 sky130_fd_sc_hd__mux2_1 _18421_ (.A0(net121),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[3] ));
 sky130_fd_sc_hd__mux2i_2 _18422_ (.A0(net122),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Y(_11120_));
 sky130_fd_sc_hd__inv_1 _18423_ (.A(_11120_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[4] ));
 sky130_fd_sc_hd__mux2_1 _18424_ (.A0(net123),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[5] ));
 sky130_fd_sc_hd__mux2_1 _18425_ (.A0(net124),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[6] ));
 sky130_fd_sc_hd__mux2i_1 _18426_ (.A0(net125),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Y(_11121_));
 sky130_fd_sc_hd__inv_1 _18427_ (.A(_11121_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[7] ));
 sky130_fd_sc_hd__mux2_1 _18428_ (.A0(net126),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[8] ));
 sky130_fd_sc_hd__mux2i_1 _18429_ (.A0(net127),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Y(_11122_));
 sky130_fd_sc_hd__inv_1 _18430_ (.A(_11122_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[9] ));
 sky130_fd_sc_hd__mux2_1 _18431_ (.A0(net97),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[10] ));
 sky130_fd_sc_hd__mux2i_1 _18432_ (.A0(net98),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Y(_11123_));
 sky130_fd_sc_hd__inv_1 _18433_ (.A(_11123_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[11] ));
 sky130_fd_sc_hd__mux2i_1 _18434_ (.A0(net99),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Y(_11124_));
 sky130_fd_sc_hd__inv_1 _18435_ (.A(_11124_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[12] ));
 sky130_fd_sc_hd__mux2_1 _18436_ (.A0(net100),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[13] ));
 sky130_fd_sc_hd__mux2i_1 _18437_ (.A0(net101),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Y(_11125_));
 sky130_fd_sc_hd__inv_1 _18438_ (.A(_11125_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[14] ));
 sky130_fd_sc_hd__mux2_1 _18439_ (.A0(net102),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[15] ));
 sky130_fd_sc_hd__clkinvlp_4 _18440_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Y(_11126_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_784 ();
 sky130_fd_sc_hd__nand2_2 _18444_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .B(net128),
    .Y(_11130_));
 sky130_fd_sc_hd__nor4_4 _18445_ (.A(_11126_),
    .B(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .C(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .D(_11130_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[2] ));
 sky130_fd_sc_hd__nor2_1 _18446_ (.A(net60),
    .B(core_busy_q),
    .Y(_11131_));
 sky130_fd_sc_hd__nand2_2 _18447_ (.A(_11030_),
    .B(_11131_),
    .Y(_11132_));
 sky130_fd_sc_hd__nand2_1 _18448_ (.A(fetch_enable_q),
    .B(_11132_),
    .Y(net150));
 sky130_fd_sc_hd__nand2b_1 _18449_ (.A_N(net149),
    .B(net150),
    .Y(_00006_));
 sky130_fd_sc_hd__nand2_1 _18450_ (.A(net103),
    .B(net104),
    .Y(_11133_));
 sky130_fd_sc_hd__nor2_1 _18451_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .B(_11133_),
    .Y(_11134_));
 sky130_fd_sc_hd__a31oi_1 _18452_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .A2(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ),
    .A3(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ),
    .B1(_11134_),
    .Y(_11135_));
 sky130_fd_sc_hd__mux2i_1 _18453_ (.A0(net94),
    .A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ),
    .S(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .Y(_11136_));
 sky130_fd_sc_hd__nand2_1 _18454_ (.A(_11135_),
    .B(_11136_),
    .Y(_11137_));
 sky130_fd_sc_hd__and2_1 _18455_ (.A(\cs_registers_i.pc_if_i[1] ),
    .B(_11137_),
    .X(_11138_));
 sky130_fd_sc_hd__nor2_2 _18456_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .B(_11130_),
    .Y(_11139_));
 sky130_fd_sc_hd__nor2_1 _18457_ (.A(_11139_),
    .B(_11138_),
    .Y(_11140_));
 sky130_fd_sc_hd__a21oi_1 _18458_ (.A1(_11126_),
    .A2(_11138_),
    .B1(_11140_),
    .Y(_11141_));
 sky130_fd_sc_hd__nand2_1 _18459_ (.A(_10935_),
    .B(_10941_),
    .Y(_11142_));
 sky130_fd_sc_hd__nand2_1 _18460_ (.A(_08158_),
    .B(_11000_),
    .Y(_11143_));
 sky130_fd_sc_hd__o21ai_1 _18461_ (.A1(_10845_),
    .A2(_10849_),
    .B1(_11143_),
    .Y(_11144_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_783 ();
 sky130_fd_sc_hd__and3_4 _18463_ (.A(net682),
    .B(_08190_),
    .C(_08206_),
    .X(_11146_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_782 ();
 sky130_fd_sc_hd__nand2_8 _18465_ (.A(net491),
    .B(_11146_),
    .Y(_11148_));
 sky130_fd_sc_hd__nor3_1 _18466_ (.A(net554),
    .B(_08124_),
    .C(_11148_),
    .Y(_11149_));
 sky130_fd_sc_hd__nand3_4 _18467_ (.A(net683),
    .B(_08190_),
    .C(_08206_),
    .Y(_11150_));
 sky130_fd_sc_hd__nor2_8 _18468_ (.A(_08254_),
    .B(_11150_),
    .Y(_11151_));
 sky130_fd_sc_hd__nor4_1 _18469_ (.A(net382),
    .B(net372),
    .C(_08118_),
    .D(_11151_),
    .Y(_11152_));
 sky130_fd_sc_hd__inv_1 _18470_ (.A(_08139_),
    .Y(_11153_));
 sky130_fd_sc_hd__o2111ai_4 _18471_ (.A1(_11149_),
    .A2(_11152_),
    .B1(\id_stage_i.controller_i.instr_valid_i ),
    .C1(_11153_),
    .D1(_10858_),
    .Y(_11154_));
 sky130_fd_sc_hd__nor4b_4 _18472_ (.A(\id_stage_i.controller_i.exc_req_d ),
    .B(_11142_),
    .C(_11144_),
    .D_N(_11154_),
    .Y(_11155_));
 sky130_fd_sc_hd__nor3_2 _18473_ (.A(\cs_registers_i.debug_mode_i ),
    .B(_11030_),
    .C(_11033_),
    .Y(_11156_));
 sky130_fd_sc_hd__a21oi_2 _18474_ (.A1(\id_stage_i.controller_i.instr_valid_i ),
    .A2(\cs_registers_i.dcsr_q[2] ),
    .B1(net60),
    .Y(_11157_));
 sky130_fd_sc_hd__nor2_4 _18475_ (.A(\cs_registers_i.debug_mode_i ),
    .B(_11157_),
    .Y(_11158_));
 sky130_fd_sc_hd__o221ai_4 _18476_ (.A1(_08104_),
    .A2(_11155_),
    .B1(_11156_),
    .B2(_11158_),
    .C1(_11036_),
    .Y(_11159_));
 sky130_fd_sc_hd__nor2_1 _18477_ (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .B(_11139_),
    .Y(_11160_));
 sky130_fd_sc_hd__inv_1 _18478_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .Y(_11161_));
 sky130_fd_sc_hd__and2_1 _18479_ (.A(_11161_),
    .B(_10944_),
    .X(_11162_));
 sky130_fd_sc_hd__a211oi_1 _18480_ (.A1(_11138_),
    .A2(_11160_),
    .B1(_11162_),
    .C1(_10946_),
    .Y(_11163_));
 sky130_fd_sc_hd__o211ai_4 _18481_ (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .A2(_11141_),
    .B1(_11159_),
    .C1(_11163_),
    .Y(_11164_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_780 ();
 sky130_fd_sc_hd__xor2_1 _18484_ (.A(_10695_),
    .B(_10724_),
    .X(_11167_));
 sky130_fd_sc_hd__o21ai_2 _18485_ (.A1(_08385_),
    .A2(_08386_),
    .B1(_08233_),
    .Y(_11168_));
 sky130_fd_sc_hd__a211oi_2 _18486_ (.A1(net1091),
    .A2(_08394_),
    .B1(_08410_),
    .C1(_08224_),
    .Y(_11169_));
 sky130_fd_sc_hd__a21oi_1 _18487_ (.A1(_08396_),
    .A2(_08400_),
    .B1(_08265_),
    .Y(_11170_));
 sky130_fd_sc_hd__nor4_4 _18488_ (.A(_11168_),
    .B(_08404_),
    .C(_11169_),
    .D(_11170_),
    .Y(_11171_));
 sky130_fd_sc_hd__xor2_1 _18489_ (.A(_08424_),
    .B(_11171_),
    .X(_11172_));
 sky130_fd_sc_hd__nor4_1 _18490_ (.A(_08410_),
    .B(_08387_),
    .C(net644),
    .D(_11172_),
    .Y(_11173_));
 sky130_fd_sc_hd__nor2_1 _18491_ (.A(_08410_),
    .B(_08387_),
    .Y(_11174_));
 sky130_fd_sc_hd__nor2b_1 _18492_ (.A(_08424_),
    .B_N(_11171_),
    .Y(_11175_));
 sky130_fd_sc_hd__o21ai_0 _18493_ (.A1(_08410_),
    .A2(_08387_),
    .B1(_08429_),
    .Y(_11176_));
 sky130_fd_sc_hd__a21boi_0 _18494_ (.A1(_11174_),
    .A2(_11175_),
    .B1_N(_11176_),
    .Y(_11177_));
 sky130_fd_sc_hd__nand3b_1 _18495_ (.A_N(_11171_),
    .B(_08423_),
    .C(net644),
    .Y(_11178_));
 sky130_fd_sc_hd__o21ai_1 _18496_ (.A1(net644),
    .A2(_11177_),
    .B1(_11178_),
    .Y(_11179_));
 sky130_fd_sc_hd__mux2_1 _18497_ (.A0(_11173_),
    .A1(_11179_),
    .S(net173),
    .X(_11180_));
 sky130_fd_sc_hd__nand2b_1 _18498_ (.A_N(net644),
    .B(_11171_),
    .Y(_11181_));
 sky130_fd_sc_hd__o21ai_1 _18499_ (.A1(_11176_),
    .A2(_11181_),
    .B1(_11178_),
    .Y(_11182_));
 sky130_fd_sc_hd__nand2_1 _18500_ (.A(_08428_),
    .B(_11181_),
    .Y(_11183_));
 sky130_fd_sc_hd__a21oi_1 _18501_ (.A1(_08423_),
    .A2(_11183_),
    .B1(_11179_),
    .Y(_11184_));
 sky130_fd_sc_hd__nand2_1 _18502_ (.A(_08423_),
    .B(_11183_),
    .Y(_11185_));
 sky130_fd_sc_hd__o2111ai_1 _18503_ (.A1(_11173_),
    .A2(_11182_),
    .B1(_11185_),
    .C1(_10724_),
    .D1(_10695_),
    .Y(_11186_));
 sky130_fd_sc_hd__o41ai_1 _18504_ (.A1(_10695_),
    .A2(_10724_),
    .A3(_11182_),
    .A4(_11184_),
    .B1(_11186_),
    .Y(_11187_));
 sky130_fd_sc_hd__a21oi_1 _18505_ (.A1(_11167_),
    .A2(_11180_),
    .B1(_11187_),
    .Y(_11188_));
 sky130_fd_sc_hd__nor3_1 _18506_ (.A(net1089),
    .B(_08416_),
    .C(_08410_),
    .Y(_11189_));
 sky130_fd_sc_hd__nor3_1 _18507_ (.A(_11173_),
    .B(_11179_),
    .C(_11189_),
    .Y(_11190_));
 sky130_fd_sc_hd__mux2i_1 _18508_ (.A0(_11189_),
    .A1(_11190_),
    .S(_10988_),
    .Y(_11191_));
 sky130_fd_sc_hd__nand2_2 _18509_ (.A(_11191_),
    .B(_11188_),
    .Y(_11192_));
 sky130_fd_sc_hd__nand2_4 _18510_ (.A(_11192_),
    .B(_08409_),
    .Y(_11193_));
 sky130_fd_sc_hd__nor4_4 _18511_ (.A(\id_stage_i.id_fsm_q ),
    .B(_08109_),
    .C(_08268_),
    .D(_11193_),
    .Y(\id_stage_i.branch_set_d ));
 sky130_fd_sc_hd__inv_1 _18512_ (.A(\id_stage_i.id_fsm_q ),
    .Y(_11194_));
 sky130_fd_sc_hd__nor2_2 _18513_ (.A(_08214_),
    .B(_08268_),
    .Y(_11195_));
 sky130_fd_sc_hd__o211ai_1 _18514_ (.A1(_11194_),
    .A2(_10849_),
    .B1(_11195_),
    .C1(\id_stage_i.controller_i.instr_valid_i ),
    .Y(_11196_));
 sky130_fd_sc_hd__a2111oi_4 _18515_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .A2(net490),
    .B1(net739),
    .C1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .D1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_valid ),
    .Y(_11197_));
 sky130_fd_sc_hd__o21ai_0 _18516_ (.A1(_11038_),
    .A2(_11197_),
    .B1(_08269_),
    .Y(_11198_));
 sky130_fd_sc_hd__nand2_2 _18517_ (.A(_11196_),
    .B(_11198_),
    .Y(_11199_));
 sky130_fd_sc_hd__nor2_8 _18518_ (.A(_11199_),
    .B(\id_stage_i.branch_set_d ),
    .Y(_11200_));
 sky130_fd_sc_hd__o21ai_4 _18519_ (.A1(_11037_),
    .A2(_11155_),
    .B1(_11200_),
    .Y(_11201_));
 sky130_fd_sc_hd__nor2_8 _18520_ (.A(_11201_),
    .B(_11164_),
    .Y(_00007_));
 sky130_fd_sc_hd__nor2_1 _18521_ (.A(\id_stage_i.id_fsm_q ),
    .B(_08109_),
    .Y(_11202_));
 sky130_fd_sc_hd__nand2_1 _18522_ (.A(_11202_),
    .B(_11195_),
    .Y(_11203_));
 sky130_fd_sc_hd__nor2_1 _18523_ (.A(\load_store_unit_i.ls_fsm_cs[1] ),
    .B(_11203_),
    .Y(_11204_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_779 ();
 sky130_fd_sc_hd__nor2b_2 _18525_ (.A(\load_store_unit_i.ls_fsm_cs[2] ),
    .B_N(net26),
    .Y(_11206_));
 sky130_fd_sc_hd__o21ai_4 _18526_ (.A1(\load_store_unit_i.ls_fsm_cs[0] ),
    .A2(_11204_),
    .B1(_11206_),
    .Y(_11207_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_778 ();
 sky130_fd_sc_hd__nand2_1 _18528_ (.A(\load_store_unit_i.data_type_q[2] ),
    .B(_11207_),
    .Y(_11209_));
 sky130_fd_sc_hd__o31ai_1 _18529_ (.A1(_08416_),
    .A2(_08214_),
    .A3(_11207_),
    .B1(_11209_),
    .Y(_00008_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_777 ();
 sky130_fd_sc_hd__nand2_1 _18531_ (.A(\load_store_unit_i.data_type_q[1] ),
    .B(_11207_),
    .Y(_11211_));
 sky130_fd_sc_hd__o41ai_1 _18532_ (.A1(net491),
    .A2(net678),
    .A3(_08214_),
    .A4(_11207_),
    .B1(_11211_),
    .Y(_00009_));
 sky130_fd_sc_hd__mux2_1 _18533_ (.A0(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .S(_08277_),
    .X(_00010_));
 sky130_fd_sc_hd__mux2_1 _18534_ (.A0(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .S(_08277_),
    .X(_00011_));
 sky130_fd_sc_hd__nand2_1 _18535_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .B(_10951_),
    .Y(_11212_));
 sky130_fd_sc_hd__o21ai_0 _18536_ (.A1(_08502_),
    .A2(_10951_),
    .B1(_11212_),
    .Y(_00012_));
 sky130_fd_sc_hd__nand2_1 _18537_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .B(_10815_),
    .Y(_11213_));
 sky130_fd_sc_hd__nand2_8 _18538_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .B(_10951_),
    .Y(_11214_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_775 ();
 sky130_fd_sc_hd__nand2_1 _18541_ (.A(_11213_),
    .B(_11214_),
    .Y(_00013_));
 sky130_fd_sc_hd__nand2_1 _18542_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .B(_10815_),
    .Y(_11217_));
 sky130_fd_sc_hd__nand2_1 _18543_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_valid ),
    .B(_10951_),
    .Y(_11218_));
 sky130_fd_sc_hd__nand2_1 _18544_ (.A(_11217_),
    .B(_11218_),
    .Y(_00014_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_772 ();
 sky130_fd_sc_hd__nor2_1 _18548_ (.A(net819),
    .B(_10854_),
    .Y(_11222_));
 sky130_fd_sc_hd__nand2_1 _18549_ (.A(net927),
    .B(_11222_),
    .Y(_11223_));
 sky130_fd_sc_hd__nor2_1 _18550_ (.A(net1138),
    .B(_11223_),
    .Y(_11224_));
 sky130_fd_sc_hd__nand3_4 _18551_ (.A(_10875_),
    .B(_10925_),
    .C(_11224_),
    .Y(_11225_));
 sky130_fd_sc_hd__nor3b_2 _18552_ (.A(_10876_),
    .B(net1145),
    .C_N(net1136),
    .Y(_11226_));
 sky130_fd_sc_hd__a31oi_1 _18553_ (.A1(\cs_registers_i.debug_mode_i ),
    .A2(_10879_),
    .A3(_11226_),
    .B1(_10880_),
    .Y(_11227_));
 sky130_fd_sc_hd__o21ai_0 _18554_ (.A1(net974),
    .A2(_11227_),
    .B1(_10882_),
    .Y(_11228_));
 sky130_fd_sc_hd__nor2_1 _18555_ (.A(net784),
    .B(_11223_),
    .Y(_11229_));
 sky130_fd_sc_hd__nand2_1 _18556_ (.A(_11228_),
    .B(_11229_),
    .Y(_11230_));
 sky130_fd_sc_hd__nand2_8 _18557_ (.A(_10903_),
    .B(_10899_),
    .Y(_11231_));
 sky130_fd_sc_hd__nand2_1 _18558_ (.A(_10896_),
    .B(_11231_),
    .Y(_11232_));
 sky130_fd_sc_hd__a41oi_1 _18559_ (.A1(_10888_),
    .A2(_11222_),
    .A3(_11226_),
    .A4(_11232_),
    .B1(_10912_),
    .Y(_11233_));
 sky130_fd_sc_hd__nand2_1 _18560_ (.A(_10898_),
    .B(_11233_),
    .Y(_11234_));
 sky130_fd_sc_hd__nor2_1 _18561_ (.A(_10876_),
    .B(_10884_),
    .Y(_11235_));
 sky130_fd_sc_hd__nor2_1 _18562_ (.A(net974),
    .B(_10854_),
    .Y(_11236_));
 sky130_fd_sc_hd__nand4_1 _18563_ (.A(_10852_),
    .B(_10856_),
    .C(_11235_),
    .D(_11236_),
    .Y(_11237_));
 sky130_fd_sc_hd__nor3_4 _18564_ (.A(_10868_),
    .B(_10893_),
    .C(_11237_),
    .Y(_11238_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_771 ();
 sky130_fd_sc_hd__nor4_1 _18566_ (.A(_10909_),
    .B(_10918_),
    .C(_11234_),
    .D(_11238_),
    .Y(_11240_));
 sky130_fd_sc_hd__a31oi_1 _18567_ (.A1(_10852_),
    .A2(_10856_),
    .A3(_10858_),
    .B1(_10863_),
    .Y(_11241_));
 sky130_fd_sc_hd__nand2_1 _18568_ (.A(_10858_),
    .B(_11241_),
    .Y(_11242_));
 sky130_fd_sc_hd__a41oi_4 _18569_ (.A1(_10926_),
    .A2(_11225_),
    .A3(_11230_),
    .A4(_11240_),
    .B1(_11242_),
    .Y(_11243_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_770 ();
 sky130_fd_sc_hd__nand2_1 _18571_ (.A(_10907_),
    .B(net271),
    .Y(_11245_));
 sky130_fd_sc_hd__inv_6 _18572_ (.A(_08745_),
    .Y(_11246_));
 sky130_fd_sc_hd__nand3_4 _18573_ (.A(_11246_),
    .B(_11226_),
    .C(_11229_),
    .Y(_11247_));
 sky130_fd_sc_hd__nor2_8 _18574_ (.A(_10896_),
    .B(_11247_),
    .Y(_11248_));
 sky130_fd_sc_hd__a221oi_4 _18575_ (.A1(net62),
    .A2(_11238_),
    .B1(_11248_),
    .B2(\cs_registers_i.dcsr_q[0] ),
    .C1(_10918_),
    .Y(_11249_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_769 ();
 sky130_fd_sc_hd__nand3_4 _18577_ (.A(_10902_),
    .B(net725),
    .C(_10899_),
    .Y(_11251_));
 sky130_fd_sc_hd__nor2_8 _18578_ (.A(_11251_),
    .B(_11247_),
    .Y(_11252_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_768 ();
 sky130_fd_sc_hd__a22oi_1 _18580_ (.A1(\cs_registers_i.mcountinhibit[0] ),
    .A2(_10907_),
    .B1(_11252_),
    .B2(\cs_registers_i.dscratch0_q[0] ),
    .Y(_11254_));
 sky130_fd_sc_hd__nor2_8 _18581_ (.A(_10896_),
    .B(_10889_),
    .Y(_11255_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_765 ();
 sky130_fd_sc_hd__nand3_4 _18585_ (.A(net641),
    .B(net723),
    .C(_10899_),
    .Y(_11259_));
 sky130_fd_sc_hd__nor2_8 _18586_ (.A(_11247_),
    .B(_11259_),
    .Y(_11260_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_764 ();
 sky130_fd_sc_hd__a22oi_1 _18588_ (.A1(\cs_registers_i.mscratch_q[0] ),
    .A2(_11255_),
    .B1(_11260_),
    .B2(\cs_registers_i.dscratch1_q[0] ),
    .Y(_11262_));
 sky130_fd_sc_hd__nand3_1 _18589_ (.A(_11249_),
    .B(_11254_),
    .C(_11262_),
    .Y(_11263_));
 sky130_fd_sc_hd__nand2_8 _18590_ (.A(_10869_),
    .B(_10906_),
    .Y(_11264_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_763 ();
 sky130_fd_sc_hd__nand3_4 _18592_ (.A(_10902_),
    .B(net726),
    .C(_10899_),
    .Y(_11266_));
 sky130_fd_sc_hd__nor2_8 _18593_ (.A(_11246_),
    .B(_11266_),
    .Y(_11267_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_762 ();
 sky130_fd_sc_hd__a22oi_2 _18595_ (.A1(\cs_registers_i.mcycle_counter_i.counter[0] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][0] ),
    .Y(_11269_));
 sky130_fd_sc_hd__nor2_8 _18596_ (.A(_10889_),
    .B(_11259_),
    .Y(_11270_));
 sky130_fd_sc_hd__nor2_4 _18597_ (.A(_10889_),
    .B(_11251_),
    .Y(_11271_));
 sky130_fd_sc_hd__nor2_8 _18598_ (.A(_10889_),
    .B(_11231_),
    .Y(_11272_));
 sky130_fd_sc_hd__a222oi_1 _18599_ (.A1(\cs_registers_i.mtval_q[0] ),
    .A2(_11270_),
    .B1(_11271_),
    .B2(\cs_registers_i.mcause_q[0] ),
    .C1(\cs_registers_i.csr_mepc_o[0] ),
    .C2(_11272_),
    .Y(_11273_));
 sky130_fd_sc_hd__o21ai_1 _18600_ (.A1(_10926_),
    .A2(_11269_),
    .B1(_11273_),
    .Y(_11274_));
 sky130_fd_sc_hd__a22oi_1 _18601_ (.A1(\cs_registers_i.mcycle_counter_i.counter[32] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][32] ),
    .Y(_11275_));
 sky130_fd_sc_hd__nor2_2 _18602_ (.A(_11225_),
    .B(_11275_),
    .Y(_11276_));
 sky130_fd_sc_hd__nor3_4 _18603_ (.A(_11263_),
    .B(_11274_),
    .C(_11276_),
    .Y(_11277_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_761 ();
 sky130_fd_sc_hd__nand2_1 _18605_ (.A(net731),
    .B(_11146_),
    .Y(_11279_));
 sky130_fd_sc_hd__o22a_4 _18606_ (.A1(net732),
    .A2(_11151_),
    .B1(_11277_),
    .B2(_11279_),
    .X(_11280_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_760 ();
 sky130_fd_sc_hd__nand2_1 _18608_ (.A(\cs_registers_i.mcountinhibit[0] ),
    .B(_11245_),
    .Y(_11282_));
 sky130_fd_sc_hd__o21ai_0 _18609_ (.A1(_11245_),
    .A2(_11280_),
    .B1(_11282_),
    .Y(_00015_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_757 ();
 sky130_fd_sc_hd__a22oi_4 _18613_ (.A1(\cs_registers_i.mcycle_counter_i.counter[2] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][2] ),
    .Y(_11286_));
 sky130_fd_sc_hd__a21oi_1 _18614_ (.A1(\cs_registers_i.csr_mepc_o[2] ),
    .A2(_10890_),
    .B1(_10887_),
    .Y(_11287_));
 sky130_fd_sc_hd__o22ai_2 _18615_ (.A1(_10926_),
    .A2(_11286_),
    .B1(_11287_),
    .B2(_11231_),
    .Y(_11288_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_756 ();
 sky130_fd_sc_hd__a22oi_4 _18617_ (.A1(\cs_registers_i.mcycle_counter_i.counter[34] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][34] ),
    .Y(_11290_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_754 ();
 sky130_fd_sc_hd__a222oi_1 _18620_ (.A1(\cs_registers_i.mcountinhibit[2] ),
    .A2(_10907_),
    .B1(_11252_),
    .B2(\cs_registers_i.dscratch0_q[2] ),
    .C1(_11260_),
    .C2(\cs_registers_i.dscratch1_q[2] ),
    .Y(_11293_));
 sky130_fd_sc_hd__o21ai_4 _18621_ (.A1(_11225_),
    .A2(_11290_),
    .B1(_11293_),
    .Y(_11294_));
 sky130_fd_sc_hd__nor2_8 _18622_ (.A(_11231_),
    .B(_11247_),
    .Y(_11295_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_751 ();
 sky130_fd_sc_hd__a222oi_1 _18626_ (.A1(\cs_registers_i.dcsr_q[2] ),
    .A2(_11248_),
    .B1(_11295_),
    .B2(\cs_registers_i.csr_depc_o[2] ),
    .C1(net84),
    .C2(_11238_),
    .Y(_11299_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_749 ();
 sky130_fd_sc_hd__nand2_1 _18629_ (.A(\cs_registers_i.mtval_q[2] ),
    .B(_11270_),
    .Y(_11302_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_747 ();
 sky130_fd_sc_hd__a22oi_1 _18632_ (.A1(\cs_registers_i.mscratch_q[2] ),
    .A2(_11255_),
    .B1(_11271_),
    .B2(\cs_registers_i.mcause_q[2] ),
    .Y(_11305_));
 sky130_fd_sc_hd__nand3_2 _18633_ (.A(_11299_),
    .B(_11302_),
    .C(_11305_),
    .Y(_11306_));
 sky130_fd_sc_hd__nor3_4 _18634_ (.A(_11288_),
    .B(_11294_),
    .C(_11306_),
    .Y(_11307_));
 sky130_fd_sc_hd__nand2_1 _18635_ (.A(_08850_),
    .B(_11146_),
    .Y(_11308_));
 sky130_fd_sc_hd__o22a_4 _18636_ (.A1(_08850_),
    .A2(_11151_),
    .B1(_11307_),
    .B2(_11308_),
    .X(_11309_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_746 ();
 sky130_fd_sc_hd__nand2_1 _18638_ (.A(\cs_registers_i.mcountinhibit[2] ),
    .B(_11245_),
    .Y(_11311_));
 sky130_fd_sc_hd__o21ai_0 _18639_ (.A1(_11245_),
    .A2(_11309_),
    .B1(_11311_),
    .Y(_00016_));
 sky130_fd_sc_hd__inv_1 _18640_ (.A(_10864_),
    .Y(_11312_));
 sky130_fd_sc_hd__nand2_8 _18641_ (.A(_10858_),
    .B(_11312_),
    .Y(_11313_));
 sky130_fd_sc_hd__nor2_2 _18642_ (.A(_10930_),
    .B(_11313_),
    .Y(_11314_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_745 ();
 sky130_fd_sc_hd__nand3_4 _18644_ (.A(_10929_),
    .B(_11314_),
    .C(_11264_),
    .Y(_11316_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_742 ();
 sky130_fd_sc_hd__nand3b_4 _18648_ (.A_N(_11313_),
    .B(_11264_),
    .C(_10929_),
    .Y(_11320_));
 sky130_fd_sc_hd__nand2_1 _18649_ (.A(\cs_registers_i.mcountinhibit[0] ),
    .B(_11320_),
    .Y(_11321_));
 sky130_fd_sc_hd__o21a_4 _18650_ (.A1(_10928_),
    .A2(_11316_),
    .B1(_11321_),
    .X(_11322_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_741 ();
 sky130_fd_sc_hd__o21ai_0 _18652_ (.A1(_11280_),
    .A2(_11316_),
    .B1(_11322_),
    .Y(_11324_));
 sky130_fd_sc_hd__o21ai_4 _18653_ (.A1(_10914_),
    .A2(_10927_),
    .B1(_10925_),
    .Y(_11325_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_739 ();
 sky130_fd_sc_hd__nor3b_4 _18656_ (.A(_11325_),
    .B(_11313_),
    .C_N(_11264_),
    .Y(_11328_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_738 ();
 sky130_fd_sc_hd__o21ai_4 _18658_ (.A1(_10928_),
    .A2(_11316_),
    .B1(_11321_),
    .Y(_11330_));
 sky130_fd_sc_hd__a211oi_1 _18659_ (.A1(_11280_),
    .A2(_11328_),
    .B1(_11330_),
    .C1(\cs_registers_i.mcycle_counter_i.counter[0] ),
    .Y(_11331_));
 sky130_fd_sc_hd__a21o_1 _18660_ (.A1(\cs_registers_i.mcycle_counter_i.counter[0] ),
    .A2(_11324_),
    .B1(_11331_),
    .X(_00017_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_737 ();
 sky130_fd_sc_hd__inv_1 _18662_ (.A(\cs_registers_i.mcycle_counter_i.counter[3] ),
    .Y(_11333_));
 sky130_fd_sc_hd__nand3_4 _18663_ (.A(\cs_registers_i.mcycle_counter_i.counter[0] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[1] ),
    .C(\cs_registers_i.mcycle_counter_i.counter[2] ),
    .Y(_11334_));
 sky130_fd_sc_hd__nor2_8 _18664_ (.A(_11333_),
    .B(_11334_),
    .Y(_11335_));
 sky130_fd_sc_hd__nand2_8 _18665_ (.A(_11320_),
    .B(_11335_),
    .Y(_11336_));
 sky130_fd_sc_hd__and3_1 _18666_ (.A(\cs_registers_i.mcycle_counter_i.counter[4] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[5] ),
    .C(\cs_registers_i.mcycle_counter_i.counter[6] ),
    .X(_11337_));
 sky130_fd_sc_hd__and3_1 _18667_ (.A(\cs_registers_i.mcycle_counter_i.counter[7] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[8] ),
    .C(_11337_),
    .X(_11338_));
 sky130_fd_sc_hd__nand3_1 _18668_ (.A(\cs_registers_i.mcycle_counter_i.counter[9] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[10] ),
    .C(_11338_),
    .Y(_11339_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_732 ();
 sky130_fd_sc_hd__a22oi_2 _18674_ (.A1(\cs_registers_i.mcycle_counter_i.counter[42] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][42] ),
    .Y(_11345_));
 sky130_fd_sc_hd__a22oi_2 _18675_ (.A1(\cs_registers_i.mcycle_counter_i.counter[10] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][10] ),
    .Y(_11346_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_731 ();
 sky130_fd_sc_hd__a222oi_1 _18677_ (.A1(\cs_registers_i.csr_mtvec_o[10] ),
    .A2(_10918_),
    .B1(_11252_),
    .B2(\cs_registers_i.dscratch0_q[10] ),
    .C1(\cs_registers_i.dscratch1_q[10] ),
    .C2(_11260_),
    .Y(_11348_));
 sky130_fd_sc_hd__o221ai_4 _18678_ (.A1(_11225_),
    .A2(_11345_),
    .B1(_11346_),
    .B2(_10926_),
    .C1(net1019),
    .Y(_11349_));
 sky130_fd_sc_hd__a221o_1 _18679_ (.A1(net63),
    .A2(_11238_),
    .B1(_11295_),
    .B2(\cs_registers_i.csr_depc_o[10] ),
    .C1(_10907_),
    .X(_11350_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_729 ();
 sky130_fd_sc_hd__a22o_1 _18682_ (.A1(\cs_registers_i.csr_mepc_o[10] ),
    .A2(_11272_),
    .B1(_11270_),
    .B2(\cs_registers_i.mtval_q[10] ),
    .X(_11353_));
 sky130_fd_sc_hd__a2111oi_4 _18683_ (.A1(\cs_registers_i.mscratch_q[10] ),
    .A2(_11255_),
    .B1(_11349_),
    .C1(_11350_),
    .D1(_11353_),
    .Y(_11354_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_728 ();
 sky130_fd_sc_hd__nand2_1 _18685_ (.A(_09385_),
    .B(_11148_),
    .Y(_11356_));
 sky130_fd_sc_hd__o31ai_4 _18686_ (.A1(_09385_),
    .A2(_11150_),
    .A3(_11354_),
    .B1(_11356_),
    .Y(_11357_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_726 ();
 sky130_fd_sc_hd__o22ai_1 _18689_ (.A1(_11336_),
    .A2(_11339_),
    .B1(_11357_),
    .B2(_11316_),
    .Y(_11360_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_722 ();
 sky130_fd_sc_hd__nand3_1 _18694_ (.A(\cs_registers_i.mcycle_counter_i.counter[9] ),
    .B(_11335_),
    .C(_11338_),
    .Y(_11365_));
 sky130_fd_sc_hd__nand2_1 _18695_ (.A(_11320_),
    .B(_11365_),
    .Y(_11366_));
 sky130_fd_sc_hd__a21oi_1 _18696_ (.A1(_11322_),
    .A2(_11366_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[10] ),
    .Y(_11367_));
 sky130_fd_sc_hd__a21oi_1 _18697_ (.A1(_11322_),
    .A2(_11360_),
    .B1(_11367_),
    .Y(_00018_));
 sky130_fd_sc_hd__a222oi_1 _18698_ (.A1(\cs_registers_i.csr_mtvec_o[11] ),
    .A2(_10918_),
    .B1(_11252_),
    .B2(\cs_registers_i.dscratch0_q[11] ),
    .C1(\cs_registers_i.dscratch1_q[11] ),
    .C2(_11260_),
    .Y(_11368_));
 sky130_fd_sc_hd__a21oi_1 _18699_ (.A1(net64),
    .A2(_11238_),
    .B1(_10907_),
    .Y(_11369_));
 sky130_fd_sc_hd__a22oi_1 _18700_ (.A1(\cs_registers_i.dcsr_q[11] ),
    .A2(_11248_),
    .B1(_11295_),
    .B2(\cs_registers_i.csr_depc_o[11] ),
    .Y(_11370_));
 sky130_fd_sc_hd__inv_1 _18701_ (.A(_10886_),
    .Y(_11371_));
 sky130_fd_sc_hd__nand2_4 _18702_ (.A(_10880_),
    .B(_11371_),
    .Y(_11372_));
 sky130_fd_sc_hd__nor2_8 _18703_ (.A(_10893_),
    .B(_11372_),
    .Y(_11373_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_721 ();
 sky130_fd_sc_hd__nor2_8 _18705_ (.A(_10896_),
    .B(_11372_),
    .Y(_11375_));
 sky130_fd_sc_hd__a22oi_1 _18706_ (.A1(\cs_registers_i.mie_q[15] ),
    .A2(_11373_),
    .B1(_11375_),
    .B2(\cs_registers_i.mstack_d[0] ),
    .Y(_11376_));
 sky130_fd_sc_hd__nand4_1 _18707_ (.A(_11368_),
    .B(_11369_),
    .C(_11370_),
    .D(_11376_),
    .Y(_11377_));
 sky130_fd_sc_hd__a22oi_2 _18708_ (.A1(\cs_registers_i.mcycle_counter_i.counter[11] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][11] ),
    .Y(_11378_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_719 ();
 sky130_fd_sc_hd__a22oi_2 _18711_ (.A1(\cs_registers_i.mcycle_counter_i.counter[43] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][43] ),
    .Y(_11381_));
 sky130_fd_sc_hd__o22ai_4 _18712_ (.A1(_10926_),
    .A2(_11378_),
    .B1(_11381_),
    .B2(_11225_),
    .Y(_11382_));
 sky130_fd_sc_hd__nor2_1 _18713_ (.A(_11377_),
    .B(_11382_),
    .Y(_11383_));
 sky130_fd_sc_hd__nor2_8 _18714_ (.A(_10893_),
    .B(_10889_),
    .Y(_11384_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_718 ();
 sky130_fd_sc_hd__a22oi_2 _18716_ (.A1(\cs_registers_i.mtval_q[11] ),
    .A2(_11270_),
    .B1(_11384_),
    .B2(net129),
    .Y(_11386_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_717 ();
 sky130_fd_sc_hd__a22oi_2 _18718_ (.A1(\cs_registers_i.mscratch_q[11] ),
    .A2(_11255_),
    .B1(_11272_),
    .B2(\cs_registers_i.csr_mepc_o[11] ),
    .Y(_11388_));
 sky130_fd_sc_hd__nand3_4 _18719_ (.A(_11383_),
    .B(_11386_),
    .C(_11388_),
    .Y(_11389_));
 sky130_fd_sc_hd__nor2_1 _18720_ (.A(net877),
    .B(_11151_),
    .Y(_11390_));
 sky130_fd_sc_hd__a31o_4 _18721_ (.A1(net877),
    .A2(_11146_),
    .A3(_11389_),
    .B1(_11390_),
    .X(_11391_));
 sky130_fd_sc_hd__nand4_4 _18722_ (.A(\cs_registers_i.mcycle_counter_i.counter[0] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[1] ),
    .C(\cs_registers_i.mcycle_counter_i.counter[2] ),
    .D(\cs_registers_i.mcycle_counter_i.counter[3] ),
    .Y(_11392_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_716 ();
 sky130_fd_sc_hd__nor2_4 _18724_ (.A(net273),
    .B(_11392_),
    .Y(_11394_));
 sky130_fd_sc_hd__inv_1 _18725_ (.A(\cs_registers_i.mcycle_counter_i.counter[11] ),
    .Y(_11395_));
 sky130_fd_sc_hd__nor2_2 _18726_ (.A(_11395_),
    .B(_11339_),
    .Y(_11396_));
 sky130_fd_sc_hd__nand2_1 _18727_ (.A(_11394_),
    .B(_11396_),
    .Y(_11397_));
 sky130_fd_sc_hd__o21ai_0 _18728_ (.A1(_11316_),
    .A2(_11391_),
    .B1(_11397_),
    .Y(_11398_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_715 ();
 sky130_fd_sc_hd__o21ai_0 _18730_ (.A1(_11392_),
    .A2(_11339_),
    .B1(_11316_),
    .Y(_11400_));
 sky130_fd_sc_hd__a21oi_1 _18731_ (.A1(_11322_),
    .A2(_11400_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[11] ),
    .Y(_11401_));
 sky130_fd_sc_hd__a21oi_1 _18732_ (.A1(_11322_),
    .A2(_11398_),
    .B1(_11401_),
    .Y(_00019_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_714 ();
 sky130_fd_sc_hd__nand2_1 _18734_ (.A(\cs_registers_i.mcycle_counter_i.counter[12] ),
    .B(_11396_),
    .Y(_11403_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_712 ();
 sky130_fd_sc_hd__a22oi_2 _18737_ (.A1(\cs_registers_i.mcycle_counter_i.counter[12] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][12] ),
    .Y(_11406_));
 sky130_fd_sc_hd__a22oi_2 _18738_ (.A1(\cs_registers_i.mcycle_counter_i.counter[44] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][44] ),
    .Y(_11407_));
 sky130_fd_sc_hd__nand3_4 _18739_ (.A(_11246_),
    .B(_10877_),
    .C(_10871_),
    .Y(_11408_));
 sky130_fd_sc_hd__nor2_8 _18740_ (.A(_11266_),
    .B(_11408_),
    .Y(_11409_));
 sky130_fd_sc_hd__nor2_4 _18741_ (.A(_10896_),
    .B(_11408_),
    .Y(_11410_));
 sky130_fd_sc_hd__o22ai_4 _18742_ (.A1(_10905_),
    .A2(_10906_),
    .B1(_11231_),
    .B2(_11372_),
    .Y(_11411_));
 sky130_fd_sc_hd__a221o_1 _18743_ (.A1(\cs_registers_i.dscratch0_q[12] ),
    .A2(_11409_),
    .B1(_11410_),
    .B2(\cs_registers_i.dcsr_q[12] ),
    .C1(_11411_),
    .X(_11412_));
 sky130_fd_sc_hd__a221oi_4 _18744_ (.A1(\cs_registers_i.csr_mtvec_o[12] ),
    .A2(_10918_),
    .B1(_11375_),
    .B2(\cs_registers_i.mstack_d[1] ),
    .C1(_11412_),
    .Y(_11413_));
 sky130_fd_sc_hd__o221ai_4 _18745_ (.A1(_10926_),
    .A2(_11406_),
    .B1(_11407_),
    .B2(_10928_),
    .C1(_11413_),
    .Y(_11414_));
 sky130_fd_sc_hd__nand3_4 _18746_ (.A(net642),
    .B(net727),
    .C(_10899_),
    .Y(_11415_));
 sky130_fd_sc_hd__nor2_8 _18747_ (.A(_11408_),
    .B(_11415_),
    .Y(_11416_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_711 ();
 sky130_fd_sc_hd__nor2_8 _18749_ (.A(_11231_),
    .B(_11408_),
    .Y(_11418_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_709 ();
 sky130_fd_sc_hd__a222oi_1 _18752_ (.A1(\cs_registers_i.dscratch1_q[12] ),
    .A2(_11416_),
    .B1(_11418_),
    .B2(\cs_registers_i.csr_depc_o[12] ),
    .C1(net65),
    .C2(net1231),
    .Y(_11421_));
 sky130_fd_sc_hd__nor2_8 _18753_ (.A(_10889_),
    .B(_11415_),
    .Y(_11422_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_708 ();
 sky130_fd_sc_hd__a22oi_1 _18755_ (.A1(\cs_registers_i.mtval_q[12] ),
    .A2(_11422_),
    .B1(_11272_),
    .B2(\cs_registers_i.csr_mepc_o[12] ),
    .Y(_11424_));
 sky130_fd_sc_hd__nand2_1 _18756_ (.A(_11421_),
    .B(_11424_),
    .Y(_11425_));
 sky130_fd_sc_hd__a211o_2 _18757_ (.A1(\cs_registers_i.mscratch_q[12] ),
    .A2(_11255_),
    .B1(_11414_),
    .C1(_11425_),
    .X(_11426_));
 sky130_fd_sc_hd__a21oi_1 _18758_ (.A1(_11146_),
    .A2(_11426_),
    .B1(_09562_),
    .Y(_11427_));
 sky130_fd_sc_hd__a21o_4 _18759_ (.A1(_09562_),
    .A2(_11151_),
    .B1(_11427_),
    .X(_11428_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_707 ();
 sky130_fd_sc_hd__nand2_1 _18761_ (.A(net273),
    .B(_11428_),
    .Y(_11430_));
 sky130_fd_sc_hd__o21ai_0 _18762_ (.A1(_11336_),
    .A2(_11403_),
    .B1(_11430_),
    .Y(_11431_));
 sky130_fd_sc_hd__nand2_1 _18763_ (.A(_11335_),
    .B(_11396_),
    .Y(_11432_));
 sky130_fd_sc_hd__nand2_1 _18764_ (.A(_11320_),
    .B(_11432_),
    .Y(_11433_));
 sky130_fd_sc_hd__a21oi_1 _18765_ (.A1(_11322_),
    .A2(_11433_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[12] ),
    .Y(_11434_));
 sky130_fd_sc_hd__a21oi_1 _18766_ (.A1(_11322_),
    .A2(_11431_),
    .B1(_11434_),
    .Y(_00020_));
 sky130_fd_sc_hd__nand3_1 _18767_ (.A(\cs_registers_i.mcycle_counter_i.counter[12] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[13] ),
    .C(_11396_),
    .Y(_11435_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_705 ();
 sky130_fd_sc_hd__a22oi_4 _18770_ (.A1(\cs_registers_i.mcycle_counter_i.counter[45] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][45] ),
    .Y(_11438_));
 sky130_fd_sc_hd__a22oi_4 _18771_ (.A1(\cs_registers_i.mcycle_counter_i.counter[13] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][13] ),
    .Y(_11439_));
 sky130_fd_sc_hd__a222oi_1 _18772_ (.A1(net66),
    .A2(net1231),
    .B1(_10918_),
    .B2(\cs_registers_i.csr_mtvec_o[13] ),
    .C1(\cs_registers_i.csr_depc_o[13] ),
    .C2(_11418_),
    .Y(_11440_));
 sky130_fd_sc_hd__a22oi_1 _18773_ (.A1(\cs_registers_i.dcsr_q[13] ),
    .A2(_11410_),
    .B1(_11416_),
    .B2(\cs_registers_i.dscratch1_q[13] ),
    .Y(_11441_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_704 ();
 sky130_fd_sc_hd__a21oi_1 _18775_ (.A1(\cs_registers_i.dscratch0_q[13] ),
    .A2(_11409_),
    .B1(_10907_),
    .Y(_11443_));
 sky130_fd_sc_hd__o2111a_1 _18776_ (.A1(_10926_),
    .A2(_11439_),
    .B1(_11440_),
    .C1(_11441_),
    .D1(_11443_),
    .X(_11444_));
 sky130_fd_sc_hd__a222oi_1 _18777_ (.A1(\cs_registers_i.mtval_q[13] ),
    .A2(_11422_),
    .B1(_11255_),
    .B2(\cs_registers_i.mscratch_q[13] ),
    .C1(_11272_),
    .C2(\cs_registers_i.csr_mepc_o[13] ),
    .Y(_11445_));
 sky130_fd_sc_hd__o211ai_4 _18778_ (.A1(_10928_),
    .A2(_11438_),
    .B1(_11444_),
    .C1(_11445_),
    .Y(_11446_));
 sky130_fd_sc_hd__a21oi_1 _18779_ (.A1(_11146_),
    .A2(_11446_),
    .B1(net737),
    .Y(_11447_));
 sky130_fd_sc_hd__a21o_4 _18780_ (.A1(net737),
    .A2(_11151_),
    .B1(_11447_),
    .X(_11448_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_703 ();
 sky130_fd_sc_hd__nand2_1 _18782_ (.A(net273),
    .B(_11448_),
    .Y(_11450_));
 sky130_fd_sc_hd__o21ai_0 _18783_ (.A1(_11336_),
    .A2(_11435_),
    .B1(_11450_),
    .Y(_11451_));
 sky130_fd_sc_hd__o21ai_0 _18784_ (.A1(_11392_),
    .A2(_11403_),
    .B1(_11316_),
    .Y(_11452_));
 sky130_fd_sc_hd__a21oi_1 _18785_ (.A1(_11322_),
    .A2(_11452_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[13] ),
    .Y(_11453_));
 sky130_fd_sc_hd__a21oi_1 _18786_ (.A1(_11322_),
    .A2(_11451_),
    .B1(_11453_),
    .Y(_00021_));
 sky130_fd_sc_hd__nand4_4 _18787_ (.A(\cs_registers_i.mcycle_counter_i.counter[12] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[13] ),
    .C(\cs_registers_i.mcycle_counter_i.counter[14] ),
    .D(_11396_),
    .Y(_11454_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_702 ();
 sky130_fd_sc_hd__a22oi_4 _18789_ (.A1(\cs_registers_i.mcycle_counter_i.counter[46] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][46] ),
    .Y(_11456_));
 sky130_fd_sc_hd__a22oi_4 _18790_ (.A1(\cs_registers_i.mcycle_counter_i.counter[14] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][14] ),
    .Y(_11457_));
 sky130_fd_sc_hd__a222oi_1 _18791_ (.A1(\cs_registers_i.dscratch0_q[14] ),
    .A2(_11409_),
    .B1(_11418_),
    .B2(\cs_registers_i.csr_depc_o[14] ),
    .C1(net67),
    .C2(net1231),
    .Y(_11458_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_701 ();
 sky130_fd_sc_hd__a221oi_4 _18793_ (.A1(\cs_registers_i.csr_mtvec_o[14] ),
    .A2(_10918_),
    .B1(_11416_),
    .B2(\cs_registers_i.dscratch1_q[14] ),
    .C1(_10907_),
    .Y(_11460_));
 sky130_fd_sc_hd__o211a_1 _18794_ (.A1(_10926_),
    .A2(_11457_),
    .B1(_11458_),
    .C1(_11460_),
    .X(_11461_));
 sky130_fd_sc_hd__a222oi_1 _18795_ (.A1(\cs_registers_i.mtval_q[14] ),
    .A2(_11422_),
    .B1(_11255_),
    .B2(\cs_registers_i.mscratch_q[14] ),
    .C1(_11272_),
    .C2(\cs_registers_i.csr_mepc_o[14] ),
    .Y(_11462_));
 sky130_fd_sc_hd__o211ai_4 _18796_ (.A1(_10928_),
    .A2(_11456_),
    .B1(_11461_),
    .C1(_11462_),
    .Y(_11463_));
 sky130_fd_sc_hd__a21oi_1 _18797_ (.A1(_11146_),
    .A2(_11463_),
    .B1(_09640_),
    .Y(_11464_));
 sky130_fd_sc_hd__a21o_4 _18798_ (.A1(_09640_),
    .A2(_11151_),
    .B1(_11464_),
    .X(_11465_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_700 ();
 sky130_fd_sc_hd__nand2_1 _18800_ (.A(net273),
    .B(_11465_),
    .Y(_11467_));
 sky130_fd_sc_hd__o21ai_0 _18801_ (.A1(_11336_),
    .A2(_11454_),
    .B1(_11467_),
    .Y(_11468_));
 sky130_fd_sc_hd__o21ai_0 _18802_ (.A1(_11392_),
    .A2(_11435_),
    .B1(_11316_),
    .Y(_11469_));
 sky130_fd_sc_hd__a21oi_1 _18803_ (.A1(_11322_),
    .A2(_11469_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[14] ),
    .Y(_11470_));
 sky130_fd_sc_hd__a21oi_1 _18804_ (.A1(_11322_),
    .A2(_11468_),
    .B1(_11470_),
    .Y(_00022_));
 sky130_fd_sc_hd__inv_1 _18805_ (.A(\cs_registers_i.mcycle_counter_i.counter[15] ),
    .Y(_11471_));
 sky130_fd_sc_hd__and3_4 _18806_ (.A(_10929_),
    .B(_11314_),
    .C(_11264_),
    .X(_11472_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_698 ();
 sky130_fd_sc_hd__nor2_1 _18809_ (.A(_11392_),
    .B(_11454_),
    .Y(_11475_));
 sky130_fd_sc_hd__o21ai_0 _18810_ (.A1(_11472_),
    .A2(_11475_),
    .B1(_11322_),
    .Y(_11476_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_696 ();
 sky130_fd_sc_hd__a22oi_4 _18813_ (.A1(\cs_registers_i.mcycle_counter_i.counter[47] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][47] ),
    .Y(_11479_));
 sky130_fd_sc_hd__a22oi_4 _18814_ (.A1(\cs_registers_i.mcycle_counter_i.counter[15] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][15] ),
    .Y(_11480_));
 sky130_fd_sc_hd__a222oi_1 _18815_ (.A1(net68),
    .A2(net1231),
    .B1(_10918_),
    .B2(\cs_registers_i.csr_mtvec_o[15] ),
    .C1(\cs_registers_i.csr_depc_o[15] ),
    .C2(_11418_),
    .Y(_11481_));
 sky130_fd_sc_hd__a22oi_2 _18816_ (.A1(\cs_registers_i.dcsr_q[15] ),
    .A2(_11410_),
    .B1(_11416_),
    .B2(\cs_registers_i.dscratch1_q[15] ),
    .Y(_11482_));
 sky130_fd_sc_hd__a21oi_1 _18817_ (.A1(\cs_registers_i.dscratch0_q[15] ),
    .A2(_11409_),
    .B1(_10907_),
    .Y(_11483_));
 sky130_fd_sc_hd__o2111a_1 _18818_ (.A1(_10926_),
    .A2(_11480_),
    .B1(_11481_),
    .C1(_11482_),
    .D1(_11483_),
    .X(_11484_));
 sky130_fd_sc_hd__a222oi_1 _18819_ (.A1(\cs_registers_i.mtval_q[15] ),
    .A2(_11422_),
    .B1(_11255_),
    .B2(\cs_registers_i.mscratch_q[15] ),
    .C1(_11272_),
    .C2(\cs_registers_i.csr_mepc_o[15] ),
    .Y(_11485_));
 sky130_fd_sc_hd__o211ai_4 _18820_ (.A1(_10928_),
    .A2(_11479_),
    .B1(_11484_),
    .C1(_11485_),
    .Y(_11486_));
 sky130_fd_sc_hd__a21oi_1 _18821_ (.A1(_11146_),
    .A2(_11486_),
    .B1(_09679_),
    .Y(_11487_));
 sky130_fd_sc_hd__a21o_4 _18822_ (.A1(_09679_),
    .A2(_11151_),
    .B1(_11487_),
    .X(_11488_));
 sky130_fd_sc_hd__nand2_1 _18823_ (.A(net273),
    .B(_11488_),
    .Y(_11489_));
 sky130_fd_sc_hd__o31a_1 _18824_ (.A1(_11471_),
    .A2(_11336_),
    .A3(_11454_),
    .B1(_11489_),
    .X(_11490_));
 sky130_fd_sc_hd__nor2_1 _18825_ (.A(_11330_),
    .B(_11490_),
    .Y(_11491_));
 sky130_fd_sc_hd__a21oi_1 _18826_ (.A1(_11471_),
    .A2(_11476_),
    .B1(_11491_),
    .Y(_00023_));
 sky130_fd_sc_hd__and3_1 _18827_ (.A(\cs_registers_i.mcycle_counter_i.counter[15] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[16] ),
    .C(_11475_),
    .X(_11492_));
 sky130_fd_sc_hd__a221oi_2 _18828_ (.A1(net69),
    .A2(net274),
    .B1(_11295_),
    .B2(\cs_registers_i.csr_depc_o[16] ),
    .C1(_10907_),
    .Y(_11493_));
 sky130_fd_sc_hd__nand2_1 _18829_ (.A(\cs_registers_i.mtval_q[16] ),
    .B(_11270_),
    .Y(_11494_));
 sky130_fd_sc_hd__a22oi_1 _18830_ (.A1(\cs_registers_i.csr_mtvec_o[16] ),
    .A2(_10918_),
    .B1(_11252_),
    .B2(\cs_registers_i.dscratch0_q[16] ),
    .Y(_11495_));
 sky130_fd_sc_hd__a22oi_1 _18831_ (.A1(\cs_registers_i.dscratch1_q[16] ),
    .A2(_11260_),
    .B1(_11373_),
    .B2(\cs_registers_i.mie_q[0] ),
    .Y(_11496_));
 sky130_fd_sc_hd__nand4_1 _18832_ (.A(_11493_),
    .B(_11494_),
    .C(_11495_),
    .D(_11496_),
    .Y(_11497_));
 sky130_fd_sc_hd__a22oi_4 _18833_ (.A1(\cs_registers_i.mcycle_counter_i.counter[16] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][16] ),
    .Y(_11498_));
 sky130_fd_sc_hd__a222oi_1 _18834_ (.A1(\cs_registers_i.mscratch_q[16] ),
    .A2(_11255_),
    .B1(_11272_),
    .B2(\cs_registers_i.csr_mepc_o[16] ),
    .C1(net130),
    .C2(_11384_),
    .Y(_11499_));
 sky130_fd_sc_hd__o21ai_1 _18835_ (.A1(_10926_),
    .A2(_11498_),
    .B1(_11499_),
    .Y(_11500_));
 sky130_fd_sc_hd__a22oi_1 _18836_ (.A1(\cs_registers_i.mcycle_counter_i.counter[48] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][48] ),
    .Y(_11501_));
 sky130_fd_sc_hd__nor2_2 _18837_ (.A(_11225_),
    .B(_11501_),
    .Y(_11502_));
 sky130_fd_sc_hd__nor3_4 _18838_ (.A(_11497_),
    .B(_11500_),
    .C(_11502_),
    .Y(_11503_));
 sky130_fd_sc_hd__nor3_1 _18839_ (.A(_09825_),
    .B(_11150_),
    .C(_11503_),
    .Y(_11504_));
 sky130_fd_sc_hd__a21oi_4 _18840_ (.A1(_09825_),
    .A2(_11148_),
    .B1(_11504_),
    .Y(_11505_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_695 ();
 sky130_fd_sc_hd__mux2i_1 _18842_ (.A0(_11492_),
    .A1(_11505_),
    .S(net273),
    .Y(_11507_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_694 ();
 sky130_fd_sc_hd__a21oi_1 _18844_ (.A1(\cs_registers_i.mcycle_counter_i.counter[15] ),
    .A2(_11475_),
    .B1(net273),
    .Y(_11509_));
 sky130_fd_sc_hd__nor2_1 _18845_ (.A(_11330_),
    .B(_11509_),
    .Y(_11510_));
 sky130_fd_sc_hd__o22a_1 _18846_ (.A1(_11330_),
    .A2(_11507_),
    .B1(_11510_),
    .B2(\cs_registers_i.mcycle_counter_i.counter[16] ),
    .X(_00024_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_693 ();
 sky130_fd_sc_hd__nand2_1 _18848_ (.A(\cs_registers_i.mcycle_counter_i.counter[17] ),
    .B(_11492_),
    .Y(_11512_));
 sky130_fd_sc_hd__a22oi_2 _18849_ (.A1(\cs_registers_i.mcycle_counter_i.counter[17] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][17] ),
    .Y(_11513_));
 sky130_fd_sc_hd__a22oi_2 _18850_ (.A1(\cs_registers_i.mcycle_counter_i.counter[49] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][49] ),
    .Y(_11514_));
 sky130_fd_sc_hd__o22ai_4 _18851_ (.A1(_10926_),
    .A2(_11513_),
    .B1(_11514_),
    .B2(_10928_),
    .Y(_11515_));
 sky130_fd_sc_hd__a22oi_1 _18852_ (.A1(\cs_registers_i.csr_mtvec_o[17] ),
    .A2(_10918_),
    .B1(_11373_),
    .B2(\cs_registers_i.mie_q[1] ),
    .Y(_11516_));
 sky130_fd_sc_hd__a222oi_1 _18853_ (.A1(\cs_registers_i.dscratch0_q[17] ),
    .A2(_11409_),
    .B1(_11375_),
    .B2(\cs_registers_i.mstatus_q[1] ),
    .C1(net70),
    .C2(net1230),
    .Y(_11517_));
 sky130_fd_sc_hd__a222oi_1 _18854_ (.A1(\cs_registers_i.mscratch_q[17] ),
    .A2(_11255_),
    .B1(_11272_),
    .B2(\cs_registers_i.csr_mepc_o[17] ),
    .C1(net136),
    .C2(_11384_),
    .Y(_11518_));
 sky130_fd_sc_hd__nand3_1 _18855_ (.A(_11516_),
    .B(_11517_),
    .C(_11518_),
    .Y(_11519_));
 sky130_fd_sc_hd__a221o_1 _18856_ (.A1(\cs_registers_i.dscratch1_q[17] ),
    .A2(_11416_),
    .B1(_11418_),
    .B2(\cs_registers_i.csr_depc_o[17] ),
    .C1(_10907_),
    .X(_11520_));
 sky130_fd_sc_hd__a2111oi_4 _18857_ (.A1(\cs_registers_i.mtval_q[17] ),
    .A2(_11422_),
    .B1(_11515_),
    .C1(_11519_),
    .D1(_11520_),
    .Y(_11521_));
 sky130_fd_sc_hd__o21ai_1 _18858_ (.A1(_11150_),
    .A2(_11521_),
    .B1(_09754_),
    .Y(_11522_));
 sky130_fd_sc_hd__o21ai_4 _18859_ (.A1(_09754_),
    .A2(_11148_),
    .B1(_11522_),
    .Y(_11523_));
 sky130_fd_sc_hd__nand2_1 _18860_ (.A(_11472_),
    .B(_11523_),
    .Y(_11524_));
 sky130_fd_sc_hd__o21ai_0 _18861_ (.A1(net273),
    .A2(_11512_),
    .B1(_11524_),
    .Y(_11525_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_692 ();
 sky130_fd_sc_hd__o21ai_0 _18863_ (.A1(net273),
    .A2(_11492_),
    .B1(_11322_),
    .Y(_11527_));
 sky130_fd_sc_hd__inv_1 _18864_ (.A(\cs_registers_i.mcycle_counter_i.counter[17] ),
    .Y(_11528_));
 sky130_fd_sc_hd__a22oi_1 _18865_ (.A1(_11322_),
    .A2(_11525_),
    .B1(_11527_),
    .B2(_11528_),
    .Y(_00025_));
 sky130_fd_sc_hd__nand2_1 _18866_ (.A(_11316_),
    .B(_11512_),
    .Y(_11529_));
 sky130_fd_sc_hd__a21oi_1 _18867_ (.A1(_11322_),
    .A2(_11529_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[18] ),
    .Y(_11530_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_691 ();
 sky130_fd_sc_hd__nand4_4 _18869_ (.A(\cs_registers_i.mcycle_counter_i.counter[15] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[16] ),
    .C(\cs_registers_i.mcycle_counter_i.counter[17] ),
    .D(\cs_registers_i.mcycle_counter_i.counter[18] ),
    .Y(_11532_));
 sky130_fd_sc_hd__nor3_1 _18870_ (.A(_11392_),
    .B(_11454_),
    .C(_11532_),
    .Y(_11533_));
 sky130_fd_sc_hd__nand2_1 _18871_ (.A(_11320_),
    .B(_11533_),
    .Y(_11534_));
 sky130_fd_sc_hd__a22o_1 _18872_ (.A1(\cs_registers_i.mtval_q[18] ),
    .A2(_11422_),
    .B1(_11255_),
    .B2(\cs_registers_i.mscratch_q[18] ),
    .X(_11535_));
 sky130_fd_sc_hd__a22oi_2 _18873_ (.A1(\cs_registers_i.mcycle_counter_i.counter[18] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][18] ),
    .Y(_11536_));
 sky130_fd_sc_hd__a22oi_2 _18874_ (.A1(\cs_registers_i.mcycle_counter_i.counter[50] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][50] ),
    .Y(_11537_));
 sky130_fd_sc_hd__o22ai_4 _18875_ (.A1(_10926_),
    .A2(_11536_),
    .B1(_11537_),
    .B2(_10928_),
    .Y(_11538_));
 sky130_fd_sc_hd__a221oi_2 _18876_ (.A1(net71),
    .A2(net1231),
    .B1(_11418_),
    .B2(\cs_registers_i.csr_depc_o[18] ),
    .C1(_10907_),
    .Y(_11539_));
 sky130_fd_sc_hd__a222oi_1 _18877_ (.A1(\cs_registers_i.dscratch0_q[18] ),
    .A2(_11409_),
    .B1(_11416_),
    .B2(\cs_registers_i.dscratch1_q[18] ),
    .C1(\cs_registers_i.mie_q[2] ),
    .C2(_11373_),
    .Y(_11540_));
 sky130_fd_sc_hd__a22oi_1 _18878_ (.A1(\cs_registers_i.csr_mtvec_o[18] ),
    .A2(_10918_),
    .B1(_11384_),
    .B2(net137),
    .Y(_11541_));
 sky130_fd_sc_hd__nand3_1 _18879_ (.A(_11539_),
    .B(_11540_),
    .C(_11541_),
    .Y(_11542_));
 sky130_fd_sc_hd__a2111oi_4 _18880_ (.A1(\cs_registers_i.csr_mepc_o[18] ),
    .A2(_11272_),
    .B1(_11535_),
    .C1(_11538_),
    .D1(_11542_),
    .Y(_11543_));
 sky130_fd_sc_hd__nor2_1 _18881_ (.A(_11150_),
    .B(_11543_),
    .Y(_11544_));
 sky130_fd_sc_hd__nand2_1 _18882_ (.A(_09898_),
    .B(_11151_),
    .Y(_11545_));
 sky130_fd_sc_hd__o21ai_4 _18883_ (.A1(_09898_),
    .A2(_11544_),
    .B1(_11545_),
    .Y(_11546_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_690 ();
 sky130_fd_sc_hd__nand2_1 _18885_ (.A(_11472_),
    .B(_11546_),
    .Y(_11548_));
 sky130_fd_sc_hd__a21oi_1 _18886_ (.A1(_11534_),
    .A2(_11548_),
    .B1(_11330_),
    .Y(_11549_));
 sky130_fd_sc_hd__nor2_1 _18887_ (.A(_11530_),
    .B(_11549_),
    .Y(_00026_));
 sky130_fd_sc_hd__nand2_1 _18888_ (.A(\cs_registers_i.mcycle_counter_i.counter[19] ),
    .B(_11533_),
    .Y(_11550_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_689 ();
 sky130_fd_sc_hd__a22o_2 _18890_ (.A1(\cs_registers_i.mtval_q[19] ),
    .A2(_11422_),
    .B1(_11255_),
    .B2(\cs_registers_i.mscratch_q[19] ),
    .X(_11552_));
 sky130_fd_sc_hd__a22oi_2 _18891_ (.A1(\cs_registers_i.mcycle_counter_i.counter[19] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][19] ),
    .Y(_11553_));
 sky130_fd_sc_hd__a22oi_2 _18892_ (.A1(\cs_registers_i.mcycle_counter_i.counter[51] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][51] ),
    .Y(_11554_));
 sky130_fd_sc_hd__o22ai_4 _18893_ (.A1(_10926_),
    .A2(_11553_),
    .B1(_11554_),
    .B2(_10928_),
    .Y(_11555_));
 sky130_fd_sc_hd__a221oi_1 _18894_ (.A1(net72),
    .A2(net1231),
    .B1(_11418_),
    .B2(\cs_registers_i.csr_depc_o[19] ),
    .C1(_10907_),
    .Y(_11556_));
 sky130_fd_sc_hd__a222oi_1 _18895_ (.A1(\cs_registers_i.dscratch0_q[19] ),
    .A2(_11409_),
    .B1(_11416_),
    .B2(\cs_registers_i.dscratch1_q[19] ),
    .C1(\cs_registers_i.mie_q[3] ),
    .C2(_11373_),
    .Y(_11557_));
 sky130_fd_sc_hd__a22oi_1 _18896_ (.A1(\cs_registers_i.csr_mtvec_o[19] ),
    .A2(_10918_),
    .B1(_11384_),
    .B2(net138),
    .Y(_11558_));
 sky130_fd_sc_hd__nand3_1 _18897_ (.A(_11556_),
    .B(_11557_),
    .C(_11558_),
    .Y(_11559_));
 sky130_fd_sc_hd__a2111oi_4 _18898_ (.A1(\cs_registers_i.csr_mepc_o[19] ),
    .A2(_11272_),
    .B1(_11552_),
    .C1(_11555_),
    .D1(_11559_),
    .Y(_11560_));
 sky130_fd_sc_hd__nor2_1 _18899_ (.A(_11150_),
    .B(_11560_),
    .Y(_11561_));
 sky130_fd_sc_hd__nand2_1 _18900_ (.A(_10008_),
    .B(_11151_),
    .Y(_11562_));
 sky130_fd_sc_hd__o21ai_4 _18901_ (.A1(_10008_),
    .A2(_11561_),
    .B1(_11562_),
    .Y(_11563_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_688 ();
 sky130_fd_sc_hd__nand2_1 _18903_ (.A(_11472_),
    .B(_11563_),
    .Y(_11565_));
 sky130_fd_sc_hd__o21ai_0 _18904_ (.A1(net273),
    .A2(_11550_),
    .B1(_11565_),
    .Y(_11566_));
 sky130_fd_sc_hd__nor2_1 _18905_ (.A(_11472_),
    .B(_11533_),
    .Y(_11567_));
 sky130_fd_sc_hd__nor2_1 _18906_ (.A(_11330_),
    .B(_11567_),
    .Y(_11568_));
 sky130_fd_sc_hd__nor2_1 _18907_ (.A(\cs_registers_i.mcycle_counter_i.counter[19] ),
    .B(_11568_),
    .Y(_11569_));
 sky130_fd_sc_hd__a21oi_1 _18908_ (.A1(_11322_),
    .A2(_11566_),
    .B1(_11569_),
    .Y(_00027_));
 sky130_fd_sc_hd__nand2_1 _18909_ (.A(\cs_registers_i.mcycle_counter_i.counter[0] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[1] ),
    .Y(_11570_));
 sky130_fd_sc_hd__a22oi_1 _18910_ (.A1(\cs_registers_i.mcycle_counter_i.counter[1] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][1] ),
    .Y(_11571_));
 sky130_fd_sc_hd__nor2_2 _18911_ (.A(_10926_),
    .B(_11571_),
    .Y(_11572_));
 sky130_fd_sc_hd__a22oi_2 _18912_ (.A1(\cs_registers_i.mcycle_counter_i.counter[33] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][33] ),
    .Y(_11573_));
 sky130_fd_sc_hd__a222oi_1 _18913_ (.A1(net73),
    .A2(_11238_),
    .B1(_11248_),
    .B2(\cs_registers_i.dcsr_q[1] ),
    .C1(\cs_registers_i.csr_depc_o[1] ),
    .C2(_11295_),
    .Y(_11574_));
 sky130_fd_sc_hd__a22oi_1 _18914_ (.A1(\cs_registers_i.dscratch0_q[1] ),
    .A2(_11252_),
    .B1(_11260_),
    .B2(\cs_registers_i.dscratch1_q[1] ),
    .Y(_11575_));
 sky130_fd_sc_hd__o211ai_2 _18915_ (.A1(_11225_),
    .A2(_11573_),
    .B1(_11574_),
    .C1(_11575_),
    .Y(_11576_));
 sky130_fd_sc_hd__a22oi_2 _18916_ (.A1(\cs_registers_i.csr_mepc_o[1] ),
    .A2(_11272_),
    .B1(_11271_),
    .B2(\cs_registers_i.mcause_q[1] ),
    .Y(_11577_));
 sky130_fd_sc_hd__a22oi_2 _18917_ (.A1(\cs_registers_i.mscratch_q[1] ),
    .A2(_11255_),
    .B1(_11270_),
    .B2(\cs_registers_i.mtval_q[1] ),
    .Y(_11578_));
 sky130_fd_sc_hd__nand2_4 _18918_ (.A(_11577_),
    .B(_11578_),
    .Y(_11579_));
 sky130_fd_sc_hd__nor3_4 _18919_ (.A(_11572_),
    .B(_11576_),
    .C(_11579_),
    .Y(_11580_));
 sky130_fd_sc_hd__nand2_1 _18920_ (.A(net778),
    .B(_11146_),
    .Y(_11581_));
 sky130_fd_sc_hd__o22a_4 _18921_ (.A1(net778),
    .A2(_11151_),
    .B1(_11580_),
    .B2(_11581_),
    .X(_11582_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_687 ();
 sky130_fd_sc_hd__nand2_1 _18923_ (.A(_11328_),
    .B(_11582_),
    .Y(_11584_));
 sky130_fd_sc_hd__o21a_1 _18924_ (.A1(_11472_),
    .A2(_11570_),
    .B1(_11584_),
    .X(_11585_));
 sky130_fd_sc_hd__nor2_1 _18925_ (.A(\cs_registers_i.mcycle_counter_i.counter[0] ),
    .B(_11328_),
    .Y(_11586_));
 sky130_fd_sc_hd__nor2_1 _18926_ (.A(_11330_),
    .B(_11586_),
    .Y(_11587_));
 sky130_fd_sc_hd__o22a_1 _18927_ (.A1(_11330_),
    .A2(_11585_),
    .B1(_11587_),
    .B2(\cs_registers_i.mcycle_counter_i.counter[1] ),
    .X(_00028_));
 sky130_fd_sc_hd__a22oi_1 _18928_ (.A1(\cs_registers_i.mcycle_counter_i.counter[20] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][20] ),
    .Y(_11588_));
 sky130_fd_sc_hd__a22oi_1 _18929_ (.A1(\cs_registers_i.mcycle_counter_i.counter[52] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][52] ),
    .Y(_11589_));
 sky130_fd_sc_hd__o22a_2 _18930_ (.A1(_10926_),
    .A2(_11588_),
    .B1(_11589_),
    .B2(_10928_),
    .X(_11590_));
 sky130_fd_sc_hd__a221oi_2 _18931_ (.A1(\cs_registers_i.csr_mtvec_o[20] ),
    .A2(_10918_),
    .B1(_11373_),
    .B2(\cs_registers_i.mie_q[4] ),
    .C1(_11411_),
    .Y(_11591_));
 sky130_fd_sc_hd__a222oi_1 _18932_ (.A1(\cs_registers_i.mtval_q[20] ),
    .A2(_11422_),
    .B1(_11255_),
    .B2(\cs_registers_i.mscratch_q[20] ),
    .C1(_11272_),
    .C2(\cs_registers_i.csr_mepc_o[20] ),
    .Y(_11592_));
 sky130_fd_sc_hd__a22oi_1 _18933_ (.A1(\cs_registers_i.dscratch0_q[20] ),
    .A2(_11409_),
    .B1(_11418_),
    .B2(\cs_registers_i.csr_depc_o[20] ),
    .Y(_11593_));
 sky130_fd_sc_hd__a22oi_1 _18934_ (.A1(net74),
    .A2(net1230),
    .B1(_11416_),
    .B2(\cs_registers_i.dscratch1_q[20] ),
    .Y(_11594_));
 sky130_fd_sc_hd__nand2_1 _18935_ (.A(_11593_),
    .B(_11594_),
    .Y(_11595_));
 sky130_fd_sc_hd__a21oi_1 _18936_ (.A1(net139),
    .A2(_11384_),
    .B1(_11595_),
    .Y(_11596_));
 sky130_fd_sc_hd__nand4_4 _18937_ (.A(_11590_),
    .B(_11591_),
    .C(_11592_),
    .D(_11596_),
    .Y(_11597_));
 sky130_fd_sc_hd__a21oi_1 _18938_ (.A1(_11146_),
    .A2(_11597_),
    .B1(_10070_),
    .Y(_11598_));
 sky130_fd_sc_hd__a21o_4 _18939_ (.A1(_10070_),
    .A2(_11151_),
    .B1(_11598_),
    .X(_11599_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_686 ();
 sky130_fd_sc_hd__nand2_1 _18941_ (.A(_11472_),
    .B(_11599_),
    .Y(_11601_));
 sky130_fd_sc_hd__nand2_1 _18942_ (.A(\cs_registers_i.mcycle_counter_i.counter[19] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[20] ),
    .Y(_11602_));
 sky130_fd_sc_hd__nor3_1 _18943_ (.A(_11454_),
    .B(_11532_),
    .C(_11602_),
    .Y(_11603_));
 sky130_fd_sc_hd__nand2_1 _18944_ (.A(_11394_),
    .B(_11603_),
    .Y(_11604_));
 sky130_fd_sc_hd__nand2_1 _18945_ (.A(_11601_),
    .B(_11604_),
    .Y(_11605_));
 sky130_fd_sc_hd__nand2_1 _18946_ (.A(_11316_),
    .B(_11550_),
    .Y(_11606_));
 sky130_fd_sc_hd__a21oi_1 _18947_ (.A1(_11322_),
    .A2(_11606_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[20] ),
    .Y(_11607_));
 sky130_fd_sc_hd__a21oi_1 _18948_ (.A1(_11322_),
    .A2(_11605_),
    .B1(_11607_),
    .Y(_00029_));
 sky130_fd_sc_hd__nor3_1 _18949_ (.A(_11454_),
    .B(_11532_),
    .C(_11602_),
    .Y(_11608_));
 sky130_fd_sc_hd__nand2_1 _18950_ (.A(\cs_registers_i.mcycle_counter_i.counter[21] ),
    .B(_11608_),
    .Y(_11609_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_685 ();
 sky130_fd_sc_hd__a22oi_1 _18952_ (.A1(\cs_registers_i.csr_mtvec_o[21] ),
    .A2(_10918_),
    .B1(_11375_),
    .B2(\cs_registers_i.csr_mstatus_tw_o ),
    .Y(_11611_));
 sky130_fd_sc_hd__a222oi_1 _18953_ (.A1(\cs_registers_i.dscratch0_q[21] ),
    .A2(_11252_),
    .B1(_11260_),
    .B2(\cs_registers_i.dscratch1_q[21] ),
    .C1(\cs_registers_i.mie_q[5] ),
    .C2(_11373_),
    .Y(_11612_));
 sky130_fd_sc_hd__a221oi_1 _18954_ (.A1(net75),
    .A2(net274),
    .B1(_11295_),
    .B2(\cs_registers_i.csr_depc_o[21] ),
    .C1(_10907_),
    .Y(_11613_));
 sky130_fd_sc_hd__nand3_1 _18955_ (.A(_11611_),
    .B(_11612_),
    .C(_11613_),
    .Y(_11614_));
 sky130_fd_sc_hd__a22oi_2 _18956_ (.A1(\cs_registers_i.mcycle_counter_i.counter[21] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][21] ),
    .Y(_11615_));
 sky130_fd_sc_hd__a22oi_4 _18957_ (.A1(\cs_registers_i.mcycle_counter_i.counter[53] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][53] ),
    .Y(_11616_));
 sky130_fd_sc_hd__o22ai_4 _18958_ (.A1(_10926_),
    .A2(_11615_),
    .B1(_11616_),
    .B2(_11225_),
    .Y(_11617_));
 sky130_fd_sc_hd__a22oi_1 _18959_ (.A1(\cs_registers_i.mscratch_q[21] ),
    .A2(_11255_),
    .B1(_11384_),
    .B2(net140),
    .Y(_11618_));
 sky130_fd_sc_hd__a22oi_1 _18960_ (.A1(\cs_registers_i.csr_mepc_o[21] ),
    .A2(_11272_),
    .B1(_11270_),
    .B2(\cs_registers_i.mtval_q[21] ),
    .Y(_11619_));
 sky130_fd_sc_hd__nand2_1 _18961_ (.A(_11618_),
    .B(_11619_),
    .Y(_11620_));
 sky130_fd_sc_hd__nor3_4 _18962_ (.A(_11614_),
    .B(_11617_),
    .C(_11620_),
    .Y(_11621_));
 sky130_fd_sc_hd__nor3_1 _18963_ (.A(_10145_),
    .B(_11150_),
    .C(_11621_),
    .Y(_11622_));
 sky130_fd_sc_hd__a21oi_4 _18964_ (.A1(_10145_),
    .A2(_11148_),
    .B1(_11622_),
    .Y(_11623_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_684 ();
 sky130_fd_sc_hd__nand2_1 _18966_ (.A(net273),
    .B(_11623_),
    .Y(_11625_));
 sky130_fd_sc_hd__o21ai_0 _18967_ (.A1(_11336_),
    .A2(_11609_),
    .B1(_11625_),
    .Y(_11626_));
 sky130_fd_sc_hd__or3_1 _18968_ (.A(_11454_),
    .B(_11532_),
    .C(_11602_),
    .X(_11627_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_683 ();
 sky130_fd_sc_hd__o21ai_0 _18970_ (.A1(_11392_),
    .A2(_11627_),
    .B1(_11320_),
    .Y(_11629_));
 sky130_fd_sc_hd__a21oi_1 _18971_ (.A1(_11322_),
    .A2(_11629_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[21] ),
    .Y(_11630_));
 sky130_fd_sc_hd__a21oi_1 _18972_ (.A1(_11322_),
    .A2(_11626_),
    .B1(_11630_),
    .Y(_00030_));
 sky130_fd_sc_hd__nand4_1 _18973_ (.A(\cs_registers_i.mcycle_counter_i.counter[21] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[22] ),
    .C(_11335_),
    .D(_11603_),
    .Y(_11631_));
 sky130_fd_sc_hd__a222oi_1 _18974_ (.A1(\cs_registers_i.mtval_q[22] ),
    .A2(_11422_),
    .B1(_11255_),
    .B2(\cs_registers_i.mscratch_q[22] ),
    .C1(_11272_),
    .C2(\cs_registers_i.csr_mepc_o[22] ),
    .Y(_11632_));
 sky130_fd_sc_hd__a22oi_2 _18975_ (.A1(\cs_registers_i.mcycle_counter_i.counter[22] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][22] ),
    .Y(_11633_));
 sky130_fd_sc_hd__a22oi_2 _18976_ (.A1(\cs_registers_i.mcycle_counter_i.counter[54] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][54] ),
    .Y(_11634_));
 sky130_fd_sc_hd__o22ai_4 _18977_ (.A1(_10926_),
    .A2(_11633_),
    .B1(_11634_),
    .B2(_10928_),
    .Y(_11635_));
 sky130_fd_sc_hd__a221oi_1 _18978_ (.A1(net76),
    .A2(net1232),
    .B1(_11418_),
    .B2(\cs_registers_i.csr_depc_o[22] ),
    .C1(_10907_),
    .Y(_11636_));
 sky130_fd_sc_hd__a222oi_1 _18979_ (.A1(\cs_registers_i.dscratch0_q[22] ),
    .A2(_11409_),
    .B1(_11416_),
    .B2(\cs_registers_i.dscratch1_q[22] ),
    .C1(\cs_registers_i.mie_q[6] ),
    .C2(_11373_),
    .Y(_11637_));
 sky130_fd_sc_hd__a22oi_1 _18980_ (.A1(\cs_registers_i.csr_mtvec_o[22] ),
    .A2(_10918_),
    .B1(_11384_),
    .B2(net141),
    .Y(_11638_));
 sky130_fd_sc_hd__nand3_1 _18981_ (.A(_11636_),
    .B(_11637_),
    .C(_11638_),
    .Y(_11639_));
 sky130_fd_sc_hd__nor2_1 _18982_ (.A(_11635_),
    .B(_11639_),
    .Y(_11640_));
 sky130_fd_sc_hd__nand2_4 _18983_ (.A(_11632_),
    .B(_11640_),
    .Y(_11641_));
 sky130_fd_sc_hd__a21oi_1 _18984_ (.A1(_11146_),
    .A2(_11641_),
    .B1(_10172_),
    .Y(_11642_));
 sky130_fd_sc_hd__a21o_4 _18985_ (.A1(_10172_),
    .A2(_11151_),
    .B1(_11642_),
    .X(_11643_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_682 ();
 sky130_fd_sc_hd__nand2_1 _18987_ (.A(_11472_),
    .B(_11643_),
    .Y(_11645_));
 sky130_fd_sc_hd__o21ai_0 _18988_ (.A1(_11472_),
    .A2(_11631_),
    .B1(_11645_),
    .Y(_11646_));
 sky130_fd_sc_hd__o21ai_0 _18989_ (.A1(_11392_),
    .A2(_11609_),
    .B1(_11320_),
    .Y(_11647_));
 sky130_fd_sc_hd__a21oi_1 _18990_ (.A1(_11322_),
    .A2(_11647_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[22] ),
    .Y(_11648_));
 sky130_fd_sc_hd__a21oi_1 _18991_ (.A1(_11322_),
    .A2(_11646_),
    .B1(_11648_),
    .Y(_00031_));
 sky130_fd_sc_hd__nor2_1 _18992_ (.A(_11392_),
    .B(_11609_),
    .Y(_11649_));
 sky130_fd_sc_hd__nand3_2 _18993_ (.A(\cs_registers_i.mcycle_counter_i.counter[22] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[23] ),
    .C(_11649_),
    .Y(_11650_));
 sky130_fd_sc_hd__a222oi_1 _18994_ (.A1(\cs_registers_i.mtval_q[23] ),
    .A2(_11422_),
    .B1(_11255_),
    .B2(\cs_registers_i.mscratch_q[23] ),
    .C1(_11272_),
    .C2(\cs_registers_i.csr_mepc_o[23] ),
    .Y(_11651_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_681 ();
 sky130_fd_sc_hd__a22oi_2 _18996_ (.A1(\cs_registers_i.mcycle_counter_i.counter[23] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][23] ),
    .Y(_11653_));
 sky130_fd_sc_hd__a22oi_2 _18997_ (.A1(\cs_registers_i.mcycle_counter_i.counter[55] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][55] ),
    .Y(_11654_));
 sky130_fd_sc_hd__o22ai_4 _18998_ (.A1(_10926_),
    .A2(_11653_),
    .B1(_11654_),
    .B2(_10928_),
    .Y(_11655_));
 sky130_fd_sc_hd__a221oi_1 _18999_ (.A1(net77),
    .A2(net1230),
    .B1(_11418_),
    .B2(\cs_registers_i.csr_depc_o[23] ),
    .C1(_10907_),
    .Y(_11656_));
 sky130_fd_sc_hd__a222oi_1 _19000_ (.A1(\cs_registers_i.dscratch0_q[23] ),
    .A2(_11409_),
    .B1(_11416_),
    .B2(\cs_registers_i.dscratch1_q[23] ),
    .C1(\cs_registers_i.mie_q[7] ),
    .C2(_11373_),
    .Y(_11657_));
 sky130_fd_sc_hd__a22oi_1 _19001_ (.A1(\cs_registers_i.csr_mtvec_o[23] ),
    .A2(_10918_),
    .B1(_11384_),
    .B2(net142),
    .Y(_11658_));
 sky130_fd_sc_hd__nand3_1 _19002_ (.A(_11656_),
    .B(_11657_),
    .C(_11658_),
    .Y(_11659_));
 sky130_fd_sc_hd__nor2_1 _19003_ (.A(_11655_),
    .B(_11659_),
    .Y(_11660_));
 sky130_fd_sc_hd__nand2_2 _19004_ (.A(_11651_),
    .B(_11660_),
    .Y(_11661_));
 sky130_fd_sc_hd__nand2_1 _19005_ (.A(_11146_),
    .B(_11661_),
    .Y(_11662_));
 sky130_fd_sc_hd__nand2_1 _19006_ (.A(net1236),
    .B(_11662_),
    .Y(_11663_));
 sky130_fd_sc_hd__o21ai_4 _19007_ (.A1(net1236),
    .A2(_11148_),
    .B1(_11663_),
    .Y(_11664_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_680 ();
 sky130_fd_sc_hd__nand2_1 _19009_ (.A(net273),
    .B(_11664_),
    .Y(_11666_));
 sky130_fd_sc_hd__o21ai_0 _19010_ (.A1(net273),
    .A2(_11650_),
    .B1(_11666_),
    .Y(_11667_));
 sky130_fd_sc_hd__nand2_1 _19011_ (.A(\cs_registers_i.mcycle_counter_i.counter[22] ),
    .B(_11649_),
    .Y(_11668_));
 sky130_fd_sc_hd__nand2_1 _19012_ (.A(_11320_),
    .B(_11668_),
    .Y(_11669_));
 sky130_fd_sc_hd__a21oi_1 _19013_ (.A1(_11322_),
    .A2(_11669_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[23] ),
    .Y(_11670_));
 sky130_fd_sc_hd__a21oi_1 _19014_ (.A1(_11322_),
    .A2(_11667_),
    .B1(_11670_),
    .Y(_00032_));
 sky130_fd_sc_hd__nand4_2 _19015_ (.A(\cs_registers_i.mcycle_counter_i.counter[22] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[23] ),
    .C(\cs_registers_i.mcycle_counter_i.counter[24] ),
    .D(_11649_),
    .Y(_11671_));
 sky130_fd_sc_hd__a221oi_4 _19016_ (.A1(net78),
    .A2(net274),
    .B1(_11295_),
    .B2(\cs_registers_i.csr_depc_o[24] ),
    .C1(_10907_),
    .Y(_11672_));
 sky130_fd_sc_hd__nand2_1 _19017_ (.A(\cs_registers_i.mtval_q[24] ),
    .B(_11270_),
    .Y(_11673_));
 sky130_fd_sc_hd__a22oi_1 _19018_ (.A1(\cs_registers_i.csr_mtvec_o[24] ),
    .A2(_10918_),
    .B1(_11252_),
    .B2(\cs_registers_i.dscratch0_q[24] ),
    .Y(_11674_));
 sky130_fd_sc_hd__a22oi_1 _19019_ (.A1(\cs_registers_i.dscratch1_q[24] ),
    .A2(_11260_),
    .B1(_11373_),
    .B2(\cs_registers_i.mie_q[8] ),
    .Y(_11675_));
 sky130_fd_sc_hd__nand4_2 _19020_ (.A(_11672_),
    .B(_11673_),
    .C(_11674_),
    .D(_11675_),
    .Y(_11676_));
 sky130_fd_sc_hd__a22oi_4 _19021_ (.A1(\cs_registers_i.mcycle_counter_i.counter[24] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][24] ),
    .Y(_11677_));
 sky130_fd_sc_hd__a222oi_1 _19022_ (.A1(\cs_registers_i.mscratch_q[24] ),
    .A2(_11255_),
    .B1(_11272_),
    .B2(\cs_registers_i.csr_mepc_o[24] ),
    .C1(net143),
    .C2(_11384_),
    .Y(_11678_));
 sky130_fd_sc_hd__o21ai_1 _19023_ (.A1(_10926_),
    .A2(_11677_),
    .B1(_11678_),
    .Y(_11679_));
 sky130_fd_sc_hd__a22oi_4 _19024_ (.A1(\cs_registers_i.mcycle_counter_i.counter[56] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][56] ),
    .Y(_11680_));
 sky130_fd_sc_hd__nor2_1 _19025_ (.A(_11225_),
    .B(_11680_),
    .Y(_11681_));
 sky130_fd_sc_hd__nor3_4 _19026_ (.A(_11676_),
    .B(_11679_),
    .C(_11681_),
    .Y(_11682_));
 sky130_fd_sc_hd__nor3_1 _19027_ (.A(_10368_),
    .B(_11150_),
    .C(_11682_),
    .Y(_11683_));
 sky130_fd_sc_hd__a21oi_4 _19028_ (.A1(_10368_),
    .A2(_11148_),
    .B1(_11683_),
    .Y(_11684_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_679 ();
 sky130_fd_sc_hd__nand2_1 _19030_ (.A(_11328_),
    .B(_11684_),
    .Y(_11686_));
 sky130_fd_sc_hd__o21ai_0 _19031_ (.A1(_11328_),
    .A2(_11671_),
    .B1(_11686_),
    .Y(_11687_));
 sky130_fd_sc_hd__nand2_1 _19032_ (.A(_11320_),
    .B(_11650_),
    .Y(_11688_));
 sky130_fd_sc_hd__a21oi_1 _19033_ (.A1(_11322_),
    .A2(_11688_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[24] ),
    .Y(_11689_));
 sky130_fd_sc_hd__a21oi_1 _19034_ (.A1(_11322_),
    .A2(_11687_),
    .B1(_11689_),
    .Y(_00033_));
 sky130_fd_sc_hd__inv_1 _19035_ (.A(\cs_registers_i.mcycle_counter_i.counter[24] ),
    .Y(_11690_));
 sky130_fd_sc_hd__nor2_1 _19036_ (.A(_11690_),
    .B(_11650_),
    .Y(_11691_));
 sky130_fd_sc_hd__nand2_1 _19037_ (.A(\cs_registers_i.mcycle_counter_i.counter[25] ),
    .B(_11691_),
    .Y(_11692_));
 sky130_fd_sc_hd__a221oi_1 _19038_ (.A1(net79),
    .A2(net274),
    .B1(_11295_),
    .B2(\cs_registers_i.csr_depc_o[25] ),
    .C1(_10907_),
    .Y(_11693_));
 sky130_fd_sc_hd__nand2_1 _19039_ (.A(\cs_registers_i.mtval_q[25] ),
    .B(_11270_),
    .Y(_11694_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_678 ();
 sky130_fd_sc_hd__a22oi_1 _19041_ (.A1(\cs_registers_i.csr_mtvec_o[25] ),
    .A2(_10918_),
    .B1(_11252_),
    .B2(\cs_registers_i.dscratch0_q[25] ),
    .Y(_11696_));
 sky130_fd_sc_hd__a22oi_4 _19042_ (.A1(\cs_registers_i.dscratch1_q[25] ),
    .A2(_11260_),
    .B1(_11373_),
    .B2(\cs_registers_i.mie_q[9] ),
    .Y(_11697_));
 sky130_fd_sc_hd__nand4_2 _19043_ (.A(_11693_),
    .B(_11694_),
    .C(_11696_),
    .D(_11697_),
    .Y(_11698_));
 sky130_fd_sc_hd__a22oi_4 _19044_ (.A1(\cs_registers_i.mcycle_counter_i.counter[25] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][25] ),
    .Y(_11699_));
 sky130_fd_sc_hd__a222oi_1 _19045_ (.A1(\cs_registers_i.mscratch_q[25] ),
    .A2(_11255_),
    .B1(_11272_),
    .B2(\cs_registers_i.csr_mepc_o[25] ),
    .C1(net144),
    .C2(_11384_),
    .Y(_11700_));
 sky130_fd_sc_hd__o21ai_1 _19046_ (.A1(_10926_),
    .A2(_11699_),
    .B1(_11700_),
    .Y(_11701_));
 sky130_fd_sc_hd__a22oi_4 _19047_ (.A1(\cs_registers_i.mcycle_counter_i.counter[57] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][57] ),
    .Y(_11702_));
 sky130_fd_sc_hd__nor2_1 _19048_ (.A(_11225_),
    .B(_11702_),
    .Y(_11703_));
 sky130_fd_sc_hd__nor3_4 _19049_ (.A(_11698_),
    .B(_11701_),
    .C(_11703_),
    .Y(_11704_));
 sky130_fd_sc_hd__nand2_1 _19050_ (.A(_10303_),
    .B(_11146_),
    .Y(_11705_));
 sky130_fd_sc_hd__o22a_4 _19051_ (.A1(_10303_),
    .A2(_11151_),
    .B1(_11704_),
    .B2(_11705_),
    .X(_11706_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_677 ();
 sky130_fd_sc_hd__nand2_1 _19053_ (.A(_11328_),
    .B(_11706_),
    .Y(_11708_));
 sky130_fd_sc_hd__o21ai_0 _19054_ (.A1(_11328_),
    .A2(_11692_),
    .B1(_11708_),
    .Y(_11709_));
 sky130_fd_sc_hd__nand2_1 _19055_ (.A(_11320_),
    .B(_11671_),
    .Y(_11710_));
 sky130_fd_sc_hd__a21oi_1 _19056_ (.A1(_11322_),
    .A2(_11710_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[25] ),
    .Y(_11711_));
 sky130_fd_sc_hd__a21oi_1 _19057_ (.A1(_11322_),
    .A2(_11709_),
    .B1(_11711_),
    .Y(_00034_));
 sky130_fd_sc_hd__nand3_1 _19058_ (.A(\cs_registers_i.mcycle_counter_i.counter[25] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[26] ),
    .C(_11691_),
    .Y(_11712_));
 sky130_fd_sc_hd__a221oi_4 _19059_ (.A1(net80),
    .A2(net274),
    .B1(_11295_),
    .B2(\cs_registers_i.csr_depc_o[26] ),
    .C1(_10907_),
    .Y(_11713_));
 sky130_fd_sc_hd__nand2_1 _19060_ (.A(\cs_registers_i.mtval_q[26] ),
    .B(_11270_),
    .Y(_11714_));
 sky130_fd_sc_hd__a22oi_1 _19061_ (.A1(\cs_registers_i.csr_mtvec_o[26] ),
    .A2(_10918_),
    .B1(_11252_),
    .B2(\cs_registers_i.dscratch0_q[26] ),
    .Y(_11715_));
 sky130_fd_sc_hd__a22oi_1 _19062_ (.A1(\cs_registers_i.dscratch1_q[26] ),
    .A2(_11260_),
    .B1(_11373_),
    .B2(\cs_registers_i.mie_q[10] ),
    .Y(_11716_));
 sky130_fd_sc_hd__nand4_1 _19063_ (.A(_11713_),
    .B(_11714_),
    .C(_11715_),
    .D(_11716_),
    .Y(_11717_));
 sky130_fd_sc_hd__a22oi_4 _19064_ (.A1(\cs_registers_i.mcycle_counter_i.counter[26] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][26] ),
    .Y(_11718_));
 sky130_fd_sc_hd__a222oi_1 _19065_ (.A1(\cs_registers_i.mscratch_q[26] ),
    .A2(_11255_),
    .B1(_11272_),
    .B2(\cs_registers_i.csr_mepc_o[26] ),
    .C1(net131),
    .C2(_11384_),
    .Y(_11719_));
 sky130_fd_sc_hd__o21ai_1 _19066_ (.A1(_10926_),
    .A2(_11718_),
    .B1(_11719_),
    .Y(_11720_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_676 ();
 sky130_fd_sc_hd__a22oi_4 _19068_ (.A1(\cs_registers_i.mcycle_counter_i.counter[58] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][58] ),
    .Y(_11722_));
 sky130_fd_sc_hd__nor2_1 _19069_ (.A(_11225_),
    .B(_11722_),
    .Y(_11723_));
 sky130_fd_sc_hd__nor3_4 _19070_ (.A(_11717_),
    .B(_11720_),
    .C(_11723_),
    .Y(_11724_));
 sky130_fd_sc_hd__nor3_1 _19071_ (.A(_10468_),
    .B(_11150_),
    .C(_11724_),
    .Y(_11725_));
 sky130_fd_sc_hd__a21oi_4 _19072_ (.A1(_10468_),
    .A2(_11148_),
    .B1(_11725_),
    .Y(_11726_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_675 ();
 sky130_fd_sc_hd__nand2_1 _19074_ (.A(_11328_),
    .B(_11726_),
    .Y(_11728_));
 sky130_fd_sc_hd__o21ai_0 _19075_ (.A1(_11328_),
    .A2(_11712_),
    .B1(_11728_),
    .Y(_11729_));
 sky130_fd_sc_hd__nand2_1 _19076_ (.A(_11320_),
    .B(_11692_),
    .Y(_11730_));
 sky130_fd_sc_hd__a21oi_1 _19077_ (.A1(_11322_),
    .A2(_11730_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[26] ),
    .Y(_11731_));
 sky130_fd_sc_hd__a21oi_1 _19078_ (.A1(_11322_),
    .A2(_11729_),
    .B1(_11731_),
    .Y(_00035_));
 sky130_fd_sc_hd__and3_1 _19079_ (.A(\cs_registers_i.mcycle_counter_i.counter[25] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[26] ),
    .C(_11691_),
    .X(_11732_));
 sky130_fd_sc_hd__nand2_1 _19080_ (.A(\cs_registers_i.mcycle_counter_i.counter[27] ),
    .B(_11732_),
    .Y(_11733_));
 sky130_fd_sc_hd__a221oi_2 _19081_ (.A1(net81),
    .A2(net274),
    .B1(_11295_),
    .B2(\cs_registers_i.csr_depc_o[27] ),
    .C1(_10907_),
    .Y(_11734_));
 sky130_fd_sc_hd__nand2_1 _19082_ (.A(\cs_registers_i.mtval_q[27] ),
    .B(_11270_),
    .Y(_11735_));
 sky130_fd_sc_hd__a22oi_1 _19083_ (.A1(\cs_registers_i.csr_mtvec_o[27] ),
    .A2(_10918_),
    .B1(_11252_),
    .B2(\cs_registers_i.dscratch0_q[27] ),
    .Y(_11736_));
 sky130_fd_sc_hd__a22oi_1 _19084_ (.A1(\cs_registers_i.dscratch1_q[27] ),
    .A2(_11260_),
    .B1(_11373_),
    .B2(\cs_registers_i.mie_q[11] ),
    .Y(_11737_));
 sky130_fd_sc_hd__nand4_1 _19085_ (.A(_11734_),
    .B(_11735_),
    .C(_11736_),
    .D(_11737_),
    .Y(_11738_));
 sky130_fd_sc_hd__a22oi_4 _19086_ (.A1(\cs_registers_i.mcycle_counter_i.counter[27] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][27] ),
    .Y(_11739_));
 sky130_fd_sc_hd__a222oi_1 _19087_ (.A1(\cs_registers_i.mscratch_q[27] ),
    .A2(_11255_),
    .B1(_11272_),
    .B2(\cs_registers_i.csr_mepc_o[27] ),
    .C1(net132),
    .C2(_11384_),
    .Y(_11740_));
 sky130_fd_sc_hd__o21ai_1 _19088_ (.A1(_10926_),
    .A2(_11739_),
    .B1(_11740_),
    .Y(_11741_));
 sky130_fd_sc_hd__a22oi_4 _19089_ (.A1(\cs_registers_i.mcycle_counter_i.counter[59] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][59] ),
    .Y(_11742_));
 sky130_fd_sc_hd__nor2_1 _19090_ (.A(_11225_),
    .B(_11742_),
    .Y(_11743_));
 sky130_fd_sc_hd__nor3_4 _19091_ (.A(_11738_),
    .B(_11741_),
    .C(_11743_),
    .Y(_11744_));
 sky130_fd_sc_hd__nor3_1 _19092_ (.A(_10497_),
    .B(_11150_),
    .C(_11744_),
    .Y(_11745_));
 sky130_fd_sc_hd__a21oi_4 _19093_ (.A1(_10497_),
    .A2(_11148_),
    .B1(_11745_),
    .Y(_11746_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_674 ();
 sky130_fd_sc_hd__nand2_1 _19095_ (.A(_11328_),
    .B(_11746_),
    .Y(_11748_));
 sky130_fd_sc_hd__o21ai_0 _19096_ (.A1(_11328_),
    .A2(_11733_),
    .B1(_11748_),
    .Y(_11749_));
 sky130_fd_sc_hd__nand2_1 _19097_ (.A(_11320_),
    .B(_11712_),
    .Y(_11750_));
 sky130_fd_sc_hd__a21oi_1 _19098_ (.A1(_11322_),
    .A2(_11750_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[27] ),
    .Y(_11751_));
 sky130_fd_sc_hd__a21oi_1 _19099_ (.A1(_11322_),
    .A2(_11749_),
    .B1(_11751_),
    .Y(_00036_));
 sky130_fd_sc_hd__nand3_1 _19100_ (.A(\cs_registers_i.mcycle_counter_i.counter[27] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[28] ),
    .C(_11732_),
    .Y(_11752_));
 sky130_fd_sc_hd__a221oi_2 _19101_ (.A1(net82),
    .A2(net274),
    .B1(_11295_),
    .B2(\cs_registers_i.csr_depc_o[28] ),
    .C1(_10907_),
    .Y(_11753_));
 sky130_fd_sc_hd__nand2_1 _19102_ (.A(\cs_registers_i.mtval_q[28] ),
    .B(_11270_),
    .Y(_11754_));
 sky130_fd_sc_hd__a22oi_1 _19103_ (.A1(\cs_registers_i.csr_mtvec_o[28] ),
    .A2(_10918_),
    .B1(_11252_),
    .B2(\cs_registers_i.dscratch0_q[28] ),
    .Y(_11755_));
 sky130_fd_sc_hd__a22oi_1 _19104_ (.A1(\cs_registers_i.dscratch1_q[28] ),
    .A2(_11260_),
    .B1(_11373_),
    .B2(\cs_registers_i.mie_q[12] ),
    .Y(_11756_));
 sky130_fd_sc_hd__nand4_1 _19105_ (.A(_11753_),
    .B(_11754_),
    .C(_11755_),
    .D(_11756_),
    .Y(_11757_));
 sky130_fd_sc_hd__a22oi_4 _19106_ (.A1(\cs_registers_i.mcycle_counter_i.counter[28] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][28] ),
    .Y(_11758_));
 sky130_fd_sc_hd__a222oi_1 _19107_ (.A1(\cs_registers_i.mscratch_q[28] ),
    .A2(_11255_),
    .B1(_11272_),
    .B2(\cs_registers_i.csr_mepc_o[28] ),
    .C1(net133),
    .C2(_11384_),
    .Y(_11759_));
 sky130_fd_sc_hd__o21ai_1 _19108_ (.A1(_10926_),
    .A2(_11758_),
    .B1(_11759_),
    .Y(_11760_));
 sky130_fd_sc_hd__a22oi_4 _19109_ (.A1(\cs_registers_i.mcycle_counter_i.counter[60] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][60] ),
    .Y(_11761_));
 sky130_fd_sc_hd__nor2_1 _19110_ (.A(_11225_),
    .B(_11761_),
    .Y(_11762_));
 sky130_fd_sc_hd__nor3_4 _19111_ (.A(_11757_),
    .B(_11760_),
    .C(_11762_),
    .Y(_11763_));
 sky130_fd_sc_hd__nor3_1 _19112_ (.A(_10655_),
    .B(_11150_),
    .C(_11763_),
    .Y(_11764_));
 sky130_fd_sc_hd__a21oi_4 _19113_ (.A1(_10655_),
    .A2(_11148_),
    .B1(_11764_),
    .Y(_11765_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_673 ();
 sky130_fd_sc_hd__nand2_1 _19115_ (.A(_11328_),
    .B(_11765_),
    .Y(_11767_));
 sky130_fd_sc_hd__o21ai_0 _19116_ (.A1(_11328_),
    .A2(_11752_),
    .B1(_11767_),
    .Y(_11768_));
 sky130_fd_sc_hd__nand2_1 _19117_ (.A(_11320_),
    .B(_11733_),
    .Y(_11769_));
 sky130_fd_sc_hd__a21oi_1 _19118_ (.A1(_11322_),
    .A2(_11769_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[28] ),
    .Y(_11770_));
 sky130_fd_sc_hd__a21oi_1 _19119_ (.A1(_11322_),
    .A2(_11768_),
    .B1(_11770_),
    .Y(_00037_));
 sky130_fd_sc_hd__nand4_1 _19120_ (.A(\cs_registers_i.mcycle_counter_i.counter[27] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[28] ),
    .C(\cs_registers_i.mcycle_counter_i.counter[29] ),
    .D(_11732_),
    .Y(_11771_));
 sky130_fd_sc_hd__nand2_1 _19121_ (.A(\cs_registers_i.csr_mepc_o[29] ),
    .B(_11272_),
    .Y(_11772_));
 sky130_fd_sc_hd__a22oi_1 _19122_ (.A1(\cs_registers_i.mtval_q[29] ),
    .A2(_11422_),
    .B1(_11255_),
    .B2(\cs_registers_i.mscratch_q[29] ),
    .Y(_11773_));
 sky130_fd_sc_hd__nand2_1 _19123_ (.A(_11772_),
    .B(_11773_),
    .Y(_11774_));
 sky130_fd_sc_hd__a22oi_2 _19124_ (.A1(\cs_registers_i.mcycle_counter_i.counter[29] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][29] ),
    .Y(_11775_));
 sky130_fd_sc_hd__a22oi_2 _19125_ (.A1(\cs_registers_i.mcycle_counter_i.counter[61] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][61] ),
    .Y(_11776_));
 sky130_fd_sc_hd__o22ai_4 _19126_ (.A1(_10926_),
    .A2(_11775_),
    .B1(_11776_),
    .B2(_10928_),
    .Y(_11777_));
 sky130_fd_sc_hd__a221oi_1 _19127_ (.A1(net83),
    .A2(net1230),
    .B1(_11418_),
    .B2(\cs_registers_i.csr_depc_o[29] ),
    .C1(_10907_),
    .Y(_11778_));
 sky130_fd_sc_hd__a222oi_1 _19128_ (.A1(\cs_registers_i.dscratch0_q[29] ),
    .A2(_11409_),
    .B1(_11416_),
    .B2(\cs_registers_i.dscratch1_q[29] ),
    .C1(\cs_registers_i.mie_q[13] ),
    .C2(_11373_),
    .Y(_11779_));
 sky130_fd_sc_hd__a22oi_1 _19129_ (.A1(\cs_registers_i.csr_mtvec_o[29] ),
    .A2(_10918_),
    .B1(_11384_),
    .B2(net134),
    .Y(_11780_));
 sky130_fd_sc_hd__nand3_2 _19130_ (.A(_11778_),
    .B(_11779_),
    .C(_11780_),
    .Y(_11781_));
 sky130_fd_sc_hd__nor3_1 _19131_ (.A(_11774_),
    .B(_11777_),
    .C(_11781_),
    .Y(_11782_));
 sky130_fd_sc_hd__nor2_1 _19132_ (.A(_11150_),
    .B(_11782_),
    .Y(_11783_));
 sky130_fd_sc_hd__nand2_1 _19133_ (.A(_10561_),
    .B(_11151_),
    .Y(_11784_));
 sky130_fd_sc_hd__o21ai_4 _19134_ (.A1(_10561_),
    .A2(_11783_),
    .B1(_11784_),
    .Y(_11785_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_672 ();
 sky130_fd_sc_hd__nand2_1 _19136_ (.A(_11328_),
    .B(_11785_),
    .Y(_11787_));
 sky130_fd_sc_hd__o21ai_0 _19137_ (.A1(_11328_),
    .A2(_11771_),
    .B1(_11787_),
    .Y(_11788_));
 sky130_fd_sc_hd__nand2_1 _19138_ (.A(_11320_),
    .B(_11752_),
    .Y(_11789_));
 sky130_fd_sc_hd__a21oi_1 _19139_ (.A1(_11322_),
    .A2(_11789_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[29] ),
    .Y(_11790_));
 sky130_fd_sc_hd__a21oi_1 _19140_ (.A1(_11322_),
    .A2(_11788_),
    .B1(_11790_),
    .Y(_00038_));
 sky130_fd_sc_hd__nand2_1 _19141_ (.A(_11309_),
    .B(_11472_),
    .Y(_11791_));
 sky130_fd_sc_hd__o21a_1 _19142_ (.A1(_11328_),
    .A2(_11334_),
    .B1(_11791_),
    .X(_11792_));
 sky130_fd_sc_hd__a21oi_1 _19143_ (.A1(_11320_),
    .A2(_11570_),
    .B1(_11330_),
    .Y(_11793_));
 sky130_fd_sc_hd__o22a_1 _19144_ (.A1(_11330_),
    .A2(_11792_),
    .B1(_11793_),
    .B2(\cs_registers_i.mcycle_counter_i.counter[2] ),
    .X(_00039_));
 sky130_fd_sc_hd__a21oi_1 _19145_ (.A1(_11320_),
    .A2(_11771_),
    .B1(_11330_),
    .Y(_11794_));
 sky130_fd_sc_hd__nor2_1 _19146_ (.A(_11328_),
    .B(_11771_),
    .Y(_11795_));
 sky130_fd_sc_hd__a22oi_2 _19147_ (.A1(\cs_registers_i.mcycle_counter_i.counter[30] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][30] ),
    .Y(_11796_));
 sky130_fd_sc_hd__a22oi_2 _19148_ (.A1(\cs_registers_i.mcycle_counter_i.counter[62] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][62] ),
    .Y(_11797_));
 sky130_fd_sc_hd__o22ai_4 _19149_ (.A1(_10926_),
    .A2(_11796_),
    .B1(_11797_),
    .B2(_10928_),
    .Y(_11798_));
 sky130_fd_sc_hd__a22oi_1 _19150_ (.A1(\cs_registers_i.csr_mtvec_o[30] ),
    .A2(_10918_),
    .B1(_11373_),
    .B2(\cs_registers_i.mie_q[14] ),
    .Y(_11799_));
 sky130_fd_sc_hd__a21oi_1 _19151_ (.A1(\cs_registers_i.dscratch1_q[30] ),
    .A2(_11416_),
    .B1(_11410_),
    .Y(_11800_));
 sky130_fd_sc_hd__a222oi_1 _19152_ (.A1(\cs_registers_i.mtval_q[30] ),
    .A2(_11422_),
    .B1(_11255_),
    .B2(\cs_registers_i.mscratch_q[30] ),
    .C1(_11272_),
    .C2(\cs_registers_i.csr_mepc_o[30] ),
    .Y(_11801_));
 sky130_fd_sc_hd__nand4_1 _19153_ (.A(_10908_),
    .B(_11799_),
    .C(_11800_),
    .D(_11801_),
    .Y(_11802_));
 sky130_fd_sc_hd__nor2_1 _19154_ (.A(_11798_),
    .B(_11802_),
    .Y(_11803_));
 sky130_fd_sc_hd__nand2_1 _19155_ (.A(net135),
    .B(_11384_),
    .Y(_11804_));
 sky130_fd_sc_hd__a222oi_1 _19156_ (.A1(\cs_registers_i.dscratch0_q[30] ),
    .A2(_11409_),
    .B1(_11418_),
    .B2(\cs_registers_i.csr_depc_o[30] ),
    .C1(net85),
    .C2(net1230),
    .Y(_11805_));
 sky130_fd_sc_hd__nand3_4 _19157_ (.A(_11803_),
    .B(_11804_),
    .C(_11805_),
    .Y(_11806_));
 sky130_fd_sc_hd__a21oi_1 _19158_ (.A1(_11146_),
    .A2(_11806_),
    .B1(_10799_),
    .Y(_11807_));
 sky130_fd_sc_hd__a21o_4 _19159_ (.A1(_10799_),
    .A2(_11151_),
    .B1(_11807_),
    .X(_11808_));
 sky130_fd_sc_hd__a22oi_1 _19160_ (.A1(\cs_registers_i.mcycle_counter_i.counter[30] ),
    .A2(_11795_),
    .B1(_11808_),
    .B2(_11328_),
    .Y(_11809_));
 sky130_fd_sc_hd__o22a_1 _19161_ (.A1(\cs_registers_i.mcycle_counter_i.counter[30] ),
    .A2(_11794_),
    .B1(_11809_),
    .B2(_11330_),
    .X(_00040_));
 sky130_fd_sc_hd__nand4_1 _19162_ (.A(\cs_registers_i.mcycle_counter_i.counter[27] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[28] ),
    .C(\cs_registers_i.mcycle_counter_i.counter[29] ),
    .D(\cs_registers_i.mcycle_counter_i.counter[30] ),
    .Y(_11810_));
 sky130_fd_sc_hd__nand2_1 _19163_ (.A(\cs_registers_i.mcycle_counter_i.counter[25] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[26] ),
    .Y(_11811_));
 sky130_fd_sc_hd__nor3_1 _19164_ (.A(_11671_),
    .B(_11810_),
    .C(_11811_),
    .Y(_11812_));
 sky130_fd_sc_hd__nor2_1 _19165_ (.A(_11328_),
    .B(_11812_),
    .Y(_11813_));
 sky130_fd_sc_hd__nor2_1 _19166_ (.A(_11330_),
    .B(_11813_),
    .Y(_11814_));
 sky130_fd_sc_hd__a221oi_4 _19167_ (.A1(net86),
    .A2(net274),
    .B1(_11295_),
    .B2(\cs_registers_i.csr_depc_o[31] ),
    .C1(_10907_),
    .Y(_11815_));
 sky130_fd_sc_hd__a22oi_1 _19168_ (.A1(\cs_registers_i.csr_mtvec_o[31] ),
    .A2(_10918_),
    .B1(_11260_),
    .B2(\cs_registers_i.dscratch1_q[31] ),
    .Y(_11816_));
 sky130_fd_sc_hd__a22oi_1 _19169_ (.A1(\cs_registers_i.mscratch_q[31] ),
    .A2(_11255_),
    .B1(_11252_),
    .B2(\cs_registers_i.dscratch0_q[31] ),
    .Y(_11817_));
 sky130_fd_sc_hd__nand3_1 _19170_ (.A(_11815_),
    .B(_11816_),
    .C(_11817_),
    .Y(_11818_));
 sky130_fd_sc_hd__a22oi_4 _19171_ (.A1(\cs_registers_i.mcycle_counter_i.counter[31] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][31] ),
    .Y(_11819_));
 sky130_fd_sc_hd__a222oi_1 _19172_ (.A1(\cs_registers_i.mtval_q[31] ),
    .A2(_11270_),
    .B1(_11271_),
    .B2(\cs_registers_i.mcause_q[5] ),
    .C1(\cs_registers_i.csr_mepc_o[31] ),
    .C2(_11272_),
    .Y(_11820_));
 sky130_fd_sc_hd__o21ai_1 _19173_ (.A1(_10926_),
    .A2(_11819_),
    .B1(_11820_),
    .Y(_11821_));
 sky130_fd_sc_hd__a22oi_4 _19174_ (.A1(\cs_registers_i.mcycle_counter_i.counter[63] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][63] ),
    .Y(_11822_));
 sky130_fd_sc_hd__nor2_1 _19175_ (.A(_11225_),
    .B(_11822_),
    .Y(_11823_));
 sky130_fd_sc_hd__nor3_4 _19176_ (.A(_11818_),
    .B(_11821_),
    .C(_11823_),
    .Y(_11824_));
 sky130_fd_sc_hd__nand2_1 _19177_ (.A(_10695_),
    .B(_11148_),
    .Y(_11825_));
 sky130_fd_sc_hd__o31a_4 _19178_ (.A1(_10695_),
    .A2(_11150_),
    .A3(_11824_),
    .B1(_11825_),
    .X(_11826_));
 sky130_fd_sc_hd__nand2_1 _19179_ (.A(\cs_registers_i.mcycle_counter_i.counter[31] ),
    .B(_11812_),
    .Y(_11827_));
 sky130_fd_sc_hd__nor2_1 _19180_ (.A(_11328_),
    .B(_11827_),
    .Y(_11828_));
 sky130_fd_sc_hd__a21oi_1 _19181_ (.A1(_11328_),
    .A2(_11826_),
    .B1(_11828_),
    .Y(_11829_));
 sky130_fd_sc_hd__o22a_1 _19182_ (.A1(\cs_registers_i.mcycle_counter_i.counter[31] ),
    .A2(_11814_),
    .B1(_11829_),
    .B2(_11330_),
    .X(_00041_));
 sky130_fd_sc_hd__nand2_1 _19183_ (.A(net271),
    .B(_11264_),
    .Y(_11830_));
 sky130_fd_sc_hd__inv_1 _19184_ (.A(\cs_registers_i.mcountinhibit[0] ),
    .Y(_11831_));
 sky130_fd_sc_hd__o21ai_1 _19185_ (.A1(_10926_),
    .A2(_11830_),
    .B1(_11831_),
    .Y(_11832_));
 sky130_fd_sc_hd__o21ai_4 _19186_ (.A1(_11225_),
    .A2(_11830_),
    .B1(_11832_),
    .Y(_11833_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_671 ();
 sky130_fd_sc_hd__a22o_1 _19188_ (.A1(_11280_),
    .A2(_11328_),
    .B1(_11828_),
    .B2(\cs_registers_i.mcycle_counter_i.counter[32] ),
    .X(_11835_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_669 ();
 sky130_fd_sc_hd__nand2_1 _19191_ (.A(_11320_),
    .B(_11827_),
    .Y(_11838_));
 sky130_fd_sc_hd__a21oi_1 _19192_ (.A1(_11833_),
    .A2(_11838_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[32] ),
    .Y(_11839_));
 sky130_fd_sc_hd__a21oi_1 _19193_ (.A1(_11833_),
    .A2(_11835_),
    .B1(_11839_),
    .Y(_00042_));
 sky130_fd_sc_hd__nor2_1 _19194_ (.A(_11810_),
    .B(_11811_),
    .Y(_11840_));
 sky130_fd_sc_hd__nand4_1 _19195_ (.A(\cs_registers_i.mcycle_counter_i.counter[32] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[24] ),
    .C(\cs_registers_i.mcycle_counter_i.counter[31] ),
    .D(_11840_),
    .Y(_11841_));
 sky130_fd_sc_hd__nand3_1 _19196_ (.A(\cs_registers_i.mcycle_counter_i.counter[33] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[22] ),
    .C(\cs_registers_i.mcycle_counter_i.counter[23] ),
    .Y(_11842_));
 sky130_fd_sc_hd__nor2_1 _19197_ (.A(_11841_),
    .B(_11842_),
    .Y(_11843_));
 sky130_fd_sc_hd__nand3_1 _19198_ (.A(\cs_registers_i.mcycle_counter_i.counter[21] ),
    .B(_11608_),
    .C(_11843_),
    .Y(_11844_));
 sky130_fd_sc_hd__o21ai_0 _19199_ (.A1(_11336_),
    .A2(_11844_),
    .B1(_11584_),
    .Y(_11845_));
 sky130_fd_sc_hd__o21ai_0 _19200_ (.A1(_11650_),
    .A2(_11841_),
    .B1(_11320_),
    .Y(_11846_));
 sky130_fd_sc_hd__a21oi_1 _19201_ (.A1(net268),
    .A2(_11846_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[33] ),
    .Y(_11847_));
 sky130_fd_sc_hd__a21oi_1 _19202_ (.A1(net268),
    .A2(_11845_),
    .B1(_11847_),
    .Y(_00043_));
 sky130_fd_sc_hd__nand4_1 _19203_ (.A(\cs_registers_i.mcycle_counter_i.counter[34] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[21] ),
    .C(_11603_),
    .D(_11843_),
    .Y(_11848_));
 sky130_fd_sc_hd__o21ai_0 _19204_ (.A1(_11336_),
    .A2(_11848_),
    .B1(_11791_),
    .Y(_11849_));
 sky130_fd_sc_hd__o21ai_0 _19205_ (.A1(_11392_),
    .A2(_11844_),
    .B1(_11320_),
    .Y(_11850_));
 sky130_fd_sc_hd__a21oi_1 _19206_ (.A1(net268),
    .A2(_11850_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[34] ),
    .Y(_11851_));
 sky130_fd_sc_hd__a21oi_1 _19207_ (.A1(net268),
    .A2(_11849_),
    .B1(_11851_),
    .Y(_00044_));
 sky130_fd_sc_hd__inv_1 _19208_ (.A(\cs_registers_i.mcause_q[3] ),
    .Y(_11852_));
 sky130_fd_sc_hd__nor3_1 _19209_ (.A(_11852_),
    .B(_10889_),
    .C(_11266_),
    .Y(_11853_));
 sky130_fd_sc_hd__a21oi_1 _19210_ (.A1(\cs_registers_i.csr_mepc_o[3] ),
    .A2(_11272_),
    .B1(_11853_),
    .Y(_11854_));
 sky130_fd_sc_hd__a22oi_2 _19211_ (.A1(\cs_registers_i.mtval_q[3] ),
    .A2(_11422_),
    .B1(_11384_),
    .B2(net146),
    .Y(_11855_));
 sky130_fd_sc_hd__a22oi_2 _19212_ (.A1(\cs_registers_i.mcycle_counter_i.counter[3] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][3] ),
    .Y(_11856_));
 sky130_fd_sc_hd__a22oi_2 _19213_ (.A1(\cs_registers_i.mcycle_counter_i.counter[35] ),
    .A2(_11264_),
    .B1(net284),
    .B2(\cs_registers_i.mhpmcounter[2][35] ),
    .Y(_11857_));
 sky130_fd_sc_hd__o22ai_4 _19214_ (.A1(_10926_),
    .A2(_11856_),
    .B1(_11857_),
    .B2(_10928_),
    .Y(_11858_));
 sky130_fd_sc_hd__a221oi_1 _19215_ (.A1(\cs_registers_i.dscratch1_q[3] ),
    .A2(_11416_),
    .B1(_11418_),
    .B2(\cs_registers_i.csr_depc_o[3] ),
    .C1(_10907_),
    .Y(_11859_));
 sky130_fd_sc_hd__a222oi_1 _19216_ (.A1(net87),
    .A2(net1229),
    .B1(_11409_),
    .B2(\cs_registers_i.dscratch0_q[3] ),
    .C1(\cs_registers_i.mie_q[17] ),
    .C2(_11373_),
    .Y(_11860_));
 sky130_fd_sc_hd__a22oi_1 _19217_ (.A1(\cs_registers_i.mscratch_q[3] ),
    .A2(_11255_),
    .B1(_11375_),
    .B2(\cs_registers_i.csr_mstatus_mie_o ),
    .Y(_11861_));
 sky130_fd_sc_hd__nand3_1 _19218_ (.A(_11859_),
    .B(_11860_),
    .C(_11861_),
    .Y(_11862_));
 sky130_fd_sc_hd__nor2_1 _19219_ (.A(_11858_),
    .B(_11862_),
    .Y(_11863_));
 sky130_fd_sc_hd__nand3_4 _19220_ (.A(_11854_),
    .B(_11855_),
    .C(_11863_),
    .Y(_11864_));
 sky130_fd_sc_hd__nand2_1 _19221_ (.A(_11146_),
    .B(_11864_),
    .Y(_11865_));
 sky130_fd_sc_hd__nand2_1 _19222_ (.A(_08636_),
    .B(_11865_),
    .Y(_11866_));
 sky130_fd_sc_hd__o21ai_4 _19223_ (.A1(_08636_),
    .A2(_11148_),
    .B1(_11866_),
    .Y(_11867_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_668 ();
 sky130_fd_sc_hd__nand2_1 _19225_ (.A(net273),
    .B(_11867_),
    .Y(_11869_));
 sky130_fd_sc_hd__nand4_1 _19226_ (.A(\cs_registers_i.mcycle_counter_i.counter[34] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[35] ),
    .C(\cs_registers_i.mcycle_counter_i.counter[21] ),
    .D(_11843_),
    .Y(_11870_));
 sky130_fd_sc_hd__nor2_2 _19227_ (.A(_11627_),
    .B(_11870_),
    .Y(_11871_));
 sky130_fd_sc_hd__nand2_1 _19228_ (.A(_11394_),
    .B(_11871_),
    .Y(_11872_));
 sky130_fd_sc_hd__nand2_1 _19229_ (.A(_11869_),
    .B(_11872_),
    .Y(_11873_));
 sky130_fd_sc_hd__o21ai_0 _19230_ (.A1(_11392_),
    .A2(_11848_),
    .B1(_11316_),
    .Y(_11874_));
 sky130_fd_sc_hd__a21oi_1 _19231_ (.A1(net268),
    .A2(_11874_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[35] ),
    .Y(_11875_));
 sky130_fd_sc_hd__a21oi_1 _19232_ (.A1(net268),
    .A2(_11873_),
    .B1(_11875_),
    .Y(_00045_));
 sky130_fd_sc_hd__nand2_1 _19233_ (.A(\cs_registers_i.mcycle_counter_i.counter[36] ),
    .B(_11871_),
    .Y(_11876_));
 sky130_fd_sc_hd__a22oi_2 _19234_ (.A1(\cs_registers_i.mcycle_counter_i.counter[36] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][36] ),
    .Y(_11877_));
 sky130_fd_sc_hd__a22oi_2 _19235_ (.A1(\cs_registers_i.mcycle_counter_i.counter[4] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][4] ),
    .Y(_11878_));
 sky130_fd_sc_hd__a221o_2 _19236_ (.A1(net88),
    .A2(net274),
    .B1(_11295_),
    .B2(\cs_registers_i.csr_depc_o[4] ),
    .C1(_10907_),
    .X(_11879_));
 sky130_fd_sc_hd__a221oi_2 _19237_ (.A1(\cs_registers_i.dscratch0_q[4] ),
    .A2(_11252_),
    .B1(_11260_),
    .B2(\cs_registers_i.dscratch1_q[4] ),
    .C1(_11879_),
    .Y(_11880_));
 sky130_fd_sc_hd__o221ai_4 _19238_ (.A1(_11225_),
    .A2(_11877_),
    .B1(_11878_),
    .B2(_10926_),
    .C1(_11880_),
    .Y(_11881_));
 sky130_fd_sc_hd__a22oi_1 _19239_ (.A1(\cs_registers_i.mscratch_q[4] ),
    .A2(_11255_),
    .B1(_11271_),
    .B2(\cs_registers_i.mcause_q[4] ),
    .Y(_11882_));
 sky130_fd_sc_hd__a22oi_1 _19240_ (.A1(\cs_registers_i.csr_mepc_o[4] ),
    .A2(_11272_),
    .B1(_11270_),
    .B2(\cs_registers_i.mtval_q[4] ),
    .Y(_11883_));
 sky130_fd_sc_hd__nand2_1 _19241_ (.A(_11882_),
    .B(_11883_),
    .Y(_11884_));
 sky130_fd_sc_hd__nor2_4 _19242_ (.A(_11881_),
    .B(_11884_),
    .Y(_11885_));
 sky130_fd_sc_hd__nand2_1 _19243_ (.A(_08585_),
    .B(_11146_),
    .Y(_11886_));
 sky130_fd_sc_hd__o22a_4 _19244_ (.A1(_08585_),
    .A2(_11151_),
    .B1(_11885_),
    .B2(_11886_),
    .X(_11887_));
 sky130_fd_sc_hd__nand2_1 _19245_ (.A(net273),
    .B(_11887_),
    .Y(_11888_));
 sky130_fd_sc_hd__o21ai_0 _19246_ (.A1(_11336_),
    .A2(_11876_),
    .B1(_11888_),
    .Y(_11889_));
 sky130_fd_sc_hd__nand2_1 _19247_ (.A(_11335_),
    .B(_11871_),
    .Y(_11890_));
 sky130_fd_sc_hd__nand2_1 _19248_ (.A(_11320_),
    .B(_11890_),
    .Y(_11891_));
 sky130_fd_sc_hd__a21oi_1 _19249_ (.A1(net268),
    .A2(_11891_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[36] ),
    .Y(_11892_));
 sky130_fd_sc_hd__a21oi_1 _19250_ (.A1(net268),
    .A2(_11889_),
    .B1(_11892_),
    .Y(_00046_));
 sky130_fd_sc_hd__a221oi_1 _19251_ (.A1(net89),
    .A2(_11238_),
    .B1(_11295_),
    .B2(\cs_registers_i.csr_depc_o[5] ),
    .C1(_10907_),
    .Y(_11893_));
 sky130_fd_sc_hd__a22oi_1 _19252_ (.A1(\cs_registers_i.dscratch0_q[5] ),
    .A2(_11252_),
    .B1(_11260_),
    .B2(\cs_registers_i.dscratch1_q[5] ),
    .Y(_11894_));
 sky130_fd_sc_hd__a222oi_1 _19253_ (.A1(\cs_registers_i.mscratch_q[5] ),
    .A2(_11255_),
    .B1(_11272_),
    .B2(\cs_registers_i.csr_mepc_o[5] ),
    .C1(\cs_registers_i.mtval_q[5] ),
    .C2(_11270_),
    .Y(_11895_));
 sky130_fd_sc_hd__nand3_1 _19254_ (.A(_11893_),
    .B(_11894_),
    .C(_11895_),
    .Y(_11896_));
 sky130_fd_sc_hd__a22oi_2 _19255_ (.A1(\cs_registers_i.mcycle_counter_i.counter[37] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][37] ),
    .Y(_11897_));
 sky130_fd_sc_hd__a22oi_2 _19256_ (.A1(\cs_registers_i.mcycle_counter_i.counter[5] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][5] ),
    .Y(_11898_));
 sky130_fd_sc_hd__o22ai_4 _19257_ (.A1(_11225_),
    .A2(_11897_),
    .B1(_11898_),
    .B2(_10926_),
    .Y(_11899_));
 sky130_fd_sc_hd__nor2_4 _19258_ (.A(_11896_),
    .B(_11899_),
    .Y(_11900_));
 sky130_fd_sc_hd__nor3_1 _19259_ (.A(net952),
    .B(_11150_),
    .C(_11900_),
    .Y(_11901_));
 sky130_fd_sc_hd__a21o_4 _19260_ (.A1(net953),
    .A2(_11148_),
    .B1(_11901_),
    .X(_11902_));
 sky130_fd_sc_hd__nand3_1 _19261_ (.A(\cs_registers_i.mcycle_counter_i.counter[36] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[37] ),
    .C(_11871_),
    .Y(_11903_));
 sky130_fd_sc_hd__o22ai_1 _19262_ (.A1(_11320_),
    .A2(_11902_),
    .B1(_11903_),
    .B2(_11336_),
    .Y(_11904_));
 sky130_fd_sc_hd__o21ai_0 _19263_ (.A1(_11392_),
    .A2(_11876_),
    .B1(_11320_),
    .Y(_11905_));
 sky130_fd_sc_hd__a21oi_1 _19264_ (.A1(net268),
    .A2(_11905_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[37] ),
    .Y(_11906_));
 sky130_fd_sc_hd__a21oi_1 _19265_ (.A1(net268),
    .A2(_11904_),
    .B1(_11906_),
    .Y(_00047_));
 sky130_fd_sc_hd__a21oi_1 _19266_ (.A1(\cs_registers_i.csr_depc_o[6] ),
    .A2(_11295_),
    .B1(_10907_),
    .Y(_11907_));
 sky130_fd_sc_hd__a22oi_1 _19267_ (.A1(net90),
    .A2(_11238_),
    .B1(_11248_),
    .B2(\cs_registers_i.dcsr_q[6] ),
    .Y(_11908_));
 sky130_fd_sc_hd__a22oi_1 _19268_ (.A1(\cs_registers_i.dscratch0_q[6] ),
    .A2(_11252_),
    .B1(_11260_),
    .B2(\cs_registers_i.dscratch1_q[6] ),
    .Y(_11909_));
 sky130_fd_sc_hd__a222oi_1 _19269_ (.A1(\cs_registers_i.mscratch_q[6] ),
    .A2(_11255_),
    .B1(_11272_),
    .B2(\cs_registers_i.csr_mepc_o[6] ),
    .C1(\cs_registers_i.mtval_q[6] ),
    .C2(_11270_),
    .Y(_11910_));
 sky130_fd_sc_hd__nand4_1 _19270_ (.A(_11907_),
    .B(_11908_),
    .C(_11909_),
    .D(_11910_),
    .Y(_11911_));
 sky130_fd_sc_hd__a22oi_2 _19271_ (.A1(\cs_registers_i.mcycle_counter_i.counter[38] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][38] ),
    .Y(_11912_));
 sky130_fd_sc_hd__a22oi_2 _19272_ (.A1(\cs_registers_i.mcycle_counter_i.counter[6] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][6] ),
    .Y(_11913_));
 sky130_fd_sc_hd__o22ai_4 _19273_ (.A1(_11225_),
    .A2(_11912_),
    .B1(_11913_),
    .B2(_10926_),
    .Y(_11914_));
 sky130_fd_sc_hd__nor2_4 _19274_ (.A(_11911_),
    .B(_11914_),
    .Y(_11915_));
 sky130_fd_sc_hd__nand2_1 _19275_ (.A(_08547_),
    .B(_11148_),
    .Y(_11916_));
 sky130_fd_sc_hd__o31ai_4 _19276_ (.A1(_08547_),
    .A2(_11150_),
    .A3(_11915_),
    .B1(_11916_),
    .Y(_11917_));
 sky130_fd_sc_hd__nand4_4 _19277_ (.A(\cs_registers_i.mcycle_counter_i.counter[36] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[37] ),
    .C(\cs_registers_i.mcycle_counter_i.counter[38] ),
    .D(_11871_),
    .Y(_11918_));
 sky130_fd_sc_hd__o22ai_1 _19278_ (.A1(_11320_),
    .A2(_11917_),
    .B1(_11918_),
    .B2(_11336_),
    .Y(_11919_));
 sky130_fd_sc_hd__o21ai_0 _19279_ (.A1(_11392_),
    .A2(_11903_),
    .B1(_11320_),
    .Y(_11920_));
 sky130_fd_sc_hd__a21oi_1 _19280_ (.A1(net268),
    .A2(_11920_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[38] ),
    .Y(_11921_));
 sky130_fd_sc_hd__a21oi_1 _19281_ (.A1(net268),
    .A2(_11919_),
    .B1(_11921_),
    .Y(_00048_));
 sky130_fd_sc_hd__a22oi_2 _19282_ (.A1(\cs_registers_i.mcycle_counter_i.counter[7] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][7] ),
    .Y(_11922_));
 sky130_fd_sc_hd__nor2_4 _19283_ (.A(_10926_),
    .B(_11922_),
    .Y(_11923_));
 sky130_fd_sc_hd__nand2_1 _19284_ (.A(\cs_registers_i.mscratch_q[7] ),
    .B(_11255_),
    .Y(_11924_));
 sky130_fd_sc_hd__a21oi_1 _19285_ (.A1(net91),
    .A2(_11238_),
    .B1(_10907_),
    .Y(_11925_));
 sky130_fd_sc_hd__a22oi_2 _19286_ (.A1(\cs_registers_i.dcsr_q[7] ),
    .A2(_11248_),
    .B1(_11295_),
    .B2(\cs_registers_i.csr_depc_o[7] ),
    .Y(_11926_));
 sky130_fd_sc_hd__a22o_1 _19287_ (.A1(\cs_registers_i.dscratch1_q[7] ),
    .A2(_11260_),
    .B1(_11375_),
    .B2(\cs_registers_i.mstack_d[2] ),
    .X(_11927_));
 sky130_fd_sc_hd__a221oi_1 _19288_ (.A1(\cs_registers_i.dscratch0_q[7] ),
    .A2(_11252_),
    .B1(_11373_),
    .B2(\cs_registers_i.mie_q[16] ),
    .C1(_11927_),
    .Y(_11928_));
 sky130_fd_sc_hd__nand4_2 _19289_ (.A(_11924_),
    .B(_11925_),
    .C(_11926_),
    .D(_11928_),
    .Y(_11929_));
 sky130_fd_sc_hd__a22oi_4 _19290_ (.A1(\cs_registers_i.mcycle_counter_i.counter[39] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][39] ),
    .Y(_11930_));
 sky130_fd_sc_hd__a222oi_1 _19291_ (.A1(\cs_registers_i.csr_mepc_o[7] ),
    .A2(_11272_),
    .B1(_11270_),
    .B2(\cs_registers_i.mtval_q[7] ),
    .C1(net147),
    .C2(_11384_),
    .Y(_11931_));
 sky130_fd_sc_hd__o21ai_1 _19292_ (.A1(_11225_),
    .A2(_11930_),
    .B1(_11931_),
    .Y(_11932_));
 sky130_fd_sc_hd__nor3_4 _19293_ (.A(_11923_),
    .B(_11929_),
    .C(_11932_),
    .Y(_11933_));
 sky130_fd_sc_hd__nor3_1 _19294_ (.A(_08375_),
    .B(_11150_),
    .C(_11933_),
    .Y(_11934_));
 sky130_fd_sc_hd__a21oi_4 _19295_ (.A1(_08375_),
    .A2(_11148_),
    .B1(_11934_),
    .Y(_11935_));
 sky130_fd_sc_hd__inv_1 _19296_ (.A(\cs_registers_i.mcycle_counter_i.counter[39] ),
    .Y(_11936_));
 sky130_fd_sc_hd__nor2_1 _19297_ (.A(_11936_),
    .B(_11918_),
    .Y(_11937_));
 sky130_fd_sc_hd__a22o_1 _19298_ (.A1(net273),
    .A2(_11935_),
    .B1(_11937_),
    .B2(_11394_),
    .X(_11938_));
 sky130_fd_sc_hd__o21ai_0 _19299_ (.A1(_11392_),
    .A2(_11918_),
    .B1(_11320_),
    .Y(_11939_));
 sky130_fd_sc_hd__a21oi_1 _19300_ (.A1(net268),
    .A2(_11939_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[39] ),
    .Y(_11940_));
 sky130_fd_sc_hd__a21oi_1 _19301_ (.A1(net268),
    .A2(_11938_),
    .B1(_11940_),
    .Y(_00049_));
 sky130_fd_sc_hd__nand2_1 _19302_ (.A(_11320_),
    .B(_11334_),
    .Y(_11941_));
 sky130_fd_sc_hd__a21oi_1 _19303_ (.A1(_11322_),
    .A2(_11941_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[3] ),
    .Y(_11942_));
 sky130_fd_sc_hd__a21oi_1 _19304_ (.A1(_11336_),
    .A2(_11869_),
    .B1(_11330_),
    .Y(_11943_));
 sky130_fd_sc_hd__nor2_1 _19305_ (.A(_11942_),
    .B(_11943_),
    .Y(_00050_));
 sky130_fd_sc_hd__nand2_1 _19306_ (.A(\cs_registers_i.mcycle_counter_i.counter[40] ),
    .B(_11937_),
    .Y(_11944_));
 sky130_fd_sc_hd__a22oi_4 _19307_ (.A1(\cs_registers_i.mcycle_counter_i.counter[8] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][8] ),
    .Y(_11945_));
 sky130_fd_sc_hd__a21oi_1 _19308_ (.A1(\cs_registers_i.dscratch0_q[8] ),
    .A2(_11252_),
    .B1(_11411_),
    .Y(_11946_));
 sky130_fd_sc_hd__a22oi_2 _19309_ (.A1(\cs_registers_i.csr_mtvec_o[8] ),
    .A2(_10918_),
    .B1(_11260_),
    .B2(\cs_registers_i.dscratch1_q[8] ),
    .Y(_11947_));
 sky130_fd_sc_hd__o211ai_2 _19310_ (.A1(_10926_),
    .A2(_11945_),
    .B1(_11946_),
    .C1(_11947_),
    .Y(_11948_));
 sky130_fd_sc_hd__a22oi_2 _19311_ (.A1(\cs_registers_i.mcycle_counter_i.counter[40] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][40] ),
    .Y(_11949_));
 sky130_fd_sc_hd__nor2_4 _19312_ (.A(_11225_),
    .B(_11949_),
    .Y(_11950_));
 sky130_fd_sc_hd__nand2_1 _19313_ (.A(\cs_registers_i.mscratch_q[8] ),
    .B(_11255_),
    .Y(_11951_));
 sky130_fd_sc_hd__a222oi_1 _19314_ (.A1(net92),
    .A2(_11238_),
    .B1(_11248_),
    .B2(\cs_registers_i.dcsr_q[8] ),
    .C1(\cs_registers_i.csr_depc_o[8] ),
    .C2(_11295_),
    .Y(_11952_));
 sky130_fd_sc_hd__a22oi_1 _19315_ (.A1(\cs_registers_i.csr_mepc_o[8] ),
    .A2(_11272_),
    .B1(_11270_),
    .B2(\cs_registers_i.mtval_q[8] ),
    .Y(_11953_));
 sky130_fd_sc_hd__nand3_2 _19316_ (.A(_11951_),
    .B(_11952_),
    .C(_11953_),
    .Y(_11954_));
 sky130_fd_sc_hd__nor3_4 _19317_ (.A(_11948_),
    .B(_11950_),
    .C(_11954_),
    .Y(_11955_));
 sky130_fd_sc_hd__nor3_1 _19318_ (.A(_09187_),
    .B(_11150_),
    .C(_11955_),
    .Y(_11956_));
 sky130_fd_sc_hd__a21oi_4 _19319_ (.A1(_09187_),
    .A2(_11148_),
    .B1(_11956_),
    .Y(_11957_));
 sky130_fd_sc_hd__nand2_1 _19320_ (.A(net273),
    .B(_11957_),
    .Y(_11958_));
 sky130_fd_sc_hd__o21ai_0 _19321_ (.A1(_11336_),
    .A2(_11944_),
    .B1(_11958_),
    .Y(_11959_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_667 ();
 sky130_fd_sc_hd__nand2_1 _19323_ (.A(_11335_),
    .B(_11937_),
    .Y(_11961_));
 sky130_fd_sc_hd__nand2_1 _19324_ (.A(_11320_),
    .B(_11961_),
    .Y(_11962_));
 sky130_fd_sc_hd__a21oi_1 _19325_ (.A1(net268),
    .A2(_11962_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[40] ),
    .Y(_11963_));
 sky130_fd_sc_hd__a21oi_1 _19326_ (.A1(net268),
    .A2(_11959_),
    .B1(_11963_),
    .Y(_00051_));
 sky130_fd_sc_hd__nand4_1 _19327_ (.A(\cs_registers_i.mcycle_counter_i.counter[40] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[41] ),
    .C(_11335_),
    .D(_11937_),
    .Y(_11964_));
 sky130_fd_sc_hd__a22oi_2 _19328_ (.A1(\cs_registers_i.mcycle_counter_i.counter[41] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][41] ),
    .Y(_11965_));
 sky130_fd_sc_hd__a22oi_2 _19329_ (.A1(\cs_registers_i.mcycle_counter_i.counter[9] ),
    .A2(_11264_),
    .B1(net285),
    .B2(\cs_registers_i.mhpmcounter[2][9] ),
    .Y(_11966_));
 sky130_fd_sc_hd__a222oi_1 _19330_ (.A1(\cs_registers_i.csr_mtvec_o[9] ),
    .A2(_10918_),
    .B1(_11252_),
    .B2(\cs_registers_i.dscratch0_q[9] ),
    .C1(\cs_registers_i.dscratch1_q[9] ),
    .C2(_11260_),
    .Y(_11967_));
 sky130_fd_sc_hd__o221ai_4 _19331_ (.A1(_11225_),
    .A2(_11965_),
    .B1(_11966_),
    .B2(_10926_),
    .C1(_11967_),
    .Y(_11968_));
 sky130_fd_sc_hd__a221o_1 _19332_ (.A1(net93),
    .A2(_11238_),
    .B1(_11295_),
    .B2(\cs_registers_i.csr_depc_o[9] ),
    .C1(_10907_),
    .X(_11969_));
 sky130_fd_sc_hd__a22o_1 _19333_ (.A1(\cs_registers_i.csr_mepc_o[9] ),
    .A2(_11272_),
    .B1(_11270_),
    .B2(\cs_registers_i.mtval_q[9] ),
    .X(_11970_));
 sky130_fd_sc_hd__a2111oi_4 _19334_ (.A1(\cs_registers_i.mscratch_q[9] ),
    .A2(_11255_),
    .B1(_11968_),
    .C1(_11969_),
    .D1(_11970_),
    .Y(_11971_));
 sky130_fd_sc_hd__nor3_1 _19335_ (.A(_09290_),
    .B(_11150_),
    .C(_11971_),
    .Y(_11972_));
 sky130_fd_sc_hd__a21oi_4 _19336_ (.A1(_09290_),
    .A2(_11148_),
    .B1(_11972_),
    .Y(_11973_));
 sky130_fd_sc_hd__nand2_1 _19337_ (.A(net273),
    .B(_11973_),
    .Y(_11974_));
 sky130_fd_sc_hd__o21ai_0 _19338_ (.A1(net273),
    .A2(_11964_),
    .B1(_11974_),
    .Y(_11975_));
 sky130_fd_sc_hd__o21ai_0 _19339_ (.A1(_11392_),
    .A2(_11944_),
    .B1(_11320_),
    .Y(_11976_));
 sky130_fd_sc_hd__a21oi_1 _19340_ (.A1(net268),
    .A2(_11976_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[41] ),
    .Y(_11977_));
 sky130_fd_sc_hd__a21oi_1 _19341_ (.A1(net268),
    .A2(_11975_),
    .B1(_11977_),
    .Y(_00052_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_666 ();
 sky130_fd_sc_hd__nand4_1 _19343_ (.A(\cs_registers_i.mcycle_counter_i.counter[39] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[40] ),
    .C(\cs_registers_i.mcycle_counter_i.counter[41] ),
    .D(\cs_registers_i.mcycle_counter_i.counter[42] ),
    .Y(_11979_));
 sky130_fd_sc_hd__nor2_2 _19344_ (.A(_11918_),
    .B(_11979_),
    .Y(_11980_));
 sky130_fd_sc_hd__nand2_1 _19345_ (.A(_11394_),
    .B(_11980_),
    .Y(_11981_));
 sky130_fd_sc_hd__o21ai_0 _19346_ (.A1(_11320_),
    .A2(_11357_),
    .B1(_11981_),
    .Y(_11982_));
 sky130_fd_sc_hd__nand3_1 _19347_ (.A(\cs_registers_i.mcycle_counter_i.counter[39] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[40] ),
    .C(\cs_registers_i.mcycle_counter_i.counter[41] ),
    .Y(_11983_));
 sky130_fd_sc_hd__o31ai_1 _19348_ (.A1(_11392_),
    .A2(_11918_),
    .A3(_11983_),
    .B1(_11320_),
    .Y(_11984_));
 sky130_fd_sc_hd__a21oi_1 _19349_ (.A1(net268),
    .A2(_11984_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[42] ),
    .Y(_11985_));
 sky130_fd_sc_hd__a21oi_1 _19350_ (.A1(net268),
    .A2(_11982_),
    .B1(_11985_),
    .Y(_00053_));
 sky130_fd_sc_hd__nand2_1 _19351_ (.A(\cs_registers_i.mcycle_counter_i.counter[43] ),
    .B(_11980_),
    .Y(_11986_));
 sky130_fd_sc_hd__o22ai_1 _19352_ (.A1(_11320_),
    .A2(_11391_),
    .B1(_11986_),
    .B2(_11336_),
    .Y(_11987_));
 sky130_fd_sc_hd__nand2_1 _19353_ (.A(_11335_),
    .B(_11980_),
    .Y(_11988_));
 sky130_fd_sc_hd__nand2_1 _19354_ (.A(_11320_),
    .B(_11988_),
    .Y(_11989_));
 sky130_fd_sc_hd__a21oi_1 _19355_ (.A1(net268),
    .A2(_11989_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[43] ),
    .Y(_11990_));
 sky130_fd_sc_hd__a21oi_1 _19356_ (.A1(net268),
    .A2(_11987_),
    .B1(_11990_),
    .Y(_00054_));
 sky130_fd_sc_hd__nand3_2 _19357_ (.A(\cs_registers_i.mcycle_counter_i.counter[44] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[43] ),
    .C(_11980_),
    .Y(_11991_));
 sky130_fd_sc_hd__o21ai_0 _19358_ (.A1(_11336_),
    .A2(_11991_),
    .B1(_11430_),
    .Y(_11992_));
 sky130_fd_sc_hd__o21ai_0 _19359_ (.A1(_11392_),
    .A2(_11986_),
    .B1(_11320_),
    .Y(_11993_));
 sky130_fd_sc_hd__a21oi_1 _19360_ (.A1(net268),
    .A2(_11993_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[44] ),
    .Y(_11994_));
 sky130_fd_sc_hd__a21oi_1 _19361_ (.A1(net268),
    .A2(_11992_),
    .B1(_11994_),
    .Y(_00055_));
 sky130_fd_sc_hd__nand4_1 _19362_ (.A(\cs_registers_i.mcycle_counter_i.counter[44] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[43] ),
    .C(\cs_registers_i.mcycle_counter_i.counter[45] ),
    .D(_11980_),
    .Y(_11995_));
 sky130_fd_sc_hd__o21ai_0 _19363_ (.A1(_11336_),
    .A2(_11995_),
    .B1(_11450_),
    .Y(_11996_));
 sky130_fd_sc_hd__o21ai_0 _19364_ (.A1(_11392_),
    .A2(_11991_),
    .B1(_11320_),
    .Y(_11997_));
 sky130_fd_sc_hd__a21oi_1 _19365_ (.A1(net268),
    .A2(_11997_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[45] ),
    .Y(_11998_));
 sky130_fd_sc_hd__a21oi_1 _19366_ (.A1(net268),
    .A2(_11996_),
    .B1(_11998_),
    .Y(_00056_));
 sky130_fd_sc_hd__nor2_1 _19367_ (.A(_11392_),
    .B(_11991_),
    .Y(_11999_));
 sky130_fd_sc_hd__nand3_1 _19368_ (.A(\cs_registers_i.mcycle_counter_i.counter[45] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[46] ),
    .C(_11999_),
    .Y(_12000_));
 sky130_fd_sc_hd__o21ai_0 _19369_ (.A1(net273),
    .A2(_12000_),
    .B1(_11467_),
    .Y(_12001_));
 sky130_fd_sc_hd__nand2_1 _19370_ (.A(\cs_registers_i.mcycle_counter_i.counter[45] ),
    .B(_11999_),
    .Y(_12002_));
 sky130_fd_sc_hd__nand2_1 _19371_ (.A(_11320_),
    .B(_12002_),
    .Y(_12003_));
 sky130_fd_sc_hd__a21oi_1 _19372_ (.A1(net268),
    .A2(_12003_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[46] ),
    .Y(_12004_));
 sky130_fd_sc_hd__a21oi_1 _19373_ (.A1(net268),
    .A2(_12001_),
    .B1(_12004_),
    .Y(_00057_));
 sky130_fd_sc_hd__nand2_1 _19374_ (.A(_11320_),
    .B(_12000_),
    .Y(_12005_));
 sky130_fd_sc_hd__a21oi_1 _19375_ (.A1(net268),
    .A2(_12005_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[47] ),
    .Y(_12006_));
 sky130_fd_sc_hd__or3b_1 _19376_ (.A(net273),
    .B(_12000_),
    .C_N(\cs_registers_i.mcycle_counter_i.counter[47] ),
    .X(_12007_));
 sky130_fd_sc_hd__a21boi_0 _19377_ (.A1(_11489_),
    .A2(_12007_),
    .B1_N(net268),
    .Y(_12008_));
 sky130_fd_sc_hd__nor2_1 _19378_ (.A(_12006_),
    .B(_12008_),
    .Y(_00058_));
 sky130_fd_sc_hd__nand4_1 _19379_ (.A(\cs_registers_i.mcycle_counter_i.counter[45] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[46] ),
    .C(\cs_registers_i.mcycle_counter_i.counter[47] ),
    .D(_11335_),
    .Y(_12009_));
 sky130_fd_sc_hd__nor2_1 _19380_ (.A(_11991_),
    .B(_12009_),
    .Y(_12010_));
 sky130_fd_sc_hd__o21ai_0 _19381_ (.A1(net273),
    .A2(_12010_),
    .B1(net268),
    .Y(_12011_));
 sky130_fd_sc_hd__nand2_1 _19382_ (.A(\cs_registers_i.mcycle_counter_i.counter[48] ),
    .B(_12011_),
    .Y(_12012_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_665 ();
 sky130_fd_sc_hd__o22ai_1 _19384_ (.A1(_11320_),
    .A2(_11505_),
    .B1(_12007_),
    .B2(\cs_registers_i.mcycle_counter_i.counter[48] ),
    .Y(_12014_));
 sky130_fd_sc_hd__nand2_1 _19385_ (.A(net268),
    .B(_12014_),
    .Y(_12015_));
 sky130_fd_sc_hd__nand2_1 _19386_ (.A(_12012_),
    .B(_12015_),
    .Y(_00059_));
 sky130_fd_sc_hd__inv_1 _19387_ (.A(\cs_registers_i.mcycle_counter_i.counter[48] ),
    .Y(_12016_));
 sky130_fd_sc_hd__inv_1 _19388_ (.A(\cs_registers_i.mcycle_counter_i.counter[44] ),
    .Y(_12017_));
 sky130_fd_sc_hd__inv_1 _19389_ (.A(\cs_registers_i.mcycle_counter_i.counter[43] ),
    .Y(_12018_));
 sky130_fd_sc_hd__nor4_1 _19390_ (.A(_11454_),
    .B(_11532_),
    .C(_11602_),
    .D(_11870_),
    .Y(_12019_));
 sky130_fd_sc_hd__nand4_1 _19391_ (.A(\cs_registers_i.mcycle_counter_i.counter[36] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[37] ),
    .C(\cs_registers_i.mcycle_counter_i.counter[38] ),
    .D(_12019_),
    .Y(_12020_));
 sky130_fd_sc_hd__or4_1 _19392_ (.A(_12017_),
    .B(_12018_),
    .C(_12020_),
    .D(_11979_),
    .X(_12021_));
 sky130_fd_sc_hd__nor3_2 _19393_ (.A(_12016_),
    .B(_12021_),
    .C(_12009_),
    .Y(_12022_));
 sky130_fd_sc_hd__o21ai_0 _19394_ (.A1(_11472_),
    .A2(_12022_),
    .B1(net268),
    .Y(_12023_));
 sky130_fd_sc_hd__nand2_1 _19395_ (.A(\cs_registers_i.mcycle_counter_i.counter[49] ),
    .B(_12023_),
    .Y(_12024_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_664 ();
 sky130_fd_sc_hd__nor2_1 _19397_ (.A(_11320_),
    .B(_11523_),
    .Y(_12026_));
 sky130_fd_sc_hd__nor3_1 _19398_ (.A(_12016_),
    .B(\cs_registers_i.mcycle_counter_i.counter[49] ),
    .C(_12007_),
    .Y(_12027_));
 sky130_fd_sc_hd__o21ai_0 _19399_ (.A1(_12026_),
    .A2(_12027_),
    .B1(net268),
    .Y(_12028_));
 sky130_fd_sc_hd__nand2_1 _19400_ (.A(_12024_),
    .B(_12028_),
    .Y(_00060_));
 sky130_fd_sc_hd__a21boi_0 _19401_ (.A1(\cs_registers_i.mcycle_counter_i.counter[4] ),
    .A2(_11394_),
    .B1_N(_11888_),
    .Y(_12029_));
 sky130_fd_sc_hd__a21oi_1 _19402_ (.A1(_11320_),
    .A2(_11392_),
    .B1(_11330_),
    .Y(_12030_));
 sky130_fd_sc_hd__o22a_1 _19403_ (.A1(_11330_),
    .A2(_12029_),
    .B1(_12030_),
    .B2(\cs_registers_i.mcycle_counter_i.counter[4] ),
    .X(_00061_));
 sky130_fd_sc_hd__nand3_1 _19404_ (.A(\cs_registers_i.mcycle_counter_i.counter[49] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[50] ),
    .C(_12022_),
    .Y(_12031_));
 sky130_fd_sc_hd__o21ai_0 _19405_ (.A1(_11472_),
    .A2(_12031_),
    .B1(_11548_),
    .Y(_12032_));
 sky130_fd_sc_hd__nand2_1 _19406_ (.A(\cs_registers_i.mcycle_counter_i.counter[49] ),
    .B(_12022_),
    .Y(_12033_));
 sky130_fd_sc_hd__nand2_1 _19407_ (.A(_11316_),
    .B(_12033_),
    .Y(_12034_));
 sky130_fd_sc_hd__a21oi_1 _19408_ (.A1(_11833_),
    .A2(_12034_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[50] ),
    .Y(_12035_));
 sky130_fd_sc_hd__a21oi_1 _19409_ (.A1(_11833_),
    .A2(_12032_),
    .B1(_12035_),
    .Y(_00062_));
 sky130_fd_sc_hd__and3_1 _19410_ (.A(\cs_registers_i.mcycle_counter_i.counter[49] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[50] ),
    .C(_12022_),
    .X(_12036_));
 sky130_fd_sc_hd__nand2_1 _19411_ (.A(\cs_registers_i.mcycle_counter_i.counter[51] ),
    .B(_12036_),
    .Y(_12037_));
 sky130_fd_sc_hd__o21ai_0 _19412_ (.A1(_11472_),
    .A2(_12037_),
    .B1(_11565_),
    .Y(_12038_));
 sky130_fd_sc_hd__nand2_1 _19413_ (.A(_11316_),
    .B(_12031_),
    .Y(_12039_));
 sky130_fd_sc_hd__a21oi_1 _19414_ (.A1(_11833_),
    .A2(_12039_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[51] ),
    .Y(_12040_));
 sky130_fd_sc_hd__a21oi_1 _19415_ (.A1(_11833_),
    .A2(_12038_),
    .B1(_12040_),
    .Y(_00063_));
 sky130_fd_sc_hd__and2_0 _19416_ (.A(\cs_registers_i.mcycle_counter_i.counter[51] ),
    .B(_12036_),
    .X(_12041_));
 sky130_fd_sc_hd__nand2_1 _19417_ (.A(\cs_registers_i.mcycle_counter_i.counter[52] ),
    .B(_12041_),
    .Y(_12042_));
 sky130_fd_sc_hd__o21ai_0 _19418_ (.A1(_11472_),
    .A2(_12042_),
    .B1(_11601_),
    .Y(_12043_));
 sky130_fd_sc_hd__nand2_1 _19419_ (.A(_11316_),
    .B(_12037_),
    .Y(_12044_));
 sky130_fd_sc_hd__a21oi_1 _19420_ (.A1(_11833_),
    .A2(_12044_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[52] ),
    .Y(_12045_));
 sky130_fd_sc_hd__a21oi_1 _19421_ (.A1(_11833_),
    .A2(_12043_),
    .B1(_12045_),
    .Y(_00064_));
 sky130_fd_sc_hd__nand3_1 _19422_ (.A(\cs_registers_i.mcycle_counter_i.counter[52] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[53] ),
    .C(_12041_),
    .Y(_12046_));
 sky130_fd_sc_hd__nand2_1 _19423_ (.A(_11472_),
    .B(_11623_),
    .Y(_12047_));
 sky130_fd_sc_hd__o21ai_0 _19424_ (.A1(_11472_),
    .A2(_12046_),
    .B1(_12047_),
    .Y(_12048_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_663 ();
 sky130_fd_sc_hd__nand2_1 _19426_ (.A(_11316_),
    .B(_12042_),
    .Y(_12050_));
 sky130_fd_sc_hd__a21oi_1 _19427_ (.A1(_11833_),
    .A2(_12050_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[53] ),
    .Y(_12051_));
 sky130_fd_sc_hd__a21oi_1 _19428_ (.A1(_11833_),
    .A2(_12048_),
    .B1(_12051_),
    .Y(_00065_));
 sky130_fd_sc_hd__and3_1 _19429_ (.A(\cs_registers_i.mcycle_counter_i.counter[52] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[53] ),
    .C(_12041_),
    .X(_12052_));
 sky130_fd_sc_hd__nand2_1 _19430_ (.A(\cs_registers_i.mcycle_counter_i.counter[54] ),
    .B(_12052_),
    .Y(_12053_));
 sky130_fd_sc_hd__o21ai_0 _19431_ (.A1(_11472_),
    .A2(_12053_),
    .B1(_11645_),
    .Y(_12054_));
 sky130_fd_sc_hd__nand2_1 _19432_ (.A(_11316_),
    .B(_12046_),
    .Y(_12055_));
 sky130_fd_sc_hd__a21oi_1 _19433_ (.A1(_11833_),
    .A2(_12055_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[54] ),
    .Y(_12056_));
 sky130_fd_sc_hd__a21oi_1 _19434_ (.A1(_11833_),
    .A2(_12054_),
    .B1(_12056_),
    .Y(_00066_));
 sky130_fd_sc_hd__nand3_1 _19435_ (.A(\cs_registers_i.mcycle_counter_i.counter[54] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[55] ),
    .C(_12052_),
    .Y(_12057_));
 sky130_fd_sc_hd__nand2_1 _19436_ (.A(_11472_),
    .B(_11664_),
    .Y(_12058_));
 sky130_fd_sc_hd__o21ai_0 _19437_ (.A1(_11472_),
    .A2(_12057_),
    .B1(_12058_),
    .Y(_12059_));
 sky130_fd_sc_hd__nand2_1 _19438_ (.A(_11316_),
    .B(_12053_),
    .Y(_12060_));
 sky130_fd_sc_hd__a21oi_1 _19439_ (.A1(_11833_),
    .A2(_12060_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[55] ),
    .Y(_12061_));
 sky130_fd_sc_hd__a21oi_1 _19440_ (.A1(_11833_),
    .A2(_12059_),
    .B1(_12061_),
    .Y(_00067_));
 sky130_fd_sc_hd__and3_1 _19441_ (.A(\cs_registers_i.mcycle_counter_i.counter[54] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[55] ),
    .C(_12052_),
    .X(_12062_));
 sky130_fd_sc_hd__nand2_1 _19442_ (.A(\cs_registers_i.mcycle_counter_i.counter[56] ),
    .B(_12062_),
    .Y(_12063_));
 sky130_fd_sc_hd__nand2_1 _19443_ (.A(_11472_),
    .B(_11684_),
    .Y(_12064_));
 sky130_fd_sc_hd__o21ai_0 _19444_ (.A1(_11472_),
    .A2(_12063_),
    .B1(_12064_),
    .Y(_12065_));
 sky130_fd_sc_hd__nand2_1 _19445_ (.A(_11316_),
    .B(_12057_),
    .Y(_12066_));
 sky130_fd_sc_hd__a21oi_1 _19446_ (.A1(_11833_),
    .A2(_12066_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[56] ),
    .Y(_12067_));
 sky130_fd_sc_hd__a21oi_1 _19447_ (.A1(_11833_),
    .A2(_12065_),
    .B1(_12067_),
    .Y(_00068_));
 sky130_fd_sc_hd__nand3_1 _19448_ (.A(\cs_registers_i.mcycle_counter_i.counter[56] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[57] ),
    .C(_12062_),
    .Y(_12068_));
 sky130_fd_sc_hd__nand2_1 _19449_ (.A(_11472_),
    .B(_11706_),
    .Y(_12069_));
 sky130_fd_sc_hd__o21ai_0 _19450_ (.A1(_11472_),
    .A2(_12068_),
    .B1(_12069_),
    .Y(_12070_));
 sky130_fd_sc_hd__nand2_1 _19451_ (.A(_11316_),
    .B(_12063_),
    .Y(_12071_));
 sky130_fd_sc_hd__a21oi_1 _19452_ (.A1(_11833_),
    .A2(_12071_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[57] ),
    .Y(_12072_));
 sky130_fd_sc_hd__a21oi_1 _19453_ (.A1(_11833_),
    .A2(_12070_),
    .B1(_12072_),
    .Y(_00069_));
 sky130_fd_sc_hd__nand4_1 _19454_ (.A(\cs_registers_i.mcycle_counter_i.counter[56] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[57] ),
    .C(\cs_registers_i.mcycle_counter_i.counter[58] ),
    .D(_12062_),
    .Y(_12073_));
 sky130_fd_sc_hd__nand2_1 _19455_ (.A(_11472_),
    .B(_11726_),
    .Y(_12074_));
 sky130_fd_sc_hd__o21ai_0 _19456_ (.A1(_11472_),
    .A2(_12073_),
    .B1(_12074_),
    .Y(_12075_));
 sky130_fd_sc_hd__nand2_1 _19457_ (.A(_11316_),
    .B(_12068_),
    .Y(_12076_));
 sky130_fd_sc_hd__a21oi_1 _19458_ (.A1(_11833_),
    .A2(_12076_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[58] ),
    .Y(_12077_));
 sky130_fd_sc_hd__a21oi_1 _19459_ (.A1(_11833_),
    .A2(_12075_),
    .B1(_12077_),
    .Y(_00070_));
 sky130_fd_sc_hd__and4_1 _19460_ (.A(\cs_registers_i.mcycle_counter_i.counter[48] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[49] ),
    .C(\cs_registers_i.mcycle_counter_i.counter[50] ),
    .D(_12010_),
    .X(_12078_));
 sky130_fd_sc_hd__and4_1 _19461_ (.A(\cs_registers_i.mcycle_counter_i.counter[51] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[52] ),
    .C(\cs_registers_i.mcycle_counter_i.counter[53] ),
    .D(_12078_),
    .X(_12079_));
 sky130_fd_sc_hd__and4_1 _19462_ (.A(\cs_registers_i.mcycle_counter_i.counter[54] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[55] ),
    .C(\cs_registers_i.mcycle_counter_i.counter[56] ),
    .D(_12079_),
    .X(_12080_));
 sky130_fd_sc_hd__and4_1 _19463_ (.A(\cs_registers_i.mcycle_counter_i.counter[57] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[58] ),
    .C(\cs_registers_i.mcycle_counter_i.counter[59] ),
    .D(_12080_),
    .X(_12081_));
 sky130_fd_sc_hd__nand2_1 _19464_ (.A(_11320_),
    .B(_12081_),
    .Y(_12082_));
 sky130_fd_sc_hd__nand2_1 _19465_ (.A(_11748_),
    .B(_12082_),
    .Y(_12083_));
 sky130_fd_sc_hd__nand2_1 _19466_ (.A(_11316_),
    .B(_12073_),
    .Y(_12084_));
 sky130_fd_sc_hd__a21oi_1 _19467_ (.A1(_11833_),
    .A2(_12084_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[59] ),
    .Y(_12085_));
 sky130_fd_sc_hd__a21oi_1 _19468_ (.A1(_11833_),
    .A2(_12083_),
    .B1(_12085_),
    .Y(_00071_));
 sky130_fd_sc_hd__nand3_1 _19469_ (.A(\cs_registers_i.mcycle_counter_i.counter[4] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[5] ),
    .C(_11394_),
    .Y(_12086_));
 sky130_fd_sc_hd__o21ai_0 _19470_ (.A1(_11316_),
    .A2(_11902_),
    .B1(_12086_),
    .Y(_12087_));
 sky130_fd_sc_hd__nand2_1 _19471_ (.A(\cs_registers_i.mcycle_counter_i.counter[4] ),
    .B(_11335_),
    .Y(_12088_));
 sky130_fd_sc_hd__nand2_1 _19472_ (.A(_11320_),
    .B(_12088_),
    .Y(_12089_));
 sky130_fd_sc_hd__a21oi_1 _19473_ (.A1(_11322_),
    .A2(_12089_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[5] ),
    .Y(_12090_));
 sky130_fd_sc_hd__a21oi_1 _19474_ (.A1(_11322_),
    .A2(_12087_),
    .B1(_12090_),
    .Y(_00072_));
 sky130_fd_sc_hd__inv_1 _19475_ (.A(\cs_registers_i.mcycle_counter_i.counter[60] ),
    .Y(_12091_));
 sky130_fd_sc_hd__o21ai_0 _19476_ (.A1(_11328_),
    .A2(_12081_),
    .B1(_11833_),
    .Y(_12092_));
 sky130_fd_sc_hd__nand2_1 _19477_ (.A(\cs_registers_i.mcycle_counter_i.counter[60] ),
    .B(_12081_),
    .Y(_12093_));
 sky130_fd_sc_hd__o21ai_0 _19478_ (.A1(_11328_),
    .A2(_12093_),
    .B1(_11767_),
    .Y(_12094_));
 sky130_fd_sc_hd__a22oi_1 _19479_ (.A1(_12091_),
    .A2(_12092_),
    .B1(_12094_),
    .B2(_11833_),
    .Y(_00073_));
 sky130_fd_sc_hd__nand3_1 _19480_ (.A(\cs_registers_i.mcycle_counter_i.counter[60] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[61] ),
    .C(_12081_),
    .Y(_12095_));
 sky130_fd_sc_hd__o21ai_0 _19481_ (.A1(_11328_),
    .A2(_12095_),
    .B1(_11787_),
    .Y(_12096_));
 sky130_fd_sc_hd__nand2_1 _19482_ (.A(_11320_),
    .B(_12093_),
    .Y(_12097_));
 sky130_fd_sc_hd__a21oi_1 _19483_ (.A1(_11833_),
    .A2(_12097_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[61] ),
    .Y(_12098_));
 sky130_fd_sc_hd__a21oi_1 _19484_ (.A1(_11833_),
    .A2(_12096_),
    .B1(_12098_),
    .Y(_00074_));
 sky130_fd_sc_hd__inv_1 _19485_ (.A(_12095_),
    .Y(_12099_));
 sky130_fd_sc_hd__nand2_1 _19486_ (.A(\cs_registers_i.mcycle_counter_i.counter[62] ),
    .B(_12099_),
    .Y(_12100_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_662 ();
 sky130_fd_sc_hd__nand2_1 _19488_ (.A(_11328_),
    .B(_11808_),
    .Y(_12102_));
 sky130_fd_sc_hd__o21ai_0 _19489_ (.A1(_11328_),
    .A2(_12100_),
    .B1(_12102_),
    .Y(_12103_));
 sky130_fd_sc_hd__nand2_1 _19490_ (.A(_11320_),
    .B(_12095_),
    .Y(_12104_));
 sky130_fd_sc_hd__a21oi_1 _19491_ (.A1(_11833_),
    .A2(_12104_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[62] ),
    .Y(_12105_));
 sky130_fd_sc_hd__a21oi_1 _19492_ (.A1(_11833_),
    .A2(_12103_),
    .B1(_12105_),
    .Y(_00075_));
 sky130_fd_sc_hd__o31ai_4 _19493_ (.A1(_10695_),
    .A2(_11150_),
    .A3(_11824_),
    .B1(_11825_),
    .Y(_12106_));
 sky130_fd_sc_hd__nand4_1 _19494_ (.A(\cs_registers_i.mcycle_counter_i.counter[62] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[63] ),
    .C(_11320_),
    .D(_12099_),
    .Y(_12107_));
 sky130_fd_sc_hd__o21ai_0 _19495_ (.A1(_11320_),
    .A2(_12106_),
    .B1(_12107_),
    .Y(_12108_));
 sky130_fd_sc_hd__nand2_1 _19496_ (.A(_11320_),
    .B(_12100_),
    .Y(_12109_));
 sky130_fd_sc_hd__a21oi_1 _19497_ (.A1(_11833_),
    .A2(_12109_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[63] ),
    .Y(_12110_));
 sky130_fd_sc_hd__a21oi_1 _19498_ (.A1(_11833_),
    .A2(_12108_),
    .B1(_12110_),
    .Y(_00076_));
 sky130_fd_sc_hd__nand3_1 _19499_ (.A(\cs_registers_i.mcycle_counter_i.counter[4] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[5] ),
    .C(_11335_),
    .Y(_12111_));
 sky130_fd_sc_hd__a21oi_1 _19500_ (.A1(_11320_),
    .A2(_12111_),
    .B1(_11330_),
    .Y(_12112_));
 sky130_fd_sc_hd__o31a_4 _19501_ (.A1(_08547_),
    .A2(_11150_),
    .A3(_11915_),
    .B1(_11916_),
    .X(_12113_));
 sky130_fd_sc_hd__a22oi_1 _19502_ (.A1(_11337_),
    .A2(_11394_),
    .B1(_12113_),
    .B2(_11472_),
    .Y(_12114_));
 sky130_fd_sc_hd__o22a_1 _19503_ (.A1(\cs_registers_i.mcycle_counter_i.counter[6] ),
    .A2(_12112_),
    .B1(_12114_),
    .B2(_11330_),
    .X(_00077_));
 sky130_fd_sc_hd__a21oi_1 _19504_ (.A1(_11335_),
    .A2(_11337_),
    .B1(net273),
    .Y(_12115_));
 sky130_fd_sc_hd__nor2_1 _19505_ (.A(_11330_),
    .B(_12115_),
    .Y(_12116_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_661 ();
 sky130_fd_sc_hd__and3_1 _19507_ (.A(\cs_registers_i.mcycle_counter_i.counter[7] ),
    .B(_11337_),
    .C(_11394_),
    .X(_12118_));
 sky130_fd_sc_hd__a21oi_1 _19508_ (.A1(_11472_),
    .A2(_11935_),
    .B1(_12118_),
    .Y(_12119_));
 sky130_fd_sc_hd__o22a_1 _19509_ (.A1(\cs_registers_i.mcycle_counter_i.counter[7] ),
    .A2(_12116_),
    .B1(_12119_),
    .B2(_11330_),
    .X(_00078_));
 sky130_fd_sc_hd__nand3_1 _19510_ (.A(\cs_registers_i.mcycle_counter_i.counter[7] ),
    .B(_11335_),
    .C(_11337_),
    .Y(_12120_));
 sky130_fd_sc_hd__a21oi_1 _19511_ (.A1(_11320_),
    .A2(_12120_),
    .B1(_11330_),
    .Y(_12121_));
 sky130_fd_sc_hd__a21boi_0 _19512_ (.A1(_11338_),
    .A2(_11394_),
    .B1_N(_11958_),
    .Y(_12122_));
 sky130_fd_sc_hd__o22a_1 _19513_ (.A1(\cs_registers_i.mcycle_counter_i.counter[8] ),
    .A2(_12121_),
    .B1(_12122_),
    .B2(_11330_),
    .X(_00079_));
 sky130_fd_sc_hd__nand2_1 _19514_ (.A(_11335_),
    .B(_11338_),
    .Y(_12123_));
 sky130_fd_sc_hd__nand2_1 _19515_ (.A(_11320_),
    .B(_12123_),
    .Y(_12124_));
 sky130_fd_sc_hd__a21oi_1 _19516_ (.A1(_11322_),
    .A2(_12124_),
    .B1(\cs_registers_i.mcycle_counter_i.counter[9] ),
    .Y(_12125_));
 sky130_fd_sc_hd__nand4_1 _19517_ (.A(\cs_registers_i.mcycle_counter_i.counter[9] ),
    .B(_11320_),
    .C(_11335_),
    .D(_11338_),
    .Y(_12126_));
 sky130_fd_sc_hd__a21oi_1 _19518_ (.A1(_11974_),
    .A2(_12126_),
    .B1(_11330_),
    .Y(_12127_));
 sky130_fd_sc_hd__nor2_1 _19519_ (.A(_12125_),
    .B(_12127_),
    .Y(_00080_));
 sky130_fd_sc_hd__nand2_4 _19520_ (.A(_08269_),
    .B(_10931_),
    .Y(_12128_));
 sky130_fd_sc_hd__nor4_4 _19521_ (.A(\cs_registers_i.mcountinhibit[2] ),
    .B(_10850_),
    .C(_10947_),
    .D(_12128_),
    .Y(_12129_));
 sky130_fd_sc_hd__nand2_8 _19522_ (.A(_11200_),
    .B(_12129_),
    .Y(_12130_));
 sky130_fd_sc_hd__nor3b_4 _19523_ (.A(_11325_),
    .B(_11313_),
    .C_N(_11267_),
    .Y(_12131_));
 sky130_fd_sc_hd__nand2_2 _19524_ (.A(_11314_),
    .B(_11267_),
    .Y(_12132_));
 sky130_fd_sc_hd__nor2_8 _19525_ (.A(_11325_),
    .B(_12132_),
    .Y(_12133_));
 sky130_fd_sc_hd__nand2_8 _19526_ (.A(_10928_),
    .B(_12133_),
    .Y(_12134_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_660 ();
 sky130_fd_sc_hd__o21ai_4 _19528_ (.A1(_12130_),
    .A2(_12131_),
    .B1(_12134_),
    .Y(_12136_));
 sky130_fd_sc_hd__nor2_2 _19529_ (.A(_12130_),
    .B(_12133_),
    .Y(_12137_));
 sky130_fd_sc_hd__nand2_1 _19530_ (.A(\cs_registers_i.mhpmcounter[2][0] ),
    .B(_12137_),
    .Y(_12138_));
 sky130_fd_sc_hd__nand3b_4 _19531_ (.A_N(_11313_),
    .B(_11267_),
    .C(_10929_),
    .Y(_12139_));
 sky130_fd_sc_hd__a21oi_4 _19532_ (.A1(_10925_),
    .A2(_10927_),
    .B1(_12139_),
    .Y(_12140_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_658 ();
 sky130_fd_sc_hd__nand2_1 _19535_ (.A(_11280_),
    .B(_12140_),
    .Y(_12143_));
 sky130_fd_sc_hd__o211a_1 _19536_ (.A1(\cs_registers_i.mhpmcounter[2][0] ),
    .A2(_12136_),
    .B1(_12138_),
    .C1(_12143_),
    .X(_00081_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_656 ();
 sky130_fd_sc_hd__and3_1 _19539_ (.A(\cs_registers_i.mhpmcounter[2][0] ),
    .B(\cs_registers_i.mhpmcounter[2][1] ),
    .C(\cs_registers_i.mhpmcounter[2][2] ),
    .X(_12146_));
 sky130_fd_sc_hd__nand2_4 _19540_ (.A(\cs_registers_i.mhpmcounter[2][3] ),
    .B(_12146_),
    .Y(_12147_));
 sky130_fd_sc_hd__nor2_4 _19541_ (.A(net272),
    .B(_12147_),
    .Y(_12148_));
 sky130_fd_sc_hd__and3_1 _19542_ (.A(\cs_registers_i.mhpmcounter[2][4] ),
    .B(\cs_registers_i.mhpmcounter[2][5] ),
    .C(\cs_registers_i.mhpmcounter[2][6] ),
    .X(_12149_));
 sky130_fd_sc_hd__and4_1 _19543_ (.A(\cs_registers_i.mhpmcounter[2][7] ),
    .B(\cs_registers_i.mhpmcounter[2][8] ),
    .C(\cs_registers_i.mhpmcounter[2][9] ),
    .D(_12149_),
    .X(_12150_));
 sky130_fd_sc_hd__and2_0 _19544_ (.A(\cs_registers_i.mhpmcounter[2][10] ),
    .B(_12150_),
    .X(_12151_));
 sky130_fd_sc_hd__nand2_1 _19545_ (.A(_12148_),
    .B(_12151_),
    .Y(_12152_));
 sky130_fd_sc_hd__o21ai_0 _19546_ (.A1(_11357_),
    .A2(_12139_),
    .B1(_12152_),
    .Y(_12153_));
 sky130_fd_sc_hd__and2_1 _19547_ (.A(\cs_registers_i.mhpmcounter[2][3] ),
    .B(_12146_),
    .X(_12154_));
 sky130_fd_sc_hd__nand2_2 _19548_ (.A(_12139_),
    .B(_12154_),
    .Y(_12155_));
 sky130_fd_sc_hd__nor2_8 _19549_ (.A(_12155_),
    .B(_12130_),
    .Y(_12156_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_655 ();
 sky130_fd_sc_hd__a211oi_1 _19551_ (.A1(_12150_),
    .A2(_12156_),
    .B1(\cs_registers_i.mhpmcounter[2][10] ),
    .C1(_12140_),
    .Y(_12158_));
 sky130_fd_sc_hd__a21oi_1 _19552_ (.A1(_12136_),
    .A2(_12153_),
    .B1(_12158_),
    .Y(_00082_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_654 ();
 sky130_fd_sc_hd__a211oi_1 _19554_ (.A1(_12156_),
    .A2(_12151_),
    .B1(\cs_registers_i.mhpmcounter[2][11] ),
    .C1(_12140_),
    .Y(_12160_));
 sky130_fd_sc_hd__nand2_8 _19555_ (.A(_10928_),
    .B(net272),
    .Y(_12161_));
 sky130_fd_sc_hd__nand3_1 _19556_ (.A(\cs_registers_i.mhpmcounter[2][11] ),
    .B(_12156_),
    .C(_12151_),
    .Y(_12162_));
 sky130_fd_sc_hd__o21ai_0 _19557_ (.A1(_11391_),
    .A2(_12161_),
    .B1(_12162_),
    .Y(_12163_));
 sky130_fd_sc_hd__nor2_1 _19558_ (.A(_12160_),
    .B(_12163_),
    .Y(_00083_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_653 ();
 sky130_fd_sc_hd__and3_2 _19560_ (.A(\cs_registers_i.mhpmcounter[2][11] ),
    .B(\cs_registers_i.mhpmcounter[2][10] ),
    .C(_12150_),
    .X(_12165_));
 sky130_fd_sc_hd__nand2_1 _19561_ (.A(_12156_),
    .B(_12165_),
    .Y(_12166_));
 sky130_fd_sc_hd__nand3_1 _19562_ (.A(\cs_registers_i.mhpmcounter[2][12] ),
    .B(_12161_),
    .C(_12166_),
    .Y(_12167_));
 sky130_fd_sc_hd__o221ai_1 _19563_ (.A1(_11428_),
    .A2(_12161_),
    .B1(_12166_),
    .B2(\cs_registers_i.mhpmcounter[2][12] ),
    .C1(_12167_),
    .Y(_00084_));
 sky130_fd_sc_hd__nand3_1 _19564_ (.A(\cs_registers_i.mhpmcounter[2][12] ),
    .B(_12156_),
    .C(_12165_),
    .Y(_12168_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_652 ();
 sky130_fd_sc_hd__nand2_1 _19566_ (.A(_11448_),
    .B(_12140_),
    .Y(_12170_));
 sky130_fd_sc_hd__o211ai_1 _19567_ (.A1(\cs_registers_i.mhpmcounter[2][13] ),
    .A2(_12140_),
    .B1(_12168_),
    .C1(_12170_),
    .Y(_12171_));
 sky130_fd_sc_hd__o21ai_0 _19568_ (.A1(\cs_registers_i.mhpmcounter[2][13] ),
    .A2(_12168_),
    .B1(_12171_),
    .Y(_00085_));
 sky130_fd_sc_hd__nor2_1 _19569_ (.A(\cs_registers_i.mhpmcounter[2][14] ),
    .B(_12140_),
    .Y(_12172_));
 sky130_fd_sc_hd__nand4_1 _19570_ (.A(\cs_registers_i.mhpmcounter[2][12] ),
    .B(\cs_registers_i.mhpmcounter[2][13] ),
    .C(_12156_),
    .D(_12165_),
    .Y(_12173_));
 sky130_fd_sc_hd__mux2_1 _19571_ (.A0(\cs_registers_i.mhpmcounter[2][14] ),
    .A1(_12172_),
    .S(_12173_),
    .X(_12174_));
 sky130_fd_sc_hd__a21oi_1 _19572_ (.A1(_11465_),
    .A2(_12140_),
    .B1(_12174_),
    .Y(_00086_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_651 ();
 sky130_fd_sc_hd__nand2_1 _19574_ (.A(\cs_registers_i.mhpmcounter[2][15] ),
    .B(_12134_),
    .Y(_12176_));
 sky130_fd_sc_hd__and3_1 _19575_ (.A(\cs_registers_i.mhpmcounter[2][12] ),
    .B(\cs_registers_i.mhpmcounter[2][13] ),
    .C(\cs_registers_i.mhpmcounter[2][14] ),
    .X(_12177_));
 sky130_fd_sc_hd__nand3_1 _19576_ (.A(_12156_),
    .B(_12165_),
    .C(_12177_),
    .Y(_12178_));
 sky130_fd_sc_hd__mux2_1 _19577_ (.A0(\cs_registers_i.mhpmcounter[2][15] ),
    .A1(_12176_),
    .S(_12178_),
    .X(_12179_));
 sky130_fd_sc_hd__o21ai_0 _19578_ (.A1(_11488_),
    .A2(_12134_),
    .B1(_12179_),
    .Y(_00087_));
 sky130_fd_sc_hd__and3_1 _19579_ (.A(\cs_registers_i.mhpmcounter[2][15] ),
    .B(_12165_),
    .C(_12177_),
    .X(_12180_));
 sky130_fd_sc_hd__nand2_1 _19580_ (.A(_12156_),
    .B(_12180_),
    .Y(_12181_));
 sky130_fd_sc_hd__o22ai_1 _19581_ (.A1(_11505_),
    .A2(_12161_),
    .B1(_12181_),
    .B2(\cs_registers_i.mhpmcounter[2][16] ),
    .Y(_12182_));
 sky130_fd_sc_hd__a31o_1 _19582_ (.A1(\cs_registers_i.mhpmcounter[2][16] ),
    .A2(_12161_),
    .A3(_12181_),
    .B1(_12182_),
    .X(_00088_));
 sky130_fd_sc_hd__and2_1 _19583_ (.A(\cs_registers_i.mhpmcounter[2][16] ),
    .B(_12180_),
    .X(_12183_));
 sky130_fd_sc_hd__a211oi_1 _19584_ (.A1(_12156_),
    .A2(_12183_),
    .B1(\cs_registers_i.mhpmcounter[2][17] ),
    .C1(_12140_),
    .Y(_12184_));
 sky130_fd_sc_hd__nand3_1 _19585_ (.A(\cs_registers_i.mhpmcounter[2][17] ),
    .B(_12156_),
    .C(_12183_),
    .Y(_12185_));
 sky130_fd_sc_hd__nand2_1 _19586_ (.A(_11523_),
    .B(_12140_),
    .Y(_12186_));
 sky130_fd_sc_hd__nand2_1 _19587_ (.A(_12185_),
    .B(_12186_),
    .Y(_12187_));
 sky130_fd_sc_hd__nor2_1 _19588_ (.A(_12184_),
    .B(_12187_),
    .Y(_00089_));
 sky130_fd_sc_hd__nand3_1 _19589_ (.A(\cs_registers_i.mhpmcounter[2][18] ),
    .B(_12134_),
    .C(_12185_),
    .Y(_12188_));
 sky130_fd_sc_hd__o221ai_1 _19590_ (.A1(_11546_),
    .A2(_12161_),
    .B1(_12185_),
    .B2(\cs_registers_i.mhpmcounter[2][18] ),
    .C1(_12188_),
    .Y(_00090_));
 sky130_fd_sc_hd__nand4_1 _19591_ (.A(\cs_registers_i.mhpmcounter[2][17] ),
    .B(\cs_registers_i.mhpmcounter[2][18] ),
    .C(_12156_),
    .D(_12183_),
    .Y(_12189_));
 sky130_fd_sc_hd__nand3_1 _19592_ (.A(\cs_registers_i.mhpmcounter[2][19] ),
    .B(_12134_),
    .C(_12189_),
    .Y(_12190_));
 sky130_fd_sc_hd__or2_0 _19593_ (.A(\cs_registers_i.mhpmcounter[2][19] ),
    .B(_12189_),
    .X(_12191_));
 sky130_fd_sc_hd__o211ai_1 _19594_ (.A1(_11563_),
    .A2(_12134_),
    .B1(_12190_),
    .C1(_12191_),
    .Y(_00091_));
 sky130_fd_sc_hd__nand3_1 _19595_ (.A(\cs_registers_i.mhpmcounter[2][1] ),
    .B(_12161_),
    .C(_12138_),
    .Y(_12192_));
 sky130_fd_sc_hd__o221ai_1 _19596_ (.A1(_11582_),
    .A2(_12161_),
    .B1(_12138_),
    .B2(\cs_registers_i.mhpmcounter[2][1] ),
    .C1(_12192_),
    .Y(_00092_));
 sky130_fd_sc_hd__and4_1 _19597_ (.A(\cs_registers_i.mhpmcounter[2][17] ),
    .B(\cs_registers_i.mhpmcounter[2][18] ),
    .C(\cs_registers_i.mhpmcounter[2][19] ),
    .D(_12183_),
    .X(_12193_));
 sky130_fd_sc_hd__and3_1 _19598_ (.A(\cs_registers_i.mhpmcounter[2][20] ),
    .B(_12156_),
    .C(_12193_),
    .X(_12194_));
 sky130_fd_sc_hd__a211oi_1 _19599_ (.A1(_12156_),
    .A2(_12193_),
    .B1(\cs_registers_i.mhpmcounter[2][20] ),
    .C1(_12140_),
    .Y(_12195_));
 sky130_fd_sc_hd__a211oi_1 _19600_ (.A1(_11599_),
    .A2(_12140_),
    .B1(_12194_),
    .C1(_12195_),
    .Y(_00093_));
 sky130_fd_sc_hd__and3_1 _19601_ (.A(\cs_registers_i.mhpmcounter[2][20] ),
    .B(\cs_registers_i.mhpmcounter[2][21] ),
    .C(_12193_),
    .X(_12196_));
 sky130_fd_sc_hd__nand2_1 _19602_ (.A(_12148_),
    .B(_12196_),
    .Y(_12197_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_650 ();
 sky130_fd_sc_hd__nand2_1 _19604_ (.A(_11623_),
    .B(net272),
    .Y(_12199_));
 sky130_fd_sc_hd__nand2_1 _19605_ (.A(_12197_),
    .B(_12199_),
    .Y(_12200_));
 sky130_fd_sc_hd__nor3_1 _19606_ (.A(\cs_registers_i.mhpmcounter[2][21] ),
    .B(_12140_),
    .C(_12194_),
    .Y(_12201_));
 sky130_fd_sc_hd__a21oi_1 _19607_ (.A1(_12136_),
    .A2(_12200_),
    .B1(_12201_),
    .Y(_00094_));
 sky130_fd_sc_hd__nand2_1 _19608_ (.A(_12156_),
    .B(_12196_),
    .Y(_12202_));
 sky130_fd_sc_hd__nor2_1 _19609_ (.A(\cs_registers_i.mhpmcounter[2][22] ),
    .B(_12202_),
    .Y(_12203_));
 sky130_fd_sc_hd__a31oi_1 _19610_ (.A1(\cs_registers_i.mhpmcounter[2][22] ),
    .A2(_12134_),
    .A3(_12202_),
    .B1(_12203_),
    .Y(_12204_));
 sky130_fd_sc_hd__o21ai_0 _19611_ (.A1(_11643_),
    .A2(_12134_),
    .B1(_12204_),
    .Y(_00095_));
 sky130_fd_sc_hd__nor2_1 _19612_ (.A(_12137_),
    .B(_12140_),
    .Y(_12205_));
 sky130_fd_sc_hd__nand2_1 _19613_ (.A(\cs_registers_i.mhpmcounter[2][22] ),
    .B(_12196_),
    .Y(_12206_));
 sky130_fd_sc_hd__nor3_1 _19614_ (.A(\cs_registers_i.mhpmcounter[2][23] ),
    .B(_12147_),
    .C(_12206_),
    .Y(_12207_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_649 ();
 sky130_fd_sc_hd__nor2_1 _19616_ (.A(_11664_),
    .B(_12139_),
    .Y(_12209_));
 sky130_fd_sc_hd__a21oi_1 _19617_ (.A1(_12139_),
    .A2(_12207_),
    .B1(_12209_),
    .Y(_12210_));
 sky130_fd_sc_hd__and2_4 _19618_ (.A(_11200_),
    .B(_12129_),
    .X(_12211_));
 sky130_fd_sc_hd__nand2_1 _19619_ (.A(_12211_),
    .B(_12148_),
    .Y(_12212_));
 sky130_fd_sc_hd__o211ai_1 _19620_ (.A1(_12212_),
    .A2(_12206_),
    .B1(\cs_registers_i.mhpmcounter[2][23] ),
    .C1(_12161_),
    .Y(_12213_));
 sky130_fd_sc_hd__o21ai_0 _19621_ (.A1(_12205_),
    .A2(_12210_),
    .B1(_12213_),
    .Y(_00096_));
 sky130_fd_sc_hd__and3_1 _19622_ (.A(\cs_registers_i.mhpmcounter[2][22] ),
    .B(\cs_registers_i.mhpmcounter[2][23] ),
    .C(_12196_),
    .X(_12214_));
 sky130_fd_sc_hd__nand2_1 _19623_ (.A(_12156_),
    .B(_12214_),
    .Y(_12215_));
 sky130_fd_sc_hd__nand3_1 _19624_ (.A(\cs_registers_i.mhpmcounter[2][24] ),
    .B(_12161_),
    .C(_12215_),
    .Y(_12216_));
 sky130_fd_sc_hd__o221ai_1 _19625_ (.A1(_11684_),
    .A2(_12161_),
    .B1(_12215_),
    .B2(\cs_registers_i.mhpmcounter[2][24] ),
    .C1(_12216_),
    .Y(_00097_));
 sky130_fd_sc_hd__and3_1 _19626_ (.A(\cs_registers_i.mhpmcounter[2][24] ),
    .B(_12156_),
    .C(_12214_),
    .X(_12217_));
 sky130_fd_sc_hd__nor3_1 _19627_ (.A(\cs_registers_i.mhpmcounter[2][25] ),
    .B(_12140_),
    .C(_12217_),
    .Y(_12218_));
 sky130_fd_sc_hd__a221oi_1 _19628_ (.A1(_11706_),
    .A2(_12140_),
    .B1(_12217_),
    .B2(\cs_registers_i.mhpmcounter[2][25] ),
    .C1(_12218_),
    .Y(_00098_));
 sky130_fd_sc_hd__nand4b_1 _19629_ (.A_N(\cs_registers_i.mhpmcounter[2][26] ),
    .B(_12214_),
    .C(\cs_registers_i.mhpmcounter[2][24] ),
    .D(\cs_registers_i.mhpmcounter[2][25] ),
    .Y(_12219_));
 sky130_fd_sc_hd__nand4_1 _19630_ (.A(\cs_registers_i.mhpmcounter[2][24] ),
    .B(\cs_registers_i.mhpmcounter[2][25] ),
    .C(_12156_),
    .D(_12214_),
    .Y(_12220_));
 sky130_fd_sc_hd__nand3_1 _19631_ (.A(\cs_registers_i.mhpmcounter[2][26] ),
    .B(_12134_),
    .C(_12220_),
    .Y(_12221_));
 sky130_fd_sc_hd__o221ai_1 _19632_ (.A1(_11726_),
    .A2(_12134_),
    .B1(_12212_),
    .B2(_12219_),
    .C1(_12221_),
    .Y(_00099_));
 sky130_fd_sc_hd__nand4_1 _19633_ (.A(\cs_registers_i.mhpmcounter[2][24] ),
    .B(\cs_registers_i.mhpmcounter[2][25] ),
    .C(\cs_registers_i.mhpmcounter[2][26] ),
    .D(_12214_),
    .Y(_12222_));
 sky130_fd_sc_hd__o32a_1 _19634_ (.A1(\cs_registers_i.mhpmcounter[2][27] ),
    .A2(_12155_),
    .A3(_12222_),
    .B1(_11746_),
    .B2(_12139_),
    .X(_12223_));
 sky130_fd_sc_hd__o211ai_1 _19635_ (.A1(_12212_),
    .A2(_12222_),
    .B1(\cs_registers_i.mhpmcounter[2][27] ),
    .C1(_12161_),
    .Y(_12224_));
 sky130_fd_sc_hd__o21ai_0 _19636_ (.A1(_12205_),
    .A2(_12223_),
    .B1(_12224_),
    .Y(_00100_));
 sky130_fd_sc_hd__and4_1 _19637_ (.A(\cs_registers_i.mhpmcounter[2][24] ),
    .B(\cs_registers_i.mhpmcounter[2][25] ),
    .C(\cs_registers_i.mhpmcounter[2][26] ),
    .D(_12214_),
    .X(_12225_));
 sky130_fd_sc_hd__nand2_1 _19638_ (.A(\cs_registers_i.mhpmcounter[2][27] ),
    .B(_12225_),
    .Y(_12226_));
 sky130_fd_sc_hd__nor3_1 _19639_ (.A(\cs_registers_i.mhpmcounter[2][28] ),
    .B(_12147_),
    .C(_12226_),
    .Y(_12227_));
 sky130_fd_sc_hd__nor2_1 _19640_ (.A(_11765_),
    .B(_12139_),
    .Y(_12228_));
 sky130_fd_sc_hd__a21oi_1 _19641_ (.A1(_12139_),
    .A2(_12227_),
    .B1(_12228_),
    .Y(_12229_));
 sky130_fd_sc_hd__o211ai_1 _19642_ (.A1(_12212_),
    .A2(_12226_),
    .B1(\cs_registers_i.mhpmcounter[2][28] ),
    .C1(_12161_),
    .Y(_12230_));
 sky130_fd_sc_hd__o21ai_0 _19643_ (.A1(_12205_),
    .A2(_12229_),
    .B1(_12230_),
    .Y(_00101_));
 sky130_fd_sc_hd__and3_1 _19644_ (.A(\cs_registers_i.mhpmcounter[2][27] ),
    .B(\cs_registers_i.mhpmcounter[2][28] ),
    .C(_12225_),
    .X(_12231_));
 sky130_fd_sc_hd__nand2_1 _19645_ (.A(_12156_),
    .B(_12231_),
    .Y(_12232_));
 sky130_fd_sc_hd__nand3_1 _19646_ (.A(\cs_registers_i.mhpmcounter[2][29] ),
    .B(_12161_),
    .C(_12232_),
    .Y(_12233_));
 sky130_fd_sc_hd__o221ai_1 _19647_ (.A1(_11785_),
    .A2(_12161_),
    .B1(_12232_),
    .B2(\cs_registers_i.mhpmcounter[2][29] ),
    .C1(_12233_),
    .Y(_00102_));
 sky130_fd_sc_hd__nand3_1 _19648_ (.A(\cs_registers_i.mhpmcounter[2][0] ),
    .B(\cs_registers_i.mhpmcounter[2][1] ),
    .C(_12137_),
    .Y(_12234_));
 sky130_fd_sc_hd__nand3_1 _19649_ (.A(\cs_registers_i.mhpmcounter[2][2] ),
    .B(_12161_),
    .C(_12234_),
    .Y(_12235_));
 sky130_fd_sc_hd__o21a_1 _19650_ (.A1(\cs_registers_i.mhpmcounter[2][2] ),
    .A2(_12234_),
    .B1(_12235_),
    .X(_12236_));
 sky130_fd_sc_hd__o21ai_0 _19651_ (.A1(_11309_),
    .A2(_12134_),
    .B1(_12236_),
    .Y(_00103_));
 sky130_fd_sc_hd__and3_1 _19652_ (.A(\cs_registers_i.mhpmcounter[2][29] ),
    .B(_12156_),
    .C(_12231_),
    .X(_12237_));
 sky130_fd_sc_hd__nor3_1 _19653_ (.A(\cs_registers_i.mhpmcounter[2][30] ),
    .B(_12140_),
    .C(_12237_),
    .Y(_12238_));
 sky130_fd_sc_hd__a221oi_1 _19654_ (.A1(_11808_),
    .A2(_12140_),
    .B1(_12237_),
    .B2(\cs_registers_i.mhpmcounter[2][30] ),
    .C1(_12238_),
    .Y(_00104_));
 sky130_fd_sc_hd__and3_1 _19655_ (.A(\cs_registers_i.mhpmcounter[2][29] ),
    .B(\cs_registers_i.mhpmcounter[2][30] ),
    .C(_12231_),
    .X(_12239_));
 sky130_fd_sc_hd__nand2_1 _19656_ (.A(\cs_registers_i.mhpmcounter[2][31] ),
    .B(_12239_),
    .Y(_12240_));
 sky130_fd_sc_hd__nor2_1 _19657_ (.A(_12147_),
    .B(_12240_),
    .Y(_12241_));
 sky130_fd_sc_hd__nor3_1 _19658_ (.A(\cs_registers_i.mhpmcounter[2][31] ),
    .B(_12140_),
    .C(_12156_),
    .Y(_12242_));
 sky130_fd_sc_hd__or3_1 _19659_ (.A(\cs_registers_i.mhpmcounter[2][31] ),
    .B(_12140_),
    .C(_12239_),
    .X(_12243_));
 sky130_fd_sc_hd__o21ai_0 _19660_ (.A1(_12106_),
    .A2(_12161_),
    .B1(_12243_),
    .Y(_12244_));
 sky130_fd_sc_hd__a211oi_1 _19661_ (.A1(_12137_),
    .A2(_12241_),
    .B1(_12242_),
    .C1(_12244_),
    .Y(_00105_));
 sky130_fd_sc_hd__nand2_4 _19662_ (.A(_12211_),
    .B(_12161_),
    .Y(_12245_));
 sky130_fd_sc_hd__nor2_2 _19663_ (.A(_11246_),
    .B(_11251_),
    .Y(_12246_));
 sky130_fd_sc_hd__nand3b_4 _19664_ (.A_N(_11225_),
    .B(_11243_),
    .C(_12246_),
    .Y(_12247_));
 sky130_fd_sc_hd__nand2_8 _19665_ (.A(_12245_),
    .B(_12247_),
    .Y(_12248_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_646 ();
 sky130_fd_sc_hd__nand2_1 _19669_ (.A(\cs_registers_i.mhpmcounter[2][32] ),
    .B(_12241_),
    .Y(_12252_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_645 ();
 sky130_fd_sc_hd__nand2_1 _19671_ (.A(_11280_),
    .B(_12131_),
    .Y(_12254_));
 sky130_fd_sc_hd__o21ai_0 _19672_ (.A1(_12131_),
    .A2(_12252_),
    .B1(_12254_),
    .Y(_12255_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_644 ();
 sky130_fd_sc_hd__o21ai_0 _19674_ (.A1(_12147_),
    .A2(_12240_),
    .B1(_12139_),
    .Y(_12257_));
 sky130_fd_sc_hd__a21oi_1 _19675_ (.A1(_12248_),
    .A2(_12257_),
    .B1(\cs_registers_i.mhpmcounter[2][32] ),
    .Y(_12258_));
 sky130_fd_sc_hd__a21oi_1 _19676_ (.A1(_12248_),
    .A2(_12255_),
    .B1(_12258_),
    .Y(_00106_));
 sky130_fd_sc_hd__and3_1 _19677_ (.A(\cs_registers_i.mhpmcounter[2][32] ),
    .B(\cs_registers_i.mhpmcounter[2][33] ),
    .C(_12241_),
    .X(_12259_));
 sky130_fd_sc_hd__nand2_1 _19678_ (.A(_12139_),
    .B(_12259_),
    .Y(_12260_));
 sky130_fd_sc_hd__nand2_1 _19679_ (.A(_11582_),
    .B(_12131_),
    .Y(_12261_));
 sky130_fd_sc_hd__nand2_1 _19680_ (.A(_12260_),
    .B(_12261_),
    .Y(_12262_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_643 ();
 sky130_fd_sc_hd__nand2_1 _19682_ (.A(_12139_),
    .B(_12252_),
    .Y(_12264_));
 sky130_fd_sc_hd__a21oi_1 _19683_ (.A1(_12248_),
    .A2(_12264_),
    .B1(\cs_registers_i.mhpmcounter[2][33] ),
    .Y(_12265_));
 sky130_fd_sc_hd__a21oi_1 _19684_ (.A1(_12248_),
    .A2(_12262_),
    .B1(_12265_),
    .Y(_00107_));
 sky130_fd_sc_hd__nand2_1 _19685_ (.A(_12211_),
    .B(_12259_),
    .Y(_12266_));
 sky130_fd_sc_hd__o21ai_0 _19686_ (.A1(_10928_),
    .A2(_12132_),
    .B1(_12266_),
    .Y(_12267_));
 sky130_fd_sc_hd__o21ai_0 _19687_ (.A1(_10926_),
    .A2(_12132_),
    .B1(_12267_),
    .Y(_12268_));
 sky130_fd_sc_hd__nand3b_1 _19688_ (.A_N(\cs_registers_i.mhpmcounter[2][34] ),
    .B(_12139_),
    .C(_12259_),
    .Y(_12269_));
 sky130_fd_sc_hd__o21ai_0 _19689_ (.A1(_11309_),
    .A2(_12139_),
    .B1(_12269_),
    .Y(_12270_));
 sky130_fd_sc_hd__a22o_1 _19690_ (.A1(\cs_registers_i.mhpmcounter[2][34] ),
    .A2(_12268_),
    .B1(_12270_),
    .B2(_12248_),
    .X(_00108_));
 sky130_fd_sc_hd__and4_1 _19691_ (.A(\cs_registers_i.mhpmcounter[2][32] ),
    .B(\cs_registers_i.mhpmcounter[2][33] ),
    .C(\cs_registers_i.mhpmcounter[2][34] ),
    .D(\cs_registers_i.mhpmcounter[2][35] ),
    .X(_12271_));
 sky130_fd_sc_hd__nand2_1 _19692_ (.A(_12241_),
    .B(_12271_),
    .Y(_12272_));
 sky130_fd_sc_hd__nand2_1 _19693_ (.A(_11867_),
    .B(_12131_),
    .Y(_12273_));
 sky130_fd_sc_hd__o21ai_0 _19694_ (.A1(_12131_),
    .A2(_12272_),
    .B1(_12273_),
    .Y(_12274_));
 sky130_fd_sc_hd__nand2_1 _19695_ (.A(\cs_registers_i.mhpmcounter[2][34] ),
    .B(_12259_),
    .Y(_12275_));
 sky130_fd_sc_hd__nand2_1 _19696_ (.A(_12139_),
    .B(_12275_),
    .Y(_12276_));
 sky130_fd_sc_hd__a21oi_1 _19697_ (.A1(_12248_),
    .A2(_12276_),
    .B1(\cs_registers_i.mhpmcounter[2][35] ),
    .Y(_12277_));
 sky130_fd_sc_hd__a21oi_1 _19698_ (.A1(_12248_),
    .A2(_12274_),
    .B1(_12277_),
    .Y(_00109_));
 sky130_fd_sc_hd__nand3_1 _19699_ (.A(\cs_registers_i.mhpmcounter[2][36] ),
    .B(_12241_),
    .C(_12271_),
    .Y(_12278_));
 sky130_fd_sc_hd__nand2_1 _19700_ (.A(_11887_),
    .B(_12131_),
    .Y(_12279_));
 sky130_fd_sc_hd__o21ai_0 _19701_ (.A1(_12131_),
    .A2(_12278_),
    .B1(_12279_),
    .Y(_12280_));
 sky130_fd_sc_hd__nand2_1 _19702_ (.A(_12139_),
    .B(_12272_),
    .Y(_12281_));
 sky130_fd_sc_hd__a21oi_1 _19703_ (.A1(_12248_),
    .A2(_12281_),
    .B1(\cs_registers_i.mhpmcounter[2][36] ),
    .Y(_12282_));
 sky130_fd_sc_hd__a21oi_1 _19704_ (.A1(_12248_),
    .A2(_12280_),
    .B1(_12282_),
    .Y(_00110_));
 sky130_fd_sc_hd__nand3_1 _19705_ (.A(\cs_registers_i.mhpmcounter[2][36] ),
    .B(\cs_registers_i.mhpmcounter[2][37] ),
    .C(_12271_),
    .Y(_12283_));
 sky130_fd_sc_hd__nor2_1 _19706_ (.A(_12240_),
    .B(_12283_),
    .Y(_12284_));
 sky130_fd_sc_hd__nand2_1 _19707_ (.A(_12148_),
    .B(_12284_),
    .Y(_12285_));
 sky130_fd_sc_hd__o21ai_0 _19708_ (.A1(_11902_),
    .A2(_12139_),
    .B1(_12285_),
    .Y(_12286_));
 sky130_fd_sc_hd__nand2_1 _19709_ (.A(_12139_),
    .B(_12278_),
    .Y(_12287_));
 sky130_fd_sc_hd__a21oi_1 _19710_ (.A1(_12248_),
    .A2(_12287_),
    .B1(\cs_registers_i.mhpmcounter[2][37] ),
    .Y(_12288_));
 sky130_fd_sc_hd__a21oi_1 _19711_ (.A1(_12248_),
    .A2(_12286_),
    .B1(_12288_),
    .Y(_00111_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_642 ();
 sky130_fd_sc_hd__nand2_1 _19713_ (.A(_12154_),
    .B(_12284_),
    .Y(_12290_));
 sky130_fd_sc_hd__nand2_1 _19714_ (.A(_12139_),
    .B(_12290_),
    .Y(_12291_));
 sky130_fd_sc_hd__a21oi_1 _19715_ (.A1(_12248_),
    .A2(_12291_),
    .B1(\cs_registers_i.mhpmcounter[2][38] ),
    .Y(_12292_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_641 ();
 sky130_fd_sc_hd__nand2_1 _19717_ (.A(\cs_registers_i.mhpmcounter[2][38] ),
    .B(_12284_),
    .Y(_12294_));
 sky130_fd_sc_hd__nor2_1 _19718_ (.A(_12155_),
    .B(_12294_),
    .Y(_12295_));
 sky130_fd_sc_hd__a21oi_1 _19719_ (.A1(_12113_),
    .A2(_12133_),
    .B1(_12295_),
    .Y(_12296_));
 sky130_fd_sc_hd__a21oi_1 _19720_ (.A1(_12245_),
    .A2(_12247_),
    .B1(_12296_),
    .Y(_12297_));
 sky130_fd_sc_hd__nor2_1 _19721_ (.A(_12292_),
    .B(_12297_),
    .Y(_00112_));
 sky130_fd_sc_hd__inv_1 _19722_ (.A(\cs_registers_i.mhpmcounter[2][39] ),
    .Y(_12298_));
 sky130_fd_sc_hd__nor3_2 _19723_ (.A(_12298_),
    .B(_12147_),
    .C(_12294_),
    .Y(_12299_));
 sky130_fd_sc_hd__nand2_1 _19724_ (.A(_12139_),
    .B(_12299_),
    .Y(_12300_));
 sky130_fd_sc_hd__nand2_1 _19725_ (.A(_11935_),
    .B(_12131_),
    .Y(_12301_));
 sky130_fd_sc_hd__nand2_1 _19726_ (.A(_12300_),
    .B(_12301_),
    .Y(_12302_));
 sky130_fd_sc_hd__o21ai_0 _19727_ (.A1(_12147_),
    .A2(_12294_),
    .B1(_12139_),
    .Y(_12303_));
 sky130_fd_sc_hd__a21oi_1 _19728_ (.A1(_12248_),
    .A2(_12303_),
    .B1(\cs_registers_i.mhpmcounter[2][39] ),
    .Y(_12304_));
 sky130_fd_sc_hd__a21oi_1 _19729_ (.A1(_12248_),
    .A2(_12302_),
    .B1(_12304_),
    .Y(_00113_));
 sky130_fd_sc_hd__a311oi_1 _19730_ (.A1(_12211_),
    .A2(_12139_),
    .A3(_12146_),
    .B1(_12140_),
    .C1(\cs_registers_i.mhpmcounter[2][3] ),
    .Y(_12305_));
 sky130_fd_sc_hd__a311oi_1 _19731_ (.A1(_10928_),
    .A2(_11867_),
    .A3(_12133_),
    .B1(_12156_),
    .C1(_12305_),
    .Y(_00114_));
 sky130_fd_sc_hd__inv_1 _19732_ (.A(\cs_registers_i.mhpmcounter[2][40] ),
    .Y(_12306_));
 sky130_fd_sc_hd__o21ai_0 _19733_ (.A1(_12133_),
    .A2(_12299_),
    .B1(_12248_),
    .Y(_12307_));
 sky130_fd_sc_hd__nand2_1 _19734_ (.A(\cs_registers_i.mhpmcounter[2][40] ),
    .B(_12299_),
    .Y(_12308_));
 sky130_fd_sc_hd__nand2_1 _19735_ (.A(_11957_),
    .B(_12131_),
    .Y(_12309_));
 sky130_fd_sc_hd__o21ai_0 _19736_ (.A1(_12131_),
    .A2(_12308_),
    .B1(_12309_),
    .Y(_12310_));
 sky130_fd_sc_hd__a22oi_1 _19737_ (.A1(_12306_),
    .A2(_12307_),
    .B1(_12310_),
    .B2(_12248_),
    .Y(_00115_));
 sky130_fd_sc_hd__nand4_2 _19738_ (.A(\cs_registers_i.mhpmcounter[2][39] ),
    .B(\cs_registers_i.mhpmcounter[2][40] ),
    .C(\cs_registers_i.mhpmcounter[2][41] ),
    .D(_12295_),
    .Y(_12311_));
 sky130_fd_sc_hd__nand2_1 _19739_ (.A(_11973_),
    .B(_12133_),
    .Y(_12312_));
 sky130_fd_sc_hd__nand2_1 _19740_ (.A(_12311_),
    .B(_12312_),
    .Y(_12313_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_640 ();
 sky130_fd_sc_hd__nand2_1 _19742_ (.A(_12139_),
    .B(_12308_),
    .Y(_12315_));
 sky130_fd_sc_hd__a21oi_1 _19743_ (.A1(_12248_),
    .A2(_12315_),
    .B1(\cs_registers_i.mhpmcounter[2][41] ),
    .Y(_12316_));
 sky130_fd_sc_hd__a21oi_1 _19744_ (.A1(_12248_),
    .A2(_12313_),
    .B1(_12316_),
    .Y(_00116_));
 sky130_fd_sc_hd__inv_1 _19745_ (.A(\cs_registers_i.mhpmcounter[2][42] ),
    .Y(_12317_));
 sky130_fd_sc_hd__o22ai_1 _19746_ (.A1(_11357_),
    .A2(_12139_),
    .B1(_12311_),
    .B2(_12317_),
    .Y(_12318_));
 sky130_fd_sc_hd__nand3_2 _19747_ (.A(\cs_registers_i.mhpmcounter[2][40] ),
    .B(\cs_registers_i.mhpmcounter[2][41] ),
    .C(_12299_),
    .Y(_12319_));
 sky130_fd_sc_hd__nand2_1 _19748_ (.A(_12139_),
    .B(_12319_),
    .Y(_12320_));
 sky130_fd_sc_hd__a21oi_1 _19749_ (.A1(_12248_),
    .A2(_12320_),
    .B1(\cs_registers_i.mhpmcounter[2][42] ),
    .Y(_12321_));
 sky130_fd_sc_hd__a21oi_1 _19750_ (.A1(_12248_),
    .A2(_12318_),
    .B1(_12321_),
    .Y(_00117_));
 sky130_fd_sc_hd__nand2_1 _19751_ (.A(\cs_registers_i.mhpmcounter[2][43] ),
    .B(\cs_registers_i.mhpmcounter[2][42] ),
    .Y(_12322_));
 sky130_fd_sc_hd__o22ai_1 _19752_ (.A1(_11391_),
    .A2(_12139_),
    .B1(_12311_),
    .B2(_12322_),
    .Y(_12323_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_639 ();
 sky130_fd_sc_hd__o21ai_0 _19754_ (.A1(_12317_),
    .A2(_12319_),
    .B1(_12139_),
    .Y(_12325_));
 sky130_fd_sc_hd__a21oi_1 _19755_ (.A1(_12248_),
    .A2(_12325_),
    .B1(\cs_registers_i.mhpmcounter[2][43] ),
    .Y(_12326_));
 sky130_fd_sc_hd__a21oi_1 _19756_ (.A1(_12248_),
    .A2(_12323_),
    .B1(_12326_),
    .Y(_00118_));
 sky130_fd_sc_hd__or2_0 _19757_ (.A(_12319_),
    .B(_12322_),
    .X(_12327_));
 sky130_fd_sc_hd__nor3_1 _19758_ (.A(\cs_registers_i.mhpmcounter[2][44] ),
    .B(_12131_),
    .C(_12327_),
    .Y(_12328_));
 sky130_fd_sc_hd__nor2_1 _19759_ (.A(_11428_),
    .B(_12139_),
    .Y(_12329_));
 sky130_fd_sc_hd__o21ai_0 _19760_ (.A1(_12328_),
    .A2(_12329_),
    .B1(_12248_),
    .Y(_12330_));
 sky130_fd_sc_hd__o211ai_1 _19761_ (.A1(_12245_),
    .A2(_12327_),
    .B1(_12247_),
    .C1(\cs_registers_i.mhpmcounter[2][44] ),
    .Y(_12331_));
 sky130_fd_sc_hd__nand2_1 _19762_ (.A(_12330_),
    .B(_12331_),
    .Y(_00119_));
 sky130_fd_sc_hd__nand4_1 _19763_ (.A(\cs_registers_i.mhpmcounter[2][44] ),
    .B(\cs_registers_i.mhpmcounter[2][43] ),
    .C(\cs_registers_i.mhpmcounter[2][42] ),
    .D(\cs_registers_i.mhpmcounter[2][45] ),
    .Y(_12332_));
 sky130_fd_sc_hd__nand2_1 _19764_ (.A(_11448_),
    .B(_12133_),
    .Y(_12333_));
 sky130_fd_sc_hd__o21ai_0 _19765_ (.A1(_12311_),
    .A2(_12332_),
    .B1(_12333_),
    .Y(_12334_));
 sky130_fd_sc_hd__inv_1 _19766_ (.A(\cs_registers_i.mhpmcounter[2][44] ),
    .Y(_12335_));
 sky130_fd_sc_hd__o21ai_0 _19767_ (.A1(_12335_),
    .A2(_12327_),
    .B1(_12139_),
    .Y(_12336_));
 sky130_fd_sc_hd__a21oi_1 _19768_ (.A1(_12248_),
    .A2(_12336_),
    .B1(\cs_registers_i.mhpmcounter[2][45] ),
    .Y(_12337_));
 sky130_fd_sc_hd__a21oi_1 _19769_ (.A1(_12248_),
    .A2(_12334_),
    .B1(_12337_),
    .Y(_00120_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_638 ();
 sky130_fd_sc_hd__nor2_1 _19771_ (.A(_12319_),
    .B(_12332_),
    .Y(_12339_));
 sky130_fd_sc_hd__nand2_1 _19772_ (.A(\cs_registers_i.mhpmcounter[2][46] ),
    .B(_12339_),
    .Y(_12340_));
 sky130_fd_sc_hd__nand2_1 _19773_ (.A(_11465_),
    .B(_12131_),
    .Y(_12341_));
 sky130_fd_sc_hd__o21ai_0 _19774_ (.A1(_12131_),
    .A2(_12340_),
    .B1(_12341_),
    .Y(_12342_));
 sky130_fd_sc_hd__o21ai_0 _19775_ (.A1(_12319_),
    .A2(_12332_),
    .B1(_12139_),
    .Y(_12343_));
 sky130_fd_sc_hd__a21oi_1 _19776_ (.A1(_12248_),
    .A2(_12343_),
    .B1(\cs_registers_i.mhpmcounter[2][46] ),
    .Y(_12344_));
 sky130_fd_sc_hd__a21oi_1 _19777_ (.A1(_12248_),
    .A2(_12342_),
    .B1(_12344_),
    .Y(_00121_));
 sky130_fd_sc_hd__nand3_1 _19778_ (.A(\cs_registers_i.mhpmcounter[2][46] ),
    .B(\cs_registers_i.mhpmcounter[2][47] ),
    .C(_12339_),
    .Y(_12345_));
 sky130_fd_sc_hd__nand2_1 _19779_ (.A(_11488_),
    .B(_12131_),
    .Y(_12346_));
 sky130_fd_sc_hd__o21ai_0 _19780_ (.A1(_12131_),
    .A2(_12345_),
    .B1(_12346_),
    .Y(_12347_));
 sky130_fd_sc_hd__nand2_1 _19781_ (.A(_12139_),
    .B(_12340_),
    .Y(_12348_));
 sky130_fd_sc_hd__a21oi_1 _19782_ (.A1(_12248_),
    .A2(_12348_),
    .B1(\cs_registers_i.mhpmcounter[2][47] ),
    .Y(_12349_));
 sky130_fd_sc_hd__a21oi_1 _19783_ (.A1(_12248_),
    .A2(_12347_),
    .B1(_12349_),
    .Y(_00122_));
 sky130_fd_sc_hd__inv_1 _19784_ (.A(_12332_),
    .Y(_12350_));
 sky130_fd_sc_hd__nand4_1 _19785_ (.A(\cs_registers_i.mhpmcounter[2][46] ),
    .B(\cs_registers_i.mhpmcounter[2][47] ),
    .C(\cs_registers_i.mhpmcounter[2][48] ),
    .D(_12350_),
    .Y(_12351_));
 sky130_fd_sc_hd__or2_1 _19786_ (.A(_12311_),
    .B(_12351_),
    .X(_12352_));
 sky130_fd_sc_hd__nand2_1 _19787_ (.A(_11505_),
    .B(_12133_),
    .Y(_12353_));
 sky130_fd_sc_hd__nand2_1 _19788_ (.A(_12352_),
    .B(_12353_),
    .Y(_12354_));
 sky130_fd_sc_hd__nand2_1 _19789_ (.A(_12139_),
    .B(_12345_),
    .Y(_12355_));
 sky130_fd_sc_hd__a21oi_1 _19790_ (.A1(_12248_),
    .A2(_12355_),
    .B1(\cs_registers_i.mhpmcounter[2][48] ),
    .Y(_12356_));
 sky130_fd_sc_hd__a21oi_1 _19791_ (.A1(_12248_),
    .A2(_12354_),
    .B1(_12356_),
    .Y(_00123_));
 sky130_fd_sc_hd__nor2_1 _19792_ (.A(_12319_),
    .B(_12351_),
    .Y(_12357_));
 sky130_fd_sc_hd__o21ai_0 _19793_ (.A1(_12133_),
    .A2(_12357_),
    .B1(_12248_),
    .Y(_12358_));
 sky130_fd_sc_hd__o22ai_1 _19794_ (.A1(_11523_),
    .A2(_12139_),
    .B1(_12352_),
    .B2(\cs_registers_i.mhpmcounter[2][49] ),
    .Y(_12359_));
 sky130_fd_sc_hd__a22o_1 _19795_ (.A1(\cs_registers_i.mhpmcounter[2][49] ),
    .A2(_12358_),
    .B1(_12359_),
    .B2(_12248_),
    .X(_00124_));
 sky130_fd_sc_hd__nor3_1 _19796_ (.A(\cs_registers_i.mhpmcounter[2][4] ),
    .B(_12140_),
    .C(_12156_),
    .Y(_12360_));
 sky130_fd_sc_hd__a221oi_1 _19797_ (.A1(_11887_),
    .A2(_12140_),
    .B1(_12156_),
    .B2(\cs_registers_i.mhpmcounter[2][4] ),
    .C1(_12360_),
    .Y(_00125_));
 sky130_fd_sc_hd__nand3_1 _19798_ (.A(\cs_registers_i.mhpmcounter[2][49] ),
    .B(\cs_registers_i.mhpmcounter[2][50] ),
    .C(_12357_),
    .Y(_12361_));
 sky130_fd_sc_hd__nand2_1 _19799_ (.A(_11546_),
    .B(net272),
    .Y(_12362_));
 sky130_fd_sc_hd__o21ai_0 _19800_ (.A1(net272),
    .A2(_12361_),
    .B1(_12362_),
    .Y(_12363_));
 sky130_fd_sc_hd__nand2_1 _19801_ (.A(\cs_registers_i.mhpmcounter[2][49] ),
    .B(_12357_),
    .Y(_12364_));
 sky130_fd_sc_hd__nand2_1 _19802_ (.A(_12139_),
    .B(_12364_),
    .Y(_12365_));
 sky130_fd_sc_hd__a21oi_1 _19803_ (.A1(_12248_),
    .A2(_12365_),
    .B1(\cs_registers_i.mhpmcounter[2][50] ),
    .Y(_12366_));
 sky130_fd_sc_hd__a21oi_1 _19804_ (.A1(_12248_),
    .A2(_12363_),
    .B1(_12366_),
    .Y(_00126_));
 sky130_fd_sc_hd__nand4_2 _19805_ (.A(\cs_registers_i.mhpmcounter[2][49] ),
    .B(\cs_registers_i.mhpmcounter[2][50] ),
    .C(\cs_registers_i.mhpmcounter[2][51] ),
    .D(_12357_),
    .Y(_12367_));
 sky130_fd_sc_hd__nand2_1 _19806_ (.A(_11563_),
    .B(_12133_),
    .Y(_12368_));
 sky130_fd_sc_hd__o21ai_0 _19807_ (.A1(net272),
    .A2(_12367_),
    .B1(_12368_),
    .Y(_12369_));
 sky130_fd_sc_hd__nand2_1 _19808_ (.A(_12139_),
    .B(_12361_),
    .Y(_12370_));
 sky130_fd_sc_hd__a21oi_1 _19809_ (.A1(_12248_),
    .A2(_12370_),
    .B1(\cs_registers_i.mhpmcounter[2][51] ),
    .Y(_12371_));
 sky130_fd_sc_hd__a21oi_1 _19810_ (.A1(_12248_),
    .A2(_12369_),
    .B1(_12371_),
    .Y(_00127_));
 sky130_fd_sc_hd__nor3_1 _19811_ (.A(\cs_registers_i.mhpmcounter[2][52] ),
    .B(_12133_),
    .C(_12367_),
    .Y(_12372_));
 sky130_fd_sc_hd__nor2_1 _19812_ (.A(_11599_),
    .B(_12139_),
    .Y(_12373_));
 sky130_fd_sc_hd__o21ai_0 _19813_ (.A1(_12372_),
    .A2(_12373_),
    .B1(_12248_),
    .Y(_12374_));
 sky130_fd_sc_hd__o211ai_1 _19814_ (.A1(_12245_),
    .A2(_12367_),
    .B1(_12247_),
    .C1(\cs_registers_i.mhpmcounter[2][52] ),
    .Y(_12375_));
 sky130_fd_sc_hd__nand2_1 _19815_ (.A(_12374_),
    .B(_12375_),
    .Y(_00128_));
 sky130_fd_sc_hd__nand2_1 _19816_ (.A(\cs_registers_i.mhpmcounter[2][49] ),
    .B(\cs_registers_i.mhpmcounter[2][50] ),
    .Y(_12376_));
 sky130_fd_sc_hd__nand3_1 _19817_ (.A(\cs_registers_i.mhpmcounter[2][51] ),
    .B(\cs_registers_i.mhpmcounter[2][52] ),
    .C(\cs_registers_i.mhpmcounter[2][53] ),
    .Y(_12377_));
 sky130_fd_sc_hd__o31ai_1 _19818_ (.A1(_12352_),
    .A2(_12376_),
    .A3(_12377_),
    .B1(_12199_),
    .Y(_12378_));
 sky130_fd_sc_hd__inv_1 _19819_ (.A(\cs_registers_i.mhpmcounter[2][52] ),
    .Y(_12379_));
 sky130_fd_sc_hd__o21ai_0 _19820_ (.A1(_12379_),
    .A2(_12367_),
    .B1(_12139_),
    .Y(_12380_));
 sky130_fd_sc_hd__a21oi_1 _19821_ (.A1(_12248_),
    .A2(_12380_),
    .B1(\cs_registers_i.mhpmcounter[2][53] ),
    .Y(_12381_));
 sky130_fd_sc_hd__a21oi_1 _19822_ (.A1(_12248_),
    .A2(_12378_),
    .B1(_12381_),
    .Y(_00129_));
 sky130_fd_sc_hd__nor2_1 _19823_ (.A(_12361_),
    .B(_12377_),
    .Y(_12382_));
 sky130_fd_sc_hd__and2_0 _19824_ (.A(\cs_registers_i.mhpmcounter[2][54] ),
    .B(_12382_),
    .X(_12383_));
 sky130_fd_sc_hd__nand2_1 _19825_ (.A(_12139_),
    .B(_12383_),
    .Y(_12384_));
 sky130_fd_sc_hd__nand2_1 _19826_ (.A(_11643_),
    .B(net272),
    .Y(_12385_));
 sky130_fd_sc_hd__nand2_1 _19827_ (.A(_12384_),
    .B(_12385_),
    .Y(_12386_));
 sky130_fd_sc_hd__o21ai_0 _19828_ (.A1(_12361_),
    .A2(_12377_),
    .B1(_12139_),
    .Y(_12387_));
 sky130_fd_sc_hd__a21oi_1 _19829_ (.A1(_12248_),
    .A2(_12387_),
    .B1(\cs_registers_i.mhpmcounter[2][54] ),
    .Y(_12388_));
 sky130_fd_sc_hd__a21oi_1 _19830_ (.A1(_12248_),
    .A2(_12386_),
    .B1(_12388_),
    .Y(_00130_));
 sky130_fd_sc_hd__inv_1 _19831_ (.A(\cs_registers_i.mhpmcounter[2][55] ),
    .Y(_12389_));
 sky130_fd_sc_hd__o21ai_0 _19832_ (.A1(_12133_),
    .A2(_12383_),
    .B1(_12248_),
    .Y(_12390_));
 sky130_fd_sc_hd__and3_1 _19833_ (.A(\cs_registers_i.mhpmcounter[2][54] ),
    .B(\cs_registers_i.mhpmcounter[2][55] ),
    .C(_12382_),
    .X(_12391_));
 sky130_fd_sc_hd__nand2_1 _19834_ (.A(_12139_),
    .B(_12391_),
    .Y(_12392_));
 sky130_fd_sc_hd__nand2_1 _19835_ (.A(_11664_),
    .B(net272),
    .Y(_12393_));
 sky130_fd_sc_hd__nand2_1 _19836_ (.A(_12392_),
    .B(_12393_),
    .Y(_12394_));
 sky130_fd_sc_hd__a22oi_1 _19837_ (.A1(_12389_),
    .A2(_12390_),
    .B1(_12394_),
    .B2(_12248_),
    .Y(_00131_));
 sky130_fd_sc_hd__nand3_1 _19838_ (.A(_12211_),
    .B(_12161_),
    .C(_12391_),
    .Y(_12395_));
 sky130_fd_sc_hd__nand3_1 _19839_ (.A(\cs_registers_i.mhpmcounter[2][56] ),
    .B(_12247_),
    .C(_12395_),
    .Y(_12396_));
 sky130_fd_sc_hd__o22ai_1 _19840_ (.A1(_11684_),
    .A2(_12139_),
    .B1(_12392_),
    .B2(\cs_registers_i.mhpmcounter[2][56] ),
    .Y(_12397_));
 sky130_fd_sc_hd__nand2_1 _19841_ (.A(_12248_),
    .B(_12397_),
    .Y(_12398_));
 sky130_fd_sc_hd__nand2_1 _19842_ (.A(_12396_),
    .B(_12398_),
    .Y(_00132_));
 sky130_fd_sc_hd__nand2_1 _19843_ (.A(\cs_registers_i.mhpmcounter[2][56] ),
    .B(\cs_registers_i.mhpmcounter[2][57] ),
    .Y(_12399_));
 sky130_fd_sc_hd__nand2_1 _19844_ (.A(_11706_),
    .B(net272),
    .Y(_12400_));
 sky130_fd_sc_hd__o21ai_0 _19845_ (.A1(_12392_),
    .A2(_12399_),
    .B1(_12400_),
    .Y(_12401_));
 sky130_fd_sc_hd__nand2_1 _19846_ (.A(\cs_registers_i.mhpmcounter[2][56] ),
    .B(_12391_),
    .Y(_12402_));
 sky130_fd_sc_hd__nand2_1 _19847_ (.A(_12139_),
    .B(_12402_),
    .Y(_12403_));
 sky130_fd_sc_hd__a21oi_1 _19848_ (.A1(_12248_),
    .A2(_12403_),
    .B1(\cs_registers_i.mhpmcounter[2][57] ),
    .Y(_12404_));
 sky130_fd_sc_hd__a21oi_1 _19849_ (.A1(_12248_),
    .A2(_12401_),
    .B1(_12404_),
    .Y(_00133_));
 sky130_fd_sc_hd__inv_1 _19850_ (.A(\cs_registers_i.mhpmcounter[2][58] ),
    .Y(_12405_));
 sky130_fd_sc_hd__and3_1 _19851_ (.A(\cs_registers_i.mhpmcounter[2][56] ),
    .B(\cs_registers_i.mhpmcounter[2][57] ),
    .C(_12391_),
    .X(_12406_));
 sky130_fd_sc_hd__o21ai_0 _19852_ (.A1(_12133_),
    .A2(_12406_),
    .B1(_12248_),
    .Y(_12407_));
 sky130_fd_sc_hd__nand2_1 _19853_ (.A(\cs_registers_i.mhpmcounter[2][58] ),
    .B(_12406_),
    .Y(_12408_));
 sky130_fd_sc_hd__nand2_1 _19854_ (.A(_11726_),
    .B(net272),
    .Y(_12409_));
 sky130_fd_sc_hd__o21ai_0 _19855_ (.A1(net272),
    .A2(_12408_),
    .B1(_12409_),
    .Y(_12410_));
 sky130_fd_sc_hd__a22oi_1 _19856_ (.A1(_12405_),
    .A2(_12407_),
    .B1(_12410_),
    .B2(_12248_),
    .Y(_00134_));
 sky130_fd_sc_hd__and3_1 _19857_ (.A(\cs_registers_i.mhpmcounter[2][58] ),
    .B(\cs_registers_i.mhpmcounter[2][59] ),
    .C(_12406_),
    .X(_12411_));
 sky130_fd_sc_hd__nand2_1 _19858_ (.A(_12139_),
    .B(_12411_),
    .Y(_12412_));
 sky130_fd_sc_hd__nand2_1 _19859_ (.A(_11746_),
    .B(net272),
    .Y(_12413_));
 sky130_fd_sc_hd__nand2_1 _19860_ (.A(_12412_),
    .B(_12413_),
    .Y(_12414_));
 sky130_fd_sc_hd__nand2_1 _19861_ (.A(_12139_),
    .B(_12408_),
    .Y(_12415_));
 sky130_fd_sc_hd__a21oi_1 _19862_ (.A1(_12248_),
    .A2(_12415_),
    .B1(\cs_registers_i.mhpmcounter[2][59] ),
    .Y(_12416_));
 sky130_fd_sc_hd__a21oi_1 _19863_ (.A1(_12248_),
    .A2(_12414_),
    .B1(_12416_),
    .Y(_00135_));
 sky130_fd_sc_hd__nand3_1 _19864_ (.A(\cs_registers_i.mhpmcounter[2][4] ),
    .B(\cs_registers_i.mhpmcounter[2][5] ),
    .C(_12148_),
    .Y(_12417_));
 sky130_fd_sc_hd__o21ai_0 _19865_ (.A1(_11902_),
    .A2(_12139_),
    .B1(_12417_),
    .Y(_12418_));
 sky130_fd_sc_hd__a211oi_1 _19866_ (.A1(\cs_registers_i.mhpmcounter[2][4] ),
    .A2(_12156_),
    .B1(_12140_),
    .C1(\cs_registers_i.mhpmcounter[2][5] ),
    .Y(_12419_));
 sky130_fd_sc_hd__a21oi_1 _19867_ (.A1(_12136_),
    .A2(_12418_),
    .B1(_12419_),
    .Y(_00136_));
 sky130_fd_sc_hd__inv_1 _19868_ (.A(\cs_registers_i.mhpmcounter[2][60] ),
    .Y(_12420_));
 sky130_fd_sc_hd__o21ai_0 _19869_ (.A1(_12133_),
    .A2(_12411_),
    .B1(_12248_),
    .Y(_12421_));
 sky130_fd_sc_hd__nand2_1 _19870_ (.A(\cs_registers_i.mhpmcounter[2][60] ),
    .B(_12411_),
    .Y(_12422_));
 sky130_fd_sc_hd__nor2_1 _19871_ (.A(_12131_),
    .B(_12422_),
    .Y(_12423_));
 sky130_fd_sc_hd__a21o_1 _19872_ (.A1(_11765_),
    .A2(_12131_),
    .B1(_12423_),
    .X(_12424_));
 sky130_fd_sc_hd__a22oi_1 _19873_ (.A1(_12420_),
    .A2(_12421_),
    .B1(_12424_),
    .B2(_12248_),
    .Y(_00137_));
 sky130_fd_sc_hd__a22o_1 _19874_ (.A1(_11785_),
    .A2(_12131_),
    .B1(_12423_),
    .B2(\cs_registers_i.mhpmcounter[2][61] ),
    .X(_12425_));
 sky130_fd_sc_hd__nand2_1 _19875_ (.A(_12139_),
    .B(_12422_),
    .Y(_12426_));
 sky130_fd_sc_hd__a21oi_1 _19876_ (.A1(_12248_),
    .A2(_12426_),
    .B1(\cs_registers_i.mhpmcounter[2][61] ),
    .Y(_12427_));
 sky130_fd_sc_hd__a21oi_1 _19877_ (.A1(_12248_),
    .A2(_12425_),
    .B1(_12427_),
    .Y(_00138_));
 sky130_fd_sc_hd__inv_1 _19878_ (.A(\cs_registers_i.mhpmcounter[2][62] ),
    .Y(_12428_));
 sky130_fd_sc_hd__and3_1 _19879_ (.A(\cs_registers_i.mhpmcounter[2][60] ),
    .B(\cs_registers_i.mhpmcounter[2][61] ),
    .C(_12411_),
    .X(_12429_));
 sky130_fd_sc_hd__o21ai_0 _19880_ (.A1(_12133_),
    .A2(_12429_),
    .B1(_12248_),
    .Y(_12430_));
 sky130_fd_sc_hd__nand2_1 _19881_ (.A(\cs_registers_i.mhpmcounter[2][62] ),
    .B(_12429_),
    .Y(_12431_));
 sky130_fd_sc_hd__nand2_1 _19882_ (.A(_11808_),
    .B(_12131_),
    .Y(_12432_));
 sky130_fd_sc_hd__o21ai_0 _19883_ (.A1(_12131_),
    .A2(_12431_),
    .B1(_12432_),
    .Y(_12433_));
 sky130_fd_sc_hd__a22oi_1 _19884_ (.A1(_12428_),
    .A2(_12430_),
    .B1(_12433_),
    .B2(_12248_),
    .Y(_00139_));
 sky130_fd_sc_hd__nand4_1 _19885_ (.A(\cs_registers_i.mhpmcounter[2][62] ),
    .B(\cs_registers_i.mhpmcounter[2][63] ),
    .C(_12139_),
    .D(_12429_),
    .Y(_12434_));
 sky130_fd_sc_hd__o21ai_0 _19886_ (.A1(_12106_),
    .A2(_12139_),
    .B1(_12434_),
    .Y(_12435_));
 sky130_fd_sc_hd__nand2_1 _19887_ (.A(_12139_),
    .B(_12431_),
    .Y(_12436_));
 sky130_fd_sc_hd__a21oi_1 _19888_ (.A1(_12248_),
    .A2(_12436_),
    .B1(\cs_registers_i.mhpmcounter[2][63] ),
    .Y(_12437_));
 sky130_fd_sc_hd__a21oi_1 _19889_ (.A1(_12248_),
    .A2(_12435_),
    .B1(_12437_),
    .Y(_00140_));
 sky130_fd_sc_hd__nor2_1 _19890_ (.A(\cs_registers_i.mhpmcounter[2][6] ),
    .B(_12140_),
    .Y(_12438_));
 sky130_fd_sc_hd__o21a_1 _19891_ (.A1(_12130_),
    .A2(_12417_),
    .B1(_12438_),
    .X(_12439_));
 sky130_fd_sc_hd__a221oi_1 _19892_ (.A1(_12113_),
    .A2(_12140_),
    .B1(_12149_),
    .B2(_12156_),
    .C1(_12439_),
    .Y(_00141_));
 sky130_fd_sc_hd__a211oi_1 _19893_ (.A1(_12149_),
    .A2(_12156_),
    .B1(\cs_registers_i.mhpmcounter[2][7] ),
    .C1(_12140_),
    .Y(_12440_));
 sky130_fd_sc_hd__and3_1 _19894_ (.A(\cs_registers_i.mhpmcounter[2][7] ),
    .B(_12149_),
    .C(_12156_),
    .X(_12441_));
 sky130_fd_sc_hd__a211oi_1 _19895_ (.A1(_11935_),
    .A2(_12140_),
    .B1(_12440_),
    .C1(_12441_),
    .Y(_00142_));
 sky130_fd_sc_hd__nor3_1 _19896_ (.A(\cs_registers_i.mhpmcounter[2][8] ),
    .B(_12140_),
    .C(_12441_),
    .Y(_12442_));
 sky130_fd_sc_hd__and2_0 _19897_ (.A(\cs_registers_i.mhpmcounter[2][8] ),
    .B(_12441_),
    .X(_12443_));
 sky130_fd_sc_hd__a211oi_1 _19898_ (.A1(_11957_),
    .A2(_12140_),
    .B1(_12442_),
    .C1(_12443_),
    .Y(_00143_));
 sky130_fd_sc_hd__nor3_1 _19899_ (.A(\cs_registers_i.mhpmcounter[2][9] ),
    .B(_12140_),
    .C(_12443_),
    .Y(_12444_));
 sky130_fd_sc_hd__o21ai_0 _19900_ (.A1(_10914_),
    .A2(_10927_),
    .B1(_11267_),
    .Y(_12445_));
 sky130_fd_sc_hd__nor2_1 _19901_ (.A(_11313_),
    .B(_12445_),
    .Y(_12446_));
 sky130_fd_sc_hd__nand2_1 _19902_ (.A(_12150_),
    .B(_12154_),
    .Y(_12447_));
 sky130_fd_sc_hd__a211oi_1 _19903_ (.A1(_10925_),
    .A2(_12446_),
    .B1(_12447_),
    .C1(_12130_),
    .Y(_12448_));
 sky130_fd_sc_hd__a211oi_1 _19904_ (.A1(_11973_),
    .A2(_12140_),
    .B1(_12444_),
    .C1(_12448_),
    .Y(_00144_));
 sky130_fd_sc_hd__and2_1 _19905_ (.A(_08143_),
    .B(_11000_),
    .X(_12449_));
 sky130_fd_sc_hd__nand3_4 _19906_ (.A(_08111_),
    .B(_08117_),
    .C(_12449_),
    .Y(_12450_));
 sky130_fd_sc_hd__nand2_8 _19907_ (.A(_10946_),
    .B(_10995_),
    .Y(_12451_));
 sky130_fd_sc_hd__nor2_8 _19908_ (.A(_12450_),
    .B(_12451_),
    .Y(_12452_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_636 ();
 sky130_fd_sc_hd__nor2_8 _19911_ (.A(_10935_),
    .B(_12451_),
    .Y(_12455_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_635 ();
 sky130_fd_sc_hd__nor2b_1 _19913_ (.A(_12455_),
    .B_N(\cs_registers_i.priv_lvl_q[0] ),
    .Y(_12457_));
 sky130_fd_sc_hd__nand2_2 _19914_ (.A(_10940_),
    .B(_12449_),
    .Y(_12458_));
 sky130_fd_sc_hd__nor2_8 _19915_ (.A(_12458_),
    .B(_12451_),
    .Y(_12459_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_633 ();
 sky130_fd_sc_hd__a211oi_1 _19918_ (.A1(\cs_registers_i.mstack_d[0] ),
    .A2(_12452_),
    .B1(_12457_),
    .C1(_12459_),
    .Y(_12462_));
 sky130_fd_sc_hd__nor3_1 _19919_ (.A(\cs_registers_i.dcsr_q[0] ),
    .B(_10941_),
    .C(_12451_),
    .Y(_12463_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_631 ();
 sky130_fd_sc_hd__a22oi_4 _19922_ (.A1(\cs_registers_i.dcsr_q[15] ),
    .A2(_10937_),
    .B1(_10997_),
    .B2(\cs_registers_i.dcsr_q[12] ),
    .Y(_12466_));
 sky130_fd_sc_hd__o22a_2 _19923_ (.A1(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .A2(_11007_),
    .B1(_11031_),
    .B2(_12466_),
    .X(_12467_));
 sky130_fd_sc_hd__nor2_8 _19924_ (.A(_11009_),
    .B(_12467_),
    .Y(_12468_));
 sky130_fd_sc_hd__nor3_4 _19925_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .B(_10945_),
    .C(_10995_),
    .Y(_12469_));
 sky130_fd_sc_hd__o21a_1 _19926_ (.A1(_10999_),
    .A2(_11002_),
    .B1(_12469_),
    .X(_12470_));
 sky130_fd_sc_hd__nor3_2 _19927_ (.A(_11034_),
    .B(_12468_),
    .C(_12470_),
    .Y(_12471_));
 sky130_fd_sc_hd__o21ai_0 _19928_ (.A1(_12462_),
    .A2(_12463_),
    .B1(_12471_),
    .Y(_00145_));
 sky130_fd_sc_hd__nor2_1 _19929_ (.A(_10859_),
    .B(_12455_),
    .Y(_12472_));
 sky130_fd_sc_hd__a211oi_1 _19930_ (.A1(\cs_registers_i.mstack_d[1] ),
    .A2(_12452_),
    .B1(_12459_),
    .C1(_12472_),
    .Y(_12473_));
 sky130_fd_sc_hd__nor3_1 _19931_ (.A(\cs_registers_i.dcsr_q[1] ),
    .B(_10941_),
    .C(_12451_),
    .Y(_12474_));
 sky130_fd_sc_hd__o21ai_0 _19932_ (.A1(_12473_),
    .A2(_12474_),
    .B1(_12471_),
    .Y(_00146_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_630 ();
 sky130_fd_sc_hd__a21oi_1 _19934_ (.A1(_11243_),
    .A2(_11248_),
    .B1(\cs_registers_i.dcsr_q[0] ),
    .Y(_12476_));
 sky130_fd_sc_hd__nand2_4 _19935_ (.A(_11243_),
    .B(_11248_),
    .Y(_12477_));
 sky130_fd_sc_hd__nand2_1 _19936_ (.A(_11280_),
    .B(_11582_),
    .Y(_12478_));
 sky130_fd_sc_hd__nor2_1 _19937_ (.A(_12477_),
    .B(_12478_),
    .Y(_12479_));
 sky130_fd_sc_hd__nand2_1 _19938_ (.A(\cs_registers_i.priv_lvl_q[0] ),
    .B(_12468_),
    .Y(_12480_));
 sky130_fd_sc_hd__o31ai_1 _19939_ (.A1(_12468_),
    .A2(_12476_),
    .A3(_12479_),
    .B1(_12480_),
    .Y(_00147_));
 sky130_fd_sc_hd__a31oi_4 _19940_ (.A1(net878),
    .A2(_11146_),
    .A3(_11389_),
    .B1(_11390_),
    .Y(_12481_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_629 ();
 sky130_fd_sc_hd__nand2_1 _19942_ (.A(\cs_registers_i.dcsr_q[11] ),
    .B(_12477_),
    .Y(_12483_));
 sky130_fd_sc_hd__o21ai_0 _19943_ (.A1(_12481_),
    .A2(_12477_),
    .B1(_12483_),
    .Y(_00148_));
 sky130_fd_sc_hd__nand2_1 _19944_ (.A(\cs_registers_i.dcsr_q[12] ),
    .B(_12477_),
    .Y(_12484_));
 sky130_fd_sc_hd__o21ai_0 _19945_ (.A1(_11428_),
    .A2(_12477_),
    .B1(_12484_),
    .Y(_00149_));
 sky130_fd_sc_hd__nand2_1 _19946_ (.A(\cs_registers_i.dcsr_q[13] ),
    .B(_12477_),
    .Y(_12485_));
 sky130_fd_sc_hd__o21ai_0 _19947_ (.A1(_11448_),
    .A2(_12477_),
    .B1(_12485_),
    .Y(_00150_));
 sky130_fd_sc_hd__nand2_1 _19948_ (.A(\cs_registers_i.dcsr_q[15] ),
    .B(_12477_),
    .Y(_12486_));
 sky130_fd_sc_hd__o21ai_0 _19949_ (.A1(_11488_),
    .A2(_12477_),
    .B1(_12486_),
    .Y(_00151_));
 sky130_fd_sc_hd__a21oi_1 _19950_ (.A1(_11243_),
    .A2(_11248_),
    .B1(\cs_registers_i.dcsr_q[1] ),
    .Y(_12487_));
 sky130_fd_sc_hd__nand2_1 _19951_ (.A(\cs_registers_i.priv_lvl_q[1] ),
    .B(_12468_),
    .Y(_12488_));
 sky130_fd_sc_hd__o31ai_1 _19952_ (.A1(_12468_),
    .A2(_12479_),
    .A3(_12487_),
    .B1(_12488_),
    .Y(_00152_));
 sky130_fd_sc_hd__nand2_1 _19953_ (.A(\cs_registers_i.dcsr_q[2] ),
    .B(_12477_),
    .Y(_12489_));
 sky130_fd_sc_hd__o21ai_0 _19954_ (.A1(_11309_),
    .A2(_12477_),
    .B1(_12489_),
    .Y(_00153_));
 sky130_fd_sc_hd__nor2_1 _19955_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .B(_11009_),
    .Y(_12490_));
 sky130_fd_sc_hd__nand2_1 _19956_ (.A(\cs_registers_i.dcsr_q[2] ),
    .B(_12490_),
    .Y(_12491_));
 sky130_fd_sc_hd__o21a_1 _19957_ (.A1(\cs_registers_i.dcsr_q[6] ),
    .A2(_12468_),
    .B1(_12491_),
    .X(_00154_));
 sky130_fd_sc_hd__o21ai_0 _19958_ (.A1(_11009_),
    .A2(_12467_),
    .B1(\cs_registers_i.dcsr_q[7] ),
    .Y(_12492_));
 sky130_fd_sc_hd__nand3b_1 _19959_ (.A_N(\cs_registers_i.dcsr_q[2] ),
    .B(net60),
    .C(_12490_),
    .Y(_12493_));
 sky130_fd_sc_hd__nand2_1 _19960_ (.A(_12492_),
    .B(_12493_),
    .Y(_00155_));
 sky130_fd_sc_hd__o21ai_0 _19961_ (.A1(_11009_),
    .A2(_12467_),
    .B1(\cs_registers_i.dcsr_q[8] ),
    .Y(_12494_));
 sky130_fd_sc_hd__nand2_1 _19962_ (.A(_12491_),
    .B(_12494_),
    .Y(_00156_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_627 ();
 sky130_fd_sc_hd__nor3_2 _19965_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .B(_11009_),
    .C(_11007_),
    .Y(_12497_));
 sky130_fd_sc_hd__nor2_8 _19966_ (.A(_11034_),
    .B(_12497_),
    .Y(_12498_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_626 ();
 sky130_fd_sc_hd__mux2i_1 _19968_ (.A0(\cs_registers_i.pc_if_i[10] ),
    .A1(\cs_registers_i.pc_id_i[10] ),
    .S(_12498_),
    .Y(_12500_));
 sky130_fd_sc_hd__nand2_8 _19969_ (.A(_11243_),
    .B(_11295_),
    .Y(_12501_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_625 ();
 sky130_fd_sc_hd__and3_1 _19971_ (.A(_11243_),
    .B(_11295_),
    .C(_11357_),
    .X(_12503_));
 sky130_fd_sc_hd__a211oi_1 _19972_ (.A1(\cs_registers_i.csr_depc_o[10] ),
    .A2(_12501_),
    .B1(_12503_),
    .C1(_12468_),
    .Y(_12504_));
 sky130_fd_sc_hd__a21oi_1 _19973_ (.A1(_12468_),
    .A2(_12500_),
    .B1(_12504_),
    .Y(_00157_));
 sky130_fd_sc_hd__mux2i_1 _19974_ (.A0(\cs_registers_i.pc_if_i[11] ),
    .A1(\cs_registers_i.pc_id_i[11] ),
    .S(_12498_),
    .Y(_12505_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_624 ();
 sky130_fd_sc_hd__nor2_1 _19976_ (.A(_12481_),
    .B(_12501_),
    .Y(_12507_));
 sky130_fd_sc_hd__a211oi_1 _19977_ (.A1(\cs_registers_i.csr_depc_o[11] ),
    .A2(_12501_),
    .B1(_12507_),
    .C1(_12468_),
    .Y(_12508_));
 sky130_fd_sc_hd__a21oi_1 _19978_ (.A1(_12468_),
    .A2(_12505_),
    .B1(_12508_),
    .Y(_00158_));
 sky130_fd_sc_hd__mux2i_1 _19979_ (.A0(\cs_registers_i.pc_if_i[12] ),
    .A1(\cs_registers_i.pc_id_i[12] ),
    .S(_12498_),
    .Y(_12509_));
 sky130_fd_sc_hd__nor2_1 _19980_ (.A(_11428_),
    .B(_12501_),
    .Y(_12510_));
 sky130_fd_sc_hd__a211oi_1 _19981_ (.A1(\cs_registers_i.csr_depc_o[12] ),
    .A2(_12501_),
    .B1(_12510_),
    .C1(_12468_),
    .Y(_12511_));
 sky130_fd_sc_hd__a21oi_1 _19982_ (.A1(_12468_),
    .A2(_12509_),
    .B1(_12511_),
    .Y(_00159_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_623 ();
 sky130_fd_sc_hd__mux2i_1 _19984_ (.A0(\cs_registers_i.pc_if_i[13] ),
    .A1(\cs_registers_i.pc_id_i[13] ),
    .S(_12498_),
    .Y(_12513_));
 sky130_fd_sc_hd__nor2_1 _19985_ (.A(_11448_),
    .B(_12501_),
    .Y(_12514_));
 sky130_fd_sc_hd__a211oi_1 _19986_ (.A1(\cs_registers_i.csr_depc_o[13] ),
    .A2(_12501_),
    .B1(_12514_),
    .C1(_12468_),
    .Y(_12515_));
 sky130_fd_sc_hd__a21oi_1 _19987_ (.A1(_12468_),
    .A2(_12513_),
    .B1(_12515_),
    .Y(_00160_));
 sky130_fd_sc_hd__mux2i_1 _19988_ (.A0(\cs_registers_i.pc_if_i[14] ),
    .A1(\cs_registers_i.pc_id_i[14] ),
    .S(_12498_),
    .Y(_12516_));
 sky130_fd_sc_hd__nor2_1 _19989_ (.A(_11465_),
    .B(_12501_),
    .Y(_12517_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_622 ();
 sky130_fd_sc_hd__a211oi_1 _19991_ (.A1(\cs_registers_i.csr_depc_o[14] ),
    .A2(_12501_),
    .B1(_12517_),
    .C1(_12468_),
    .Y(_12519_));
 sky130_fd_sc_hd__a21oi_1 _19992_ (.A1(_12468_),
    .A2(_12516_),
    .B1(_12519_),
    .Y(_00161_));
 sky130_fd_sc_hd__mux2i_1 _19993_ (.A0(\cs_registers_i.pc_if_i[15] ),
    .A1(\cs_registers_i.pc_id_i[15] ),
    .S(_12498_),
    .Y(_12520_));
 sky130_fd_sc_hd__nor2_1 _19994_ (.A(_11488_),
    .B(_12501_),
    .Y(_12521_));
 sky130_fd_sc_hd__a211oi_1 _19995_ (.A1(\cs_registers_i.csr_depc_o[15] ),
    .A2(_12501_),
    .B1(_12521_),
    .C1(_12468_),
    .Y(_12522_));
 sky130_fd_sc_hd__a21oi_1 _19996_ (.A1(_12468_),
    .A2(_12520_),
    .B1(_12522_),
    .Y(_00162_));
 sky130_fd_sc_hd__mux2i_2 _19997_ (.A0(\cs_registers_i.pc_if_i[16] ),
    .A1(\cs_registers_i.pc_id_i[16] ),
    .S(_12498_),
    .Y(_12523_));
 sky130_fd_sc_hd__nor2_1 _19998_ (.A(_11505_),
    .B(_12501_),
    .Y(_12524_));
 sky130_fd_sc_hd__a211oi_1 _19999_ (.A1(\cs_registers_i.csr_depc_o[16] ),
    .A2(_12501_),
    .B1(_12524_),
    .C1(_12468_),
    .Y(_12525_));
 sky130_fd_sc_hd__a21oi_1 _20000_ (.A1(_12468_),
    .A2(_12523_),
    .B1(_12525_),
    .Y(_00163_));
 sky130_fd_sc_hd__mux2i_2 _20001_ (.A0(\cs_registers_i.pc_if_i[17] ),
    .A1(\cs_registers_i.pc_id_i[17] ),
    .S(_12498_),
    .Y(_12526_));
 sky130_fd_sc_hd__nor2_1 _20002_ (.A(_11523_),
    .B(_12501_),
    .Y(_12527_));
 sky130_fd_sc_hd__a211oi_1 _20003_ (.A1(\cs_registers_i.csr_depc_o[17] ),
    .A2(_12501_),
    .B1(_12527_),
    .C1(_12468_),
    .Y(_12528_));
 sky130_fd_sc_hd__a21oi_1 _20004_ (.A1(_12468_),
    .A2(_12526_),
    .B1(_12528_),
    .Y(_00164_));
 sky130_fd_sc_hd__mux2i_1 _20005_ (.A0(\cs_registers_i.pc_if_i[18] ),
    .A1(\cs_registers_i.pc_id_i[18] ),
    .S(_12498_),
    .Y(_12529_));
 sky130_fd_sc_hd__nor2_1 _20006_ (.A(_11546_),
    .B(_12501_),
    .Y(_12530_));
 sky130_fd_sc_hd__a211oi_1 _20007_ (.A1(\cs_registers_i.csr_depc_o[18] ),
    .A2(_12501_),
    .B1(_12530_),
    .C1(_12468_),
    .Y(_12531_));
 sky130_fd_sc_hd__a21oi_1 _20008_ (.A1(_12468_),
    .A2(_12529_),
    .B1(_12531_),
    .Y(_00165_));
 sky130_fd_sc_hd__mux2i_2 _20009_ (.A0(\cs_registers_i.pc_if_i[19] ),
    .A1(\cs_registers_i.pc_id_i[19] ),
    .S(_12498_),
    .Y(_12532_));
 sky130_fd_sc_hd__nor2_1 _20010_ (.A(_11563_),
    .B(_12501_),
    .Y(_12533_));
 sky130_fd_sc_hd__a211oi_1 _20011_ (.A1(\cs_registers_i.csr_depc_o[19] ),
    .A2(_12501_),
    .B1(_12533_),
    .C1(_12468_),
    .Y(_12534_));
 sky130_fd_sc_hd__a21oi_1 _20012_ (.A1(_12468_),
    .A2(_12532_),
    .B1(_12534_),
    .Y(_00166_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_619 ();
 sky130_fd_sc_hd__mux2i_1 _20016_ (.A0(\cs_registers_i.pc_if_i[1] ),
    .A1(\cs_registers_i.pc_id_i[1] ),
    .S(_12498_),
    .Y(_12538_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_617 ();
 sky130_fd_sc_hd__nor2_1 _20019_ (.A(_11582_),
    .B(_12501_),
    .Y(_12541_));
 sky130_fd_sc_hd__a211oi_1 _20020_ (.A1(\cs_registers_i.csr_depc_o[1] ),
    .A2(_12501_),
    .B1(_12541_),
    .C1(_12468_),
    .Y(_12542_));
 sky130_fd_sc_hd__a21oi_1 _20021_ (.A1(_12468_),
    .A2(_12538_),
    .B1(_12542_),
    .Y(_00167_));
 sky130_fd_sc_hd__mux2i_1 _20022_ (.A0(\cs_registers_i.pc_if_i[20] ),
    .A1(\cs_registers_i.pc_id_i[20] ),
    .S(_12498_),
    .Y(_12543_));
 sky130_fd_sc_hd__nor2_1 _20023_ (.A(_11599_),
    .B(_12501_),
    .Y(_12544_));
 sky130_fd_sc_hd__a211oi_1 _20024_ (.A1(\cs_registers_i.csr_depc_o[20] ),
    .A2(_12501_),
    .B1(_12544_),
    .C1(_12468_),
    .Y(_12545_));
 sky130_fd_sc_hd__a21oi_1 _20025_ (.A1(_12468_),
    .A2(_12543_),
    .B1(_12545_),
    .Y(_00168_));
 sky130_fd_sc_hd__mux2i_1 _20026_ (.A0(\cs_registers_i.pc_if_i[21] ),
    .A1(\cs_registers_i.pc_id_i[21] ),
    .S(_12498_),
    .Y(_12546_));
 sky130_fd_sc_hd__nor2_1 _20027_ (.A(_11623_),
    .B(_12501_),
    .Y(_12547_));
 sky130_fd_sc_hd__a211oi_1 _20028_ (.A1(\cs_registers_i.csr_depc_o[21] ),
    .A2(_12501_),
    .B1(_12547_),
    .C1(_12468_),
    .Y(_12548_));
 sky130_fd_sc_hd__a21oi_1 _20029_ (.A1(_12468_),
    .A2(_12546_),
    .B1(_12548_),
    .Y(_00169_));
 sky130_fd_sc_hd__mux2i_2 _20030_ (.A0(\cs_registers_i.pc_if_i[22] ),
    .A1(\cs_registers_i.pc_id_i[22] ),
    .S(_12498_),
    .Y(_12549_));
 sky130_fd_sc_hd__nor2_1 _20031_ (.A(_11643_),
    .B(_12501_),
    .Y(_12550_));
 sky130_fd_sc_hd__a211oi_1 _20032_ (.A1(\cs_registers_i.csr_depc_o[22] ),
    .A2(_12501_),
    .B1(_12550_),
    .C1(_12468_),
    .Y(_12551_));
 sky130_fd_sc_hd__a21oi_1 _20033_ (.A1(_12468_),
    .A2(_12549_),
    .B1(_12551_),
    .Y(_00170_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_616 ();
 sky130_fd_sc_hd__mux2i_2 _20035_ (.A0(\cs_registers_i.pc_if_i[23] ),
    .A1(\cs_registers_i.pc_id_i[23] ),
    .S(_12498_),
    .Y(_12553_));
 sky130_fd_sc_hd__nor2_1 _20036_ (.A(_11664_),
    .B(_12501_),
    .Y(_12554_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_615 ();
 sky130_fd_sc_hd__a211oi_1 _20038_ (.A1(\cs_registers_i.csr_depc_o[23] ),
    .A2(_12501_),
    .B1(_12554_),
    .C1(_12468_),
    .Y(_12556_));
 sky130_fd_sc_hd__a21oi_1 _20039_ (.A1(_12468_),
    .A2(_12553_),
    .B1(_12556_),
    .Y(_00171_));
 sky130_fd_sc_hd__mux2i_4 _20040_ (.A0(\cs_registers_i.pc_if_i[24] ),
    .A1(\cs_registers_i.pc_id_i[24] ),
    .S(_12498_),
    .Y(_12557_));
 sky130_fd_sc_hd__nor2_1 _20041_ (.A(_11684_),
    .B(_12501_),
    .Y(_12558_));
 sky130_fd_sc_hd__a211oi_1 _20042_ (.A1(\cs_registers_i.csr_depc_o[24] ),
    .A2(_12501_),
    .B1(_12558_),
    .C1(_12468_),
    .Y(_12559_));
 sky130_fd_sc_hd__a21oi_1 _20043_ (.A1(_12468_),
    .A2(_12557_),
    .B1(_12559_),
    .Y(_00172_));
 sky130_fd_sc_hd__mux2i_2 _20044_ (.A0(\cs_registers_i.pc_if_i[25] ),
    .A1(\cs_registers_i.pc_id_i[25] ),
    .S(_12498_),
    .Y(_12560_));
 sky130_fd_sc_hd__nor2_1 _20045_ (.A(_11706_),
    .B(_12501_),
    .Y(_12561_));
 sky130_fd_sc_hd__a211oi_1 _20046_ (.A1(\cs_registers_i.csr_depc_o[25] ),
    .A2(_12501_),
    .B1(_12561_),
    .C1(_12468_),
    .Y(_12562_));
 sky130_fd_sc_hd__a21oi_1 _20047_ (.A1(_12468_),
    .A2(_12560_),
    .B1(_12562_),
    .Y(_00173_));
 sky130_fd_sc_hd__mux2i_2 _20048_ (.A0(\cs_registers_i.pc_if_i[26] ),
    .A1(\cs_registers_i.pc_id_i[26] ),
    .S(_12498_),
    .Y(_12563_));
 sky130_fd_sc_hd__nor2_1 _20049_ (.A(_11726_),
    .B(_12501_),
    .Y(_12564_));
 sky130_fd_sc_hd__a211oi_1 _20050_ (.A1(\cs_registers_i.csr_depc_o[26] ),
    .A2(_12501_),
    .B1(_12564_),
    .C1(_12468_),
    .Y(_12565_));
 sky130_fd_sc_hd__a21oi_1 _20051_ (.A1(_12468_),
    .A2(_12563_),
    .B1(_12565_),
    .Y(_00174_));
 sky130_fd_sc_hd__mux2i_4 _20052_ (.A0(\cs_registers_i.pc_if_i[27] ),
    .A1(\cs_registers_i.pc_id_i[27] ),
    .S(_12498_),
    .Y(_12566_));
 sky130_fd_sc_hd__nor2_1 _20053_ (.A(_11746_),
    .B(_12501_),
    .Y(_12567_));
 sky130_fd_sc_hd__a211oi_1 _20054_ (.A1(\cs_registers_i.csr_depc_o[27] ),
    .A2(_12501_),
    .B1(_12567_),
    .C1(_12468_),
    .Y(_12568_));
 sky130_fd_sc_hd__a21oi_1 _20055_ (.A1(_12468_),
    .A2(_12566_),
    .B1(_12568_),
    .Y(_00175_));
 sky130_fd_sc_hd__mux2i_4 _20056_ (.A0(\cs_registers_i.pc_if_i[28] ),
    .A1(\cs_registers_i.pc_id_i[28] ),
    .S(_12498_),
    .Y(_12569_));
 sky130_fd_sc_hd__nor2_1 _20057_ (.A(_11765_),
    .B(_12501_),
    .Y(_12570_));
 sky130_fd_sc_hd__a211oi_1 _20058_ (.A1(\cs_registers_i.csr_depc_o[28] ),
    .A2(_12501_),
    .B1(_12570_),
    .C1(_12468_),
    .Y(_12571_));
 sky130_fd_sc_hd__a21oi_1 _20059_ (.A1(_12468_),
    .A2(_12569_),
    .B1(_12571_),
    .Y(_00176_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_614 ();
 sky130_fd_sc_hd__mux2i_2 _20061_ (.A0(\cs_registers_i.pc_if_i[29] ),
    .A1(\cs_registers_i.pc_id_i[29] ),
    .S(_12498_),
    .Y(_12573_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_612 ();
 sky130_fd_sc_hd__nor2_1 _20064_ (.A(_11785_),
    .B(_12501_),
    .Y(_12576_));
 sky130_fd_sc_hd__a211oi_1 _20065_ (.A1(\cs_registers_i.csr_depc_o[29] ),
    .A2(_12501_),
    .B1(_12576_),
    .C1(_12468_),
    .Y(_12577_));
 sky130_fd_sc_hd__a21oi_1 _20066_ (.A1(_12468_),
    .A2(_12573_),
    .B1(_12577_),
    .Y(_00177_));
 sky130_fd_sc_hd__mux2i_2 _20067_ (.A0(\cs_registers_i.pc_if_i[2] ),
    .A1(\cs_registers_i.pc_id_i[2] ),
    .S(_12498_),
    .Y(_12578_));
 sky130_fd_sc_hd__nor2_1 _20068_ (.A(_11309_),
    .B(_12501_),
    .Y(_12579_));
 sky130_fd_sc_hd__a211oi_1 _20069_ (.A1(\cs_registers_i.csr_depc_o[2] ),
    .A2(_12501_),
    .B1(_12579_),
    .C1(_12468_),
    .Y(_12580_));
 sky130_fd_sc_hd__a21oi_1 _20070_ (.A1(_12468_),
    .A2(_12578_),
    .B1(_12580_),
    .Y(_00178_));
 sky130_fd_sc_hd__mux2i_1 _20071_ (.A0(\cs_registers_i.pc_if_i[30] ),
    .A1(\cs_registers_i.pc_id_i[30] ),
    .S(_12498_),
    .Y(_12581_));
 sky130_fd_sc_hd__nor2_1 _20072_ (.A(_11808_),
    .B(_12501_),
    .Y(_12582_));
 sky130_fd_sc_hd__a211oi_1 _20073_ (.A1(\cs_registers_i.csr_depc_o[30] ),
    .A2(_12501_),
    .B1(_12582_),
    .C1(_12468_),
    .Y(_12583_));
 sky130_fd_sc_hd__a21oi_1 _20074_ (.A1(_12468_),
    .A2(_12581_),
    .B1(_12583_),
    .Y(_00179_));
 sky130_fd_sc_hd__mux2i_1 _20075_ (.A0(\cs_registers_i.pc_if_i[31] ),
    .A1(\cs_registers_i.pc_id_i[31] ),
    .S(_12498_),
    .Y(_12584_));
 sky130_fd_sc_hd__nor2_1 _20076_ (.A(_11826_),
    .B(_12501_),
    .Y(_12585_));
 sky130_fd_sc_hd__a211oi_1 _20077_ (.A1(\cs_registers_i.csr_depc_o[31] ),
    .A2(_12501_),
    .B1(_12585_),
    .C1(_12468_),
    .Y(_12586_));
 sky130_fd_sc_hd__a21oi_1 _20078_ (.A1(_12468_),
    .A2(_12584_),
    .B1(_12586_),
    .Y(_00180_));
 sky130_fd_sc_hd__mux2i_4 _20079_ (.A0(\cs_registers_i.pc_if_i[3] ),
    .A1(\cs_registers_i.pc_id_i[3] ),
    .S(_12498_),
    .Y(_12587_));
 sky130_fd_sc_hd__nor2_1 _20080_ (.A(_11867_),
    .B(_12501_),
    .Y(_12588_));
 sky130_fd_sc_hd__a211oi_1 _20081_ (.A1(\cs_registers_i.csr_depc_o[3] ),
    .A2(_12501_),
    .B1(_12588_),
    .C1(_12468_),
    .Y(_12589_));
 sky130_fd_sc_hd__a21oi_1 _20082_ (.A1(_12468_),
    .A2(_12587_),
    .B1(_12589_),
    .Y(_00181_));
 sky130_fd_sc_hd__mux2i_2 _20083_ (.A0(\cs_registers_i.pc_if_i[4] ),
    .A1(\cs_registers_i.pc_id_i[4] ),
    .S(_12498_),
    .Y(_12590_));
 sky130_fd_sc_hd__nor2_1 _20084_ (.A(_11887_),
    .B(_12501_),
    .Y(_12591_));
 sky130_fd_sc_hd__a211oi_1 _20085_ (.A1(\cs_registers_i.csr_depc_o[4] ),
    .A2(_12501_),
    .B1(_12591_),
    .C1(_12468_),
    .Y(_12592_));
 sky130_fd_sc_hd__a21oi_1 _20086_ (.A1(_12468_),
    .A2(_12590_),
    .B1(_12592_),
    .Y(_00182_));
 sky130_fd_sc_hd__mux2i_2 _20087_ (.A0(\cs_registers_i.pc_if_i[5] ),
    .A1(\cs_registers_i.pc_id_i[5] ),
    .S(_12498_),
    .Y(_12593_));
 sky130_fd_sc_hd__a21oi_2 _20088_ (.A1(net952),
    .A2(_11148_),
    .B1(_11901_),
    .Y(_12594_));
 sky130_fd_sc_hd__nor2_1 _20089_ (.A(_12594_),
    .B(_12501_),
    .Y(_12595_));
 sky130_fd_sc_hd__a211oi_1 _20090_ (.A1(\cs_registers_i.csr_depc_o[5] ),
    .A2(_12501_),
    .B1(_12595_),
    .C1(_12468_),
    .Y(_12596_));
 sky130_fd_sc_hd__a21oi_1 _20091_ (.A1(_12468_),
    .A2(_12593_),
    .B1(_12596_),
    .Y(_00183_));
 sky130_fd_sc_hd__mux2i_1 _20092_ (.A0(\cs_registers_i.pc_if_i[6] ),
    .A1(\cs_registers_i.pc_id_i[6] ),
    .S(_12498_),
    .Y(_12597_));
 sky130_fd_sc_hd__nor2_1 _20093_ (.A(_12113_),
    .B(_12501_),
    .Y(_12598_));
 sky130_fd_sc_hd__a211oi_1 _20094_ (.A1(\cs_registers_i.csr_depc_o[6] ),
    .A2(_12501_),
    .B1(_12598_),
    .C1(_12468_),
    .Y(_12599_));
 sky130_fd_sc_hd__a21oi_1 _20095_ (.A1(_12468_),
    .A2(_12597_),
    .B1(_12599_),
    .Y(_00184_));
 sky130_fd_sc_hd__mux2i_2 _20096_ (.A0(\cs_registers_i.pc_if_i[7] ),
    .A1(\cs_registers_i.pc_id_i[7] ),
    .S(_12498_),
    .Y(_12600_));
 sky130_fd_sc_hd__nor2_1 _20097_ (.A(_11935_),
    .B(_12501_),
    .Y(_12601_));
 sky130_fd_sc_hd__a211oi_1 _20098_ (.A1(\cs_registers_i.csr_depc_o[7] ),
    .A2(_12501_),
    .B1(_12601_),
    .C1(_12468_),
    .Y(_12602_));
 sky130_fd_sc_hd__a21oi_1 _20099_ (.A1(_12468_),
    .A2(_12600_),
    .B1(_12602_),
    .Y(_00185_));
 sky130_fd_sc_hd__mux2i_1 _20100_ (.A0(\cs_registers_i.pc_if_i[8] ),
    .A1(\cs_registers_i.pc_id_i[8] ),
    .S(_12498_),
    .Y(_12603_));
 sky130_fd_sc_hd__nor2_1 _20101_ (.A(_11957_),
    .B(_12501_),
    .Y(_12604_));
 sky130_fd_sc_hd__a211oi_1 _20102_ (.A1(\cs_registers_i.csr_depc_o[8] ),
    .A2(_12501_),
    .B1(_12604_),
    .C1(_12468_),
    .Y(_12605_));
 sky130_fd_sc_hd__a21oi_1 _20103_ (.A1(_12468_),
    .A2(_12603_),
    .B1(_12605_),
    .Y(_00186_));
 sky130_fd_sc_hd__mux2i_1 _20104_ (.A0(\cs_registers_i.pc_if_i[9] ),
    .A1(\cs_registers_i.pc_id_i[9] ),
    .S(_12498_),
    .Y(_12606_));
 sky130_fd_sc_hd__nor2_1 _20105_ (.A(_11973_),
    .B(_12501_),
    .Y(_12607_));
 sky130_fd_sc_hd__a211oi_1 _20106_ (.A1(\cs_registers_i.csr_depc_o[9] ),
    .A2(_12501_),
    .B1(_12607_),
    .C1(_12468_),
    .Y(_12608_));
 sky130_fd_sc_hd__a21oi_1 _20107_ (.A1(_12468_),
    .A2(_12606_),
    .B1(_12608_),
    .Y(_00187_));
 sky130_fd_sc_hd__nand2_8 _20108_ (.A(net271),
    .B(_11252_),
    .Y(_12609_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_610 ();
 sky130_fd_sc_hd__nand2_1 _20111_ (.A(\cs_registers_i.dscratch0_q[0] ),
    .B(_12609_),
    .Y(_12612_));
 sky130_fd_sc_hd__o21ai_0 _20112_ (.A1(_11280_),
    .A2(_12609_),
    .B1(_12612_),
    .Y(_00188_));
 sky130_fd_sc_hd__mux2_1 _20113_ (.A0(_11357_),
    .A1(\cs_registers_i.dscratch0_q[10] ),
    .S(_12609_),
    .X(_00189_));
 sky130_fd_sc_hd__nand2_1 _20114_ (.A(\cs_registers_i.dscratch0_q[11] ),
    .B(_12609_),
    .Y(_12613_));
 sky130_fd_sc_hd__o21ai_0 _20115_ (.A1(_12481_),
    .A2(_12609_),
    .B1(_12613_),
    .Y(_00190_));
 sky130_fd_sc_hd__nand2_1 _20116_ (.A(\cs_registers_i.dscratch0_q[12] ),
    .B(_12609_),
    .Y(_12614_));
 sky130_fd_sc_hd__o21ai_0 _20117_ (.A1(_11428_),
    .A2(_12609_),
    .B1(_12614_),
    .Y(_00191_));
 sky130_fd_sc_hd__nand2_1 _20118_ (.A(\cs_registers_i.dscratch0_q[13] ),
    .B(_12609_),
    .Y(_12615_));
 sky130_fd_sc_hd__o21ai_0 _20119_ (.A1(_11448_),
    .A2(_12609_),
    .B1(_12615_),
    .Y(_00192_));
 sky130_fd_sc_hd__nand2_1 _20120_ (.A(\cs_registers_i.dscratch0_q[14] ),
    .B(_12609_),
    .Y(_12616_));
 sky130_fd_sc_hd__o21ai_0 _20121_ (.A1(_11465_),
    .A2(_12609_),
    .B1(_12616_),
    .Y(_00193_));
 sky130_fd_sc_hd__nand2_1 _20122_ (.A(\cs_registers_i.dscratch0_q[15] ),
    .B(_12609_),
    .Y(_12617_));
 sky130_fd_sc_hd__o21ai_0 _20123_ (.A1(_11488_),
    .A2(_12609_),
    .B1(_12617_),
    .Y(_00194_));
 sky130_fd_sc_hd__nand2_1 _20124_ (.A(\cs_registers_i.dscratch0_q[16] ),
    .B(_12609_),
    .Y(_12618_));
 sky130_fd_sc_hd__o21ai_0 _20125_ (.A1(_11505_),
    .A2(_12609_),
    .B1(_12618_),
    .Y(_00195_));
 sky130_fd_sc_hd__nand2_1 _20126_ (.A(\cs_registers_i.dscratch0_q[17] ),
    .B(_12609_),
    .Y(_12619_));
 sky130_fd_sc_hd__o21ai_0 _20127_ (.A1(_11523_),
    .A2(_12609_),
    .B1(_12619_),
    .Y(_00196_));
 sky130_fd_sc_hd__nand2_1 _20128_ (.A(\cs_registers_i.dscratch0_q[18] ),
    .B(_12609_),
    .Y(_12620_));
 sky130_fd_sc_hd__o21ai_0 _20129_ (.A1(_11546_),
    .A2(_12609_),
    .B1(_12620_),
    .Y(_00197_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_609 ();
 sky130_fd_sc_hd__nand2_1 _20131_ (.A(\cs_registers_i.dscratch0_q[19] ),
    .B(_12609_),
    .Y(_12622_));
 sky130_fd_sc_hd__o21ai_0 _20132_ (.A1(_11563_),
    .A2(_12609_),
    .B1(_12622_),
    .Y(_00198_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_608 ();
 sky130_fd_sc_hd__nand2_1 _20134_ (.A(\cs_registers_i.dscratch0_q[1] ),
    .B(_12609_),
    .Y(_12624_));
 sky130_fd_sc_hd__o21ai_0 _20135_ (.A1(_11582_),
    .A2(_12609_),
    .B1(_12624_),
    .Y(_00199_));
 sky130_fd_sc_hd__nand2_1 _20136_ (.A(\cs_registers_i.dscratch0_q[20] ),
    .B(_12609_),
    .Y(_12625_));
 sky130_fd_sc_hd__o21ai_0 _20137_ (.A1(_11599_),
    .A2(_12609_),
    .B1(_12625_),
    .Y(_00200_));
 sky130_fd_sc_hd__nand2_1 _20138_ (.A(\cs_registers_i.dscratch0_q[21] ),
    .B(_12609_),
    .Y(_12626_));
 sky130_fd_sc_hd__o21ai_0 _20139_ (.A1(_11623_),
    .A2(_12609_),
    .B1(_12626_),
    .Y(_00201_));
 sky130_fd_sc_hd__nand2_1 _20140_ (.A(\cs_registers_i.dscratch0_q[22] ),
    .B(_12609_),
    .Y(_12627_));
 sky130_fd_sc_hd__o21ai_0 _20141_ (.A1(_11643_),
    .A2(_12609_),
    .B1(_12627_),
    .Y(_00202_));
 sky130_fd_sc_hd__nand2_1 _20142_ (.A(\cs_registers_i.dscratch0_q[23] ),
    .B(_12609_),
    .Y(_12628_));
 sky130_fd_sc_hd__o21ai_0 _20143_ (.A1(_11664_),
    .A2(_12609_),
    .B1(_12628_),
    .Y(_00203_));
 sky130_fd_sc_hd__nand2_1 _20144_ (.A(\cs_registers_i.dscratch0_q[24] ),
    .B(_12609_),
    .Y(_12629_));
 sky130_fd_sc_hd__o21ai_0 _20145_ (.A1(_11684_),
    .A2(_12609_),
    .B1(_12629_),
    .Y(_00204_));
 sky130_fd_sc_hd__nand2_1 _20146_ (.A(\cs_registers_i.dscratch0_q[25] ),
    .B(_12609_),
    .Y(_12630_));
 sky130_fd_sc_hd__o21ai_0 _20147_ (.A1(_11706_),
    .A2(_12609_),
    .B1(_12630_),
    .Y(_00205_));
 sky130_fd_sc_hd__nand2_1 _20148_ (.A(\cs_registers_i.dscratch0_q[26] ),
    .B(_12609_),
    .Y(_12631_));
 sky130_fd_sc_hd__o21ai_0 _20149_ (.A1(_11726_),
    .A2(_12609_),
    .B1(_12631_),
    .Y(_00206_));
 sky130_fd_sc_hd__nand2_1 _20150_ (.A(\cs_registers_i.dscratch0_q[27] ),
    .B(_12609_),
    .Y(_12632_));
 sky130_fd_sc_hd__o21ai_0 _20151_ (.A1(_11746_),
    .A2(_12609_),
    .B1(_12632_),
    .Y(_00207_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_607 ();
 sky130_fd_sc_hd__nand2_1 _20153_ (.A(\cs_registers_i.dscratch0_q[28] ),
    .B(_12609_),
    .Y(_12634_));
 sky130_fd_sc_hd__o21ai_0 _20154_ (.A1(_11765_),
    .A2(_12609_),
    .B1(_12634_),
    .Y(_00208_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_606 ();
 sky130_fd_sc_hd__nand2_1 _20156_ (.A(\cs_registers_i.dscratch0_q[29] ),
    .B(_12609_),
    .Y(_12636_));
 sky130_fd_sc_hd__o21ai_0 _20157_ (.A1(_11785_),
    .A2(_12609_),
    .B1(_12636_),
    .Y(_00209_));
 sky130_fd_sc_hd__nand2_1 _20158_ (.A(\cs_registers_i.dscratch0_q[2] ),
    .B(_12609_),
    .Y(_12637_));
 sky130_fd_sc_hd__o21ai_0 _20159_ (.A1(_11309_),
    .A2(_12609_),
    .B1(_12637_),
    .Y(_00210_));
 sky130_fd_sc_hd__nand2_1 _20160_ (.A(\cs_registers_i.dscratch0_q[30] ),
    .B(_12609_),
    .Y(_12638_));
 sky130_fd_sc_hd__o21ai_0 _20161_ (.A1(_11808_),
    .A2(_12609_),
    .B1(_12638_),
    .Y(_00211_));
 sky130_fd_sc_hd__nand2_1 _20162_ (.A(\cs_registers_i.dscratch0_q[31] ),
    .B(_12609_),
    .Y(_12639_));
 sky130_fd_sc_hd__o21ai_0 _20163_ (.A1(_11826_),
    .A2(_12609_),
    .B1(_12639_),
    .Y(_00212_));
 sky130_fd_sc_hd__nand2_1 _20164_ (.A(\cs_registers_i.dscratch0_q[3] ),
    .B(_12609_),
    .Y(_12640_));
 sky130_fd_sc_hd__o21ai_0 _20165_ (.A1(_11867_),
    .A2(_12609_),
    .B1(_12640_),
    .Y(_00213_));
 sky130_fd_sc_hd__nand2_1 _20166_ (.A(\cs_registers_i.dscratch0_q[4] ),
    .B(_12609_),
    .Y(_12641_));
 sky130_fd_sc_hd__o21ai_0 _20167_ (.A1(_11887_),
    .A2(_12609_),
    .B1(_12641_),
    .Y(_00214_));
 sky130_fd_sc_hd__nand2_1 _20168_ (.A(\cs_registers_i.dscratch0_q[5] ),
    .B(_12609_),
    .Y(_12642_));
 sky130_fd_sc_hd__o21ai_0 _20169_ (.A1(_12594_),
    .A2(_12609_),
    .B1(_12642_),
    .Y(_00215_));
 sky130_fd_sc_hd__nand2_1 _20170_ (.A(\cs_registers_i.dscratch0_q[6] ),
    .B(_12609_),
    .Y(_12643_));
 sky130_fd_sc_hd__o21ai_0 _20171_ (.A1(_12113_),
    .A2(_12609_),
    .B1(_12643_),
    .Y(_00216_));
 sky130_fd_sc_hd__nand2_1 _20172_ (.A(\cs_registers_i.dscratch0_q[7] ),
    .B(_12609_),
    .Y(_12644_));
 sky130_fd_sc_hd__o21ai_0 _20173_ (.A1(_11935_),
    .A2(_12609_),
    .B1(_12644_),
    .Y(_00217_));
 sky130_fd_sc_hd__nand2_1 _20174_ (.A(\cs_registers_i.dscratch0_q[8] ),
    .B(_12609_),
    .Y(_12645_));
 sky130_fd_sc_hd__o21ai_0 _20175_ (.A1(_11957_),
    .A2(_12609_),
    .B1(_12645_),
    .Y(_00218_));
 sky130_fd_sc_hd__nand2_1 _20176_ (.A(\cs_registers_i.dscratch0_q[9] ),
    .B(_12609_),
    .Y(_12646_));
 sky130_fd_sc_hd__o21ai_0 _20177_ (.A1(_11973_),
    .A2(_12609_),
    .B1(_12646_),
    .Y(_00219_));
 sky130_fd_sc_hd__nand2_8 _20178_ (.A(net271),
    .B(_11260_),
    .Y(_12647_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_604 ();
 sky130_fd_sc_hd__nand2_1 _20181_ (.A(\cs_registers_i.dscratch1_q[0] ),
    .B(_12647_),
    .Y(_12650_));
 sky130_fd_sc_hd__o21ai_0 _20182_ (.A1(_11280_),
    .A2(_12647_),
    .B1(_12650_),
    .Y(_00220_));
 sky130_fd_sc_hd__mux2_1 _20183_ (.A0(_11357_),
    .A1(\cs_registers_i.dscratch1_q[10] ),
    .S(_12647_),
    .X(_00221_));
 sky130_fd_sc_hd__nand2_1 _20184_ (.A(\cs_registers_i.dscratch1_q[11] ),
    .B(_12647_),
    .Y(_12651_));
 sky130_fd_sc_hd__o21ai_0 _20185_ (.A1(_12481_),
    .A2(_12647_),
    .B1(_12651_),
    .Y(_00222_));
 sky130_fd_sc_hd__nand2_1 _20186_ (.A(\cs_registers_i.dscratch1_q[12] ),
    .B(_12647_),
    .Y(_12652_));
 sky130_fd_sc_hd__o21ai_0 _20187_ (.A1(_11428_),
    .A2(_12647_),
    .B1(_12652_),
    .Y(_00223_));
 sky130_fd_sc_hd__nand2_1 _20188_ (.A(\cs_registers_i.dscratch1_q[13] ),
    .B(_12647_),
    .Y(_12653_));
 sky130_fd_sc_hd__o21ai_0 _20189_ (.A1(_11448_),
    .A2(_12647_),
    .B1(_12653_),
    .Y(_00224_));
 sky130_fd_sc_hd__nand2_1 _20190_ (.A(\cs_registers_i.dscratch1_q[14] ),
    .B(_12647_),
    .Y(_12654_));
 sky130_fd_sc_hd__o21ai_0 _20191_ (.A1(_11465_),
    .A2(_12647_),
    .B1(_12654_),
    .Y(_00225_));
 sky130_fd_sc_hd__nand2_1 _20192_ (.A(\cs_registers_i.dscratch1_q[15] ),
    .B(_12647_),
    .Y(_12655_));
 sky130_fd_sc_hd__o21ai_0 _20193_ (.A1(_11488_),
    .A2(_12647_),
    .B1(_12655_),
    .Y(_00226_));
 sky130_fd_sc_hd__nand2_1 _20194_ (.A(\cs_registers_i.dscratch1_q[16] ),
    .B(_12647_),
    .Y(_12656_));
 sky130_fd_sc_hd__o21ai_0 _20195_ (.A1(_11505_),
    .A2(_12647_),
    .B1(_12656_),
    .Y(_00227_));
 sky130_fd_sc_hd__nand2_1 _20196_ (.A(\cs_registers_i.dscratch1_q[17] ),
    .B(_12647_),
    .Y(_12657_));
 sky130_fd_sc_hd__o21ai_0 _20197_ (.A1(_11523_),
    .A2(_12647_),
    .B1(_12657_),
    .Y(_00228_));
 sky130_fd_sc_hd__nand2_1 _20198_ (.A(\cs_registers_i.dscratch1_q[18] ),
    .B(_12647_),
    .Y(_12658_));
 sky130_fd_sc_hd__o21ai_0 _20199_ (.A1(_11546_),
    .A2(_12647_),
    .B1(_12658_),
    .Y(_00229_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_603 ();
 sky130_fd_sc_hd__nand2_1 _20201_ (.A(\cs_registers_i.dscratch1_q[19] ),
    .B(_12647_),
    .Y(_12660_));
 sky130_fd_sc_hd__o21ai_0 _20202_ (.A1(_11563_),
    .A2(_12647_),
    .B1(_12660_),
    .Y(_00230_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_602 ();
 sky130_fd_sc_hd__nand2_1 _20204_ (.A(\cs_registers_i.dscratch1_q[1] ),
    .B(_12647_),
    .Y(_12662_));
 sky130_fd_sc_hd__o21ai_0 _20205_ (.A1(_11582_),
    .A2(_12647_),
    .B1(_12662_),
    .Y(_00231_));
 sky130_fd_sc_hd__nand2_1 _20206_ (.A(\cs_registers_i.dscratch1_q[20] ),
    .B(_12647_),
    .Y(_12663_));
 sky130_fd_sc_hd__o21ai_0 _20207_ (.A1(_11599_),
    .A2(_12647_),
    .B1(_12663_),
    .Y(_00232_));
 sky130_fd_sc_hd__nand2_1 _20208_ (.A(\cs_registers_i.dscratch1_q[21] ),
    .B(_12647_),
    .Y(_12664_));
 sky130_fd_sc_hd__o21ai_0 _20209_ (.A1(_11623_),
    .A2(_12647_),
    .B1(_12664_),
    .Y(_00233_));
 sky130_fd_sc_hd__nand2_1 _20210_ (.A(\cs_registers_i.dscratch1_q[22] ),
    .B(_12647_),
    .Y(_12665_));
 sky130_fd_sc_hd__o21ai_0 _20211_ (.A1(_11643_),
    .A2(_12647_),
    .B1(_12665_),
    .Y(_00234_));
 sky130_fd_sc_hd__nand2_1 _20212_ (.A(\cs_registers_i.dscratch1_q[23] ),
    .B(_12647_),
    .Y(_12666_));
 sky130_fd_sc_hd__o21ai_0 _20213_ (.A1(_11664_),
    .A2(_12647_),
    .B1(_12666_),
    .Y(_00235_));
 sky130_fd_sc_hd__nand2_1 _20214_ (.A(\cs_registers_i.dscratch1_q[24] ),
    .B(_12647_),
    .Y(_12667_));
 sky130_fd_sc_hd__o21ai_0 _20215_ (.A1(_11684_),
    .A2(_12647_),
    .B1(_12667_),
    .Y(_00236_));
 sky130_fd_sc_hd__nand2_1 _20216_ (.A(\cs_registers_i.dscratch1_q[25] ),
    .B(_12647_),
    .Y(_12668_));
 sky130_fd_sc_hd__o21ai_0 _20217_ (.A1(_11706_),
    .A2(_12647_),
    .B1(_12668_),
    .Y(_00237_));
 sky130_fd_sc_hd__nand2_1 _20218_ (.A(\cs_registers_i.dscratch1_q[26] ),
    .B(_12647_),
    .Y(_12669_));
 sky130_fd_sc_hd__o21ai_0 _20219_ (.A1(_11726_),
    .A2(_12647_),
    .B1(_12669_),
    .Y(_00238_));
 sky130_fd_sc_hd__nand2_1 _20220_ (.A(\cs_registers_i.dscratch1_q[27] ),
    .B(_12647_),
    .Y(_12670_));
 sky130_fd_sc_hd__o21ai_0 _20221_ (.A1(_11746_),
    .A2(_12647_),
    .B1(_12670_),
    .Y(_00239_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_601 ();
 sky130_fd_sc_hd__nand2_1 _20223_ (.A(\cs_registers_i.dscratch1_q[28] ),
    .B(_12647_),
    .Y(_12672_));
 sky130_fd_sc_hd__o21ai_0 _20224_ (.A1(_11765_),
    .A2(_12647_),
    .B1(_12672_),
    .Y(_00240_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_600 ();
 sky130_fd_sc_hd__nand2_1 _20226_ (.A(\cs_registers_i.dscratch1_q[29] ),
    .B(_12647_),
    .Y(_12674_));
 sky130_fd_sc_hd__o21ai_0 _20227_ (.A1(_11785_),
    .A2(_12647_),
    .B1(_12674_),
    .Y(_00241_));
 sky130_fd_sc_hd__nand2_1 _20228_ (.A(\cs_registers_i.dscratch1_q[2] ),
    .B(_12647_),
    .Y(_12675_));
 sky130_fd_sc_hd__o21ai_0 _20229_ (.A1(_11309_),
    .A2(_12647_),
    .B1(_12675_),
    .Y(_00242_));
 sky130_fd_sc_hd__nand2_1 _20230_ (.A(\cs_registers_i.dscratch1_q[30] ),
    .B(_12647_),
    .Y(_12676_));
 sky130_fd_sc_hd__o21ai_0 _20231_ (.A1(_11808_),
    .A2(_12647_),
    .B1(_12676_),
    .Y(_00243_));
 sky130_fd_sc_hd__nand2_1 _20232_ (.A(\cs_registers_i.dscratch1_q[31] ),
    .B(_12647_),
    .Y(_12677_));
 sky130_fd_sc_hd__o21ai_0 _20233_ (.A1(_11826_),
    .A2(_12647_),
    .B1(_12677_),
    .Y(_00244_));
 sky130_fd_sc_hd__nand2_1 _20234_ (.A(\cs_registers_i.dscratch1_q[3] ),
    .B(_12647_),
    .Y(_12678_));
 sky130_fd_sc_hd__o21ai_0 _20235_ (.A1(_11867_),
    .A2(_12647_),
    .B1(_12678_),
    .Y(_00245_));
 sky130_fd_sc_hd__nand2_1 _20236_ (.A(\cs_registers_i.dscratch1_q[4] ),
    .B(_12647_),
    .Y(_12679_));
 sky130_fd_sc_hd__o21ai_0 _20237_ (.A1(_11887_),
    .A2(_12647_),
    .B1(_12679_),
    .Y(_00246_));
 sky130_fd_sc_hd__nand2_1 _20238_ (.A(\cs_registers_i.dscratch1_q[5] ),
    .B(_12647_),
    .Y(_12680_));
 sky130_fd_sc_hd__o21ai_0 _20239_ (.A1(_12594_),
    .A2(_12647_),
    .B1(_12680_),
    .Y(_00247_));
 sky130_fd_sc_hd__nand2_1 _20240_ (.A(\cs_registers_i.dscratch1_q[6] ),
    .B(_12647_),
    .Y(_12681_));
 sky130_fd_sc_hd__o21ai_0 _20241_ (.A1(_12113_),
    .A2(_12647_),
    .B1(_12681_),
    .Y(_00248_));
 sky130_fd_sc_hd__nand2_1 _20242_ (.A(\cs_registers_i.dscratch1_q[7] ),
    .B(_12647_),
    .Y(_12682_));
 sky130_fd_sc_hd__o21ai_0 _20243_ (.A1(_11935_),
    .A2(_12647_),
    .B1(_12682_),
    .Y(_00249_));
 sky130_fd_sc_hd__nand2_1 _20244_ (.A(\cs_registers_i.dscratch1_q[8] ),
    .B(_12647_),
    .Y(_12683_));
 sky130_fd_sc_hd__o21ai_0 _20245_ (.A1(_11957_),
    .A2(_12647_),
    .B1(_12683_),
    .Y(_00250_));
 sky130_fd_sc_hd__nand2_1 _20246_ (.A(\cs_registers_i.dscratch1_q[9] ),
    .B(_12647_),
    .Y(_12684_));
 sky130_fd_sc_hd__o21ai_0 _20247_ (.A1(_11973_),
    .A2(_12647_),
    .B1(_12684_),
    .Y(_00251_));
 sky130_fd_sc_hd__nor3_4 _20248_ (.A(\cs_registers_i.debug_mode_i ),
    .B(_12468_),
    .C(_12471_),
    .Y(_12685_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_599 ();
 sky130_fd_sc_hd__nor3_4 _20250_ (.A(_11032_),
    .B(_12450_),
    .C(_12451_),
    .Y(_12687_));
 sky130_fd_sc_hd__nor2_8 _20251_ (.A(net282),
    .B(_12687_),
    .Y(_12688_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_598 ();
 sky130_fd_sc_hd__nand2_8 _20253_ (.A(\cs_registers_i.nmi_mode_i ),
    .B(_12455_),
    .Y(_12690_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_597 ();
 sky130_fd_sc_hd__nor2_1 _20255_ (.A(\id_stage_i.controller_i.store_err_q ),
    .B(\id_stage_i.controller_i.load_err_q ),
    .Y(_12692_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_596 ();
 sky130_fd_sc_hd__a211oi_4 _20257_ (.A1(\id_stage_i.controller_i.instr_valid_i ),
    .A2(_10947_),
    .B1(_12692_),
    .C1(\id_stage_i.controller_i.illegal_insn_q ),
    .Y(_12694_));
 sky130_fd_sc_hd__nor3_1 _20258_ (.A(net372),
    .B(_08160_),
    .C(_08163_),
    .Y(_12695_));
 sky130_fd_sc_hd__nor4_1 _20259_ (.A(net382),
    .B(net553),
    .C(\id_stage_i.controller_i.instr_fetch_err_i ),
    .D(\id_stage_i.controller_i.illegal_insn_q ),
    .Y(_12696_));
 sky130_fd_sc_hd__nand4_1 _20260_ (.A(_12695_),
    .B(_11000_),
    .C(_10937_),
    .D(_12696_),
    .Y(_12697_));
 sky130_fd_sc_hd__o31ai_1 _20261_ (.A1(\cs_registers_i.debug_mode_i ),
    .A2(_10998_),
    .A3(_11002_),
    .B1(_12697_),
    .Y(_12698_));
 sky130_fd_sc_hd__o31ai_1 _20262_ (.A1(_11040_),
    .A2(_12694_),
    .A3(_12698_),
    .B1(_12469_),
    .Y(_12699_));
 sky130_fd_sc_hd__nand2_1 _20263_ (.A(\cs_registers_i.mie_q[8] ),
    .B(net143),
    .Y(_12700_));
 sky130_fd_sc_hd__nand2_1 _20264_ (.A(\cs_registers_i.mie_q[2] ),
    .B(net137),
    .Y(_12701_));
 sky130_fd_sc_hd__a32oi_1 _20265_ (.A1(\cs_registers_i.mie_q[1] ),
    .A2(net136),
    .A3(_12701_),
    .B1(net138),
    .B2(\cs_registers_i.mie_q[3] ),
    .Y(_12702_));
 sky130_fd_sc_hd__a21oi_1 _20266_ (.A1(\cs_registers_i.mie_q[4] ),
    .A2(net139),
    .B1(_12702_),
    .Y(_12703_));
 sky130_fd_sc_hd__a21oi_1 _20267_ (.A1(\cs_registers_i.mie_q[5] ),
    .A2(net140),
    .B1(_12703_),
    .Y(_12704_));
 sky130_fd_sc_hd__nand2_1 _20268_ (.A(\cs_registers_i.mie_q[7] ),
    .B(net142),
    .Y(_12705_));
 sky130_fd_sc_hd__o21ai_1 _20269_ (.A1(_11014_),
    .A2(_12704_),
    .B1(_12705_),
    .Y(_12706_));
 sky130_fd_sc_hd__a22oi_1 _20270_ (.A1(\cs_registers_i.mie_q[9] ),
    .A2(net144),
    .B1(_12700_),
    .B2(_12706_),
    .Y(_12707_));
 sky130_fd_sc_hd__a21oi_1 _20271_ (.A1(\cs_registers_i.mie_q[10] ),
    .A2(net131),
    .B1(_12707_),
    .Y(_12708_));
 sky130_fd_sc_hd__o21ai_1 _20272_ (.A1(_11022_),
    .A2(_12708_),
    .B1(_11020_),
    .Y(_12709_));
 sky130_fd_sc_hd__a21oi_4 _20273_ (.A1(_11019_),
    .A2(_12709_),
    .B1(_11012_),
    .Y(_12710_));
 sky130_fd_sc_hd__nor2b_2 _20274_ (.A(\cs_registers_i.nmi_mode_i ),
    .B_N(net145),
    .Y(_12711_));
 sky130_fd_sc_hd__o31ai_4 _20275_ (.A1(_11026_),
    .A2(_12710_),
    .A3(_12711_),
    .B1(_11034_),
    .Y(_12712_));
 sky130_fd_sc_hd__nand3_1 _20276_ (.A(net282),
    .B(_12699_),
    .C(_12712_),
    .Y(_12713_));
 sky130_fd_sc_hd__o21ai_0 _20277_ (.A1(\cs_registers_i.mstack_cause_q[0] ),
    .A2(_12690_),
    .B1(_12713_),
    .Y(_12714_));
 sky130_fd_sc_hd__a21oi_1 _20278_ (.A1(_11280_),
    .A2(_12688_),
    .B1(_12714_),
    .Y(_12715_));
 sky130_fd_sc_hd__nand2_1 _20279_ (.A(_11243_),
    .B(_11271_),
    .Y(_12716_));
 sky130_fd_sc_hd__nand2_4 _20280_ (.A(_12688_),
    .B(_12716_),
    .Y(_12717_));
 sky130_fd_sc_hd__mux2_1 _20281_ (.A0(\cs_registers_i.mcause_q[0] ),
    .A1(_12715_),
    .S(_12717_),
    .X(_00252_));
 sky130_fd_sc_hd__inv_1 _20282_ (.A(\cs_registers_i.mcause_q[1] ),
    .Y(_12718_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_594 ();
 sky130_fd_sc_hd__nand2_1 _20285_ (.A(_11582_),
    .B(_12688_),
    .Y(_12721_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_593 ();
 sky130_fd_sc_hd__or3_1 _20287_ (.A(_11012_),
    .B(_11018_),
    .C(_11025_),
    .X(_12723_));
 sky130_fd_sc_hd__nand2b_1 _20288_ (.A_N(_11016_),
    .B(_11013_),
    .Y(_12724_));
 sky130_fd_sc_hd__a222oi_1 _20289_ (.A1(\cs_registers_i.mie_q[8] ),
    .A2(net143),
    .B1(\cs_registers_i.mie_q[9] ),
    .B2(net144),
    .C1(_11015_),
    .C2(_12724_),
    .Y(_12725_));
 sky130_fd_sc_hd__o21ai_2 _20290_ (.A1(_11023_),
    .A2(_12725_),
    .B1(_11021_),
    .Y(_12726_));
 sky130_fd_sc_hd__nor2_1 _20291_ (.A(_11012_),
    .B(_12711_),
    .Y(_12727_));
 sky130_fd_sc_hd__nand3_1 _20292_ (.A(_12723_),
    .B(_12726_),
    .C(_12727_),
    .Y(_12728_));
 sky130_fd_sc_hd__nand2_1 _20293_ (.A(_11034_),
    .B(_12728_),
    .Y(_12729_));
 sky130_fd_sc_hd__a21boi_0 _20294_ (.A1(_08164_),
    .A2(_10934_),
    .B1_N(\id_stage_i.controller_i.store_err_q ),
    .Y(_12730_));
 sky130_fd_sc_hd__nand2_2 _20295_ (.A(\id_stage_i.controller_i.instr_valid_i ),
    .B(\id_stage_i.controller_i.instr_fetch_err_i ),
    .Y(_12731_));
 sky130_fd_sc_hd__o311ai_1 _20296_ (.A1(\id_stage_i.controller_i.illegal_insn_q ),
    .A2(_12698_),
    .A3(_12730_),
    .B1(_12731_),
    .C1(_12469_),
    .Y(_12732_));
 sky130_fd_sc_hd__nand3_1 _20297_ (.A(net283),
    .B(_12729_),
    .C(_12732_),
    .Y(_12733_));
 sky130_fd_sc_hd__o2111ai_1 _20298_ (.A1(\cs_registers_i.mstack_cause_q[1] ),
    .A2(_12690_),
    .B1(_12717_),
    .C1(_12721_),
    .D1(_12733_),
    .Y(_12734_));
 sky130_fd_sc_hd__o21ai_0 _20299_ (.A1(_12718_),
    .A2(_12717_),
    .B1(_12734_),
    .Y(_00253_));
 sky130_fd_sc_hd__inv_1 _20300_ (.A(\cs_registers_i.mcause_q[2] ),
    .Y(_12735_));
 sky130_fd_sc_hd__nand2_1 _20301_ (.A(_11309_),
    .B(_12688_),
    .Y(_12736_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_592 ();
 sky130_fd_sc_hd__nand3_1 _20303_ (.A(_12731_),
    .B(_12469_),
    .C(_12694_),
    .Y(_12738_));
 sky130_fd_sc_hd__nand2_2 _20304_ (.A(_11013_),
    .B(_11015_),
    .Y(_12739_));
 sky130_fd_sc_hd__nand2_1 _20305_ (.A(_12739_),
    .B(_11024_),
    .Y(_12740_));
 sky130_fd_sc_hd__nand4_2 _20306_ (.A(_11021_),
    .B(_11029_),
    .C(_12727_),
    .D(_12740_),
    .Y(_12741_));
 sky130_fd_sc_hd__nand2_1 _20307_ (.A(_11034_),
    .B(_12741_),
    .Y(_12742_));
 sky130_fd_sc_hd__nand3_1 _20308_ (.A(net283),
    .B(_12738_),
    .C(_12742_),
    .Y(_12743_));
 sky130_fd_sc_hd__o2111ai_1 _20309_ (.A1(\cs_registers_i.mstack_cause_q[2] ),
    .A2(_12690_),
    .B1(_12717_),
    .C1(_12736_),
    .D1(_12743_),
    .Y(_12744_));
 sky130_fd_sc_hd__o21ai_0 _20310_ (.A1(_12735_),
    .A2(_12717_),
    .B1(_12744_),
    .Y(_00254_));
 sky130_fd_sc_hd__nand2_1 _20311_ (.A(_11867_),
    .B(_12688_),
    .Y(_12745_));
 sky130_fd_sc_hd__o2111ai_1 _20312_ (.A1(_11018_),
    .A2(_11027_),
    .B1(_12727_),
    .C1(_11021_),
    .D1(_11024_),
    .Y(_12746_));
 sky130_fd_sc_hd__nand2_1 _20313_ (.A(_11034_),
    .B(_12746_),
    .Y(_12747_));
 sky130_fd_sc_hd__nand4_1 _20314_ (.A(_12695_),
    .B(_10934_),
    .C(_12469_),
    .D(_12696_),
    .Y(_12748_));
 sky130_fd_sc_hd__nand3_1 _20315_ (.A(net281),
    .B(_12747_),
    .C(_12748_),
    .Y(_12749_));
 sky130_fd_sc_hd__o2111ai_1 _20316_ (.A1(\cs_registers_i.mstack_cause_q[3] ),
    .A2(_12690_),
    .B1(_12717_),
    .C1(_12745_),
    .D1(_12749_),
    .Y(_12750_));
 sky130_fd_sc_hd__o21ai_0 _20317_ (.A1(_11852_),
    .A2(_12717_),
    .B1(_12750_),
    .Y(_00255_));
 sky130_fd_sc_hd__inv_1 _20318_ (.A(\cs_registers_i.mcause_q[4] ),
    .Y(_12751_));
 sky130_fd_sc_hd__nand2_1 _20319_ (.A(_11887_),
    .B(_12688_),
    .Y(_12752_));
 sky130_fd_sc_hd__o21ai_4 _20320_ (.A1(_12723_),
    .A2(_12711_),
    .B1(_11034_),
    .Y(_12753_));
 sky130_fd_sc_hd__nand2_1 _20321_ (.A(net277),
    .B(_12753_),
    .Y(_12754_));
 sky130_fd_sc_hd__o2111ai_1 _20322_ (.A1(\cs_registers_i.mstack_cause_q[4] ),
    .A2(_12690_),
    .B1(_12717_),
    .C1(_12752_),
    .D1(_12754_),
    .Y(_12755_));
 sky130_fd_sc_hd__o21ai_0 _20323_ (.A1(_12751_),
    .A2(_12717_),
    .B1(_12755_),
    .Y(_00256_));
 sky130_fd_sc_hd__a221oi_1 _20324_ (.A1(\cs_registers_i.mstack_cause_q[5] ),
    .A2(_12687_),
    .B1(_12688_),
    .B2(_12106_),
    .C1(_11034_),
    .Y(_12756_));
 sky130_fd_sc_hd__nor2_1 _20325_ (.A(\cs_registers_i.mcause_q[5] ),
    .B(_12717_),
    .Y(_12757_));
 sky130_fd_sc_hd__a21oi_1 _20326_ (.A1(_12717_),
    .A2(_12756_),
    .B1(_12757_),
    .Y(_00257_));
 sky130_fd_sc_hd__or2_4 _20327_ (.A(net280),
    .B(_12687_),
    .X(_12758_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_591 ();
 sky130_fd_sc_hd__a21oi_4 _20329_ (.A1(_11243_),
    .A2(_11272_),
    .B1(_12758_),
    .Y(_12760_));
 sky130_fd_sc_hd__a22o_1 _20330_ (.A1(\cs_registers_i.mstack_epc_q[0] ),
    .A2(_12687_),
    .B1(net269),
    .B2(\cs_registers_i.csr_mepc_o[0] ),
    .X(_00258_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_589 ();
 sky130_fd_sc_hd__nand2_1 _20333_ (.A(_12500_),
    .B(net277),
    .Y(_12763_));
 sky130_fd_sc_hd__o221ai_1 _20334_ (.A1(\cs_registers_i.mstack_epc_q[10] ),
    .A2(_12690_),
    .B1(_12758_),
    .B2(_11357_),
    .C1(_12763_),
    .Y(_12764_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_588 ();
 sky130_fd_sc_hd__nand2_1 _20336_ (.A(\cs_registers_i.csr_mepc_o[10] ),
    .B(net269),
    .Y(_12766_));
 sky130_fd_sc_hd__o21ai_0 _20337_ (.A1(net269),
    .A2(_12764_),
    .B1(_12766_),
    .Y(_00259_));
 sky130_fd_sc_hd__nand2_1 _20338_ (.A(_12505_),
    .B(net281),
    .Y(_12767_));
 sky130_fd_sc_hd__o221ai_1 _20339_ (.A1(\cs_registers_i.mstack_epc_q[11] ),
    .A2(_12690_),
    .B1(_12758_),
    .B2(_11391_),
    .C1(_12767_),
    .Y(_12768_));
 sky130_fd_sc_hd__nand2_1 _20340_ (.A(\cs_registers_i.csr_mepc_o[11] ),
    .B(net269),
    .Y(_12769_));
 sky130_fd_sc_hd__o21ai_0 _20341_ (.A1(net269),
    .A2(_12768_),
    .B1(_12769_),
    .Y(_00260_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_587 ();
 sky130_fd_sc_hd__nand2_1 _20343_ (.A(_12509_),
    .B(net281),
    .Y(_12771_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_586 ();
 sky130_fd_sc_hd__nand2_1 _20345_ (.A(_11428_),
    .B(_12688_),
    .Y(_12773_));
 sky130_fd_sc_hd__o211ai_1 _20346_ (.A1(\cs_registers_i.mstack_epc_q[12] ),
    .A2(_12690_),
    .B1(_12771_),
    .C1(_12773_),
    .Y(_12774_));
 sky130_fd_sc_hd__nand2_1 _20347_ (.A(\cs_registers_i.csr_mepc_o[12] ),
    .B(net269),
    .Y(_12775_));
 sky130_fd_sc_hd__o21ai_0 _20348_ (.A1(net269),
    .A2(_12774_),
    .B1(_12775_),
    .Y(_00261_));
 sky130_fd_sc_hd__nand2_1 _20349_ (.A(_12513_),
    .B(net281),
    .Y(_12776_));
 sky130_fd_sc_hd__nand2_1 _20350_ (.A(_11448_),
    .B(_12688_),
    .Y(_12777_));
 sky130_fd_sc_hd__o211ai_1 _20351_ (.A1(\cs_registers_i.mstack_epc_q[13] ),
    .A2(_12690_),
    .B1(_12776_),
    .C1(_12777_),
    .Y(_12778_));
 sky130_fd_sc_hd__nand2_1 _20352_ (.A(\cs_registers_i.csr_mepc_o[13] ),
    .B(net269),
    .Y(_12779_));
 sky130_fd_sc_hd__o21ai_0 _20353_ (.A1(net269),
    .A2(_12778_),
    .B1(_12779_),
    .Y(_00262_));
 sky130_fd_sc_hd__nand2_1 _20354_ (.A(_12516_),
    .B(net281),
    .Y(_12780_));
 sky130_fd_sc_hd__nand2_1 _20355_ (.A(_11465_),
    .B(_12688_),
    .Y(_12781_));
 sky130_fd_sc_hd__o211ai_1 _20356_ (.A1(\cs_registers_i.mstack_epc_q[14] ),
    .A2(_12690_),
    .B1(_12780_),
    .C1(_12781_),
    .Y(_12782_));
 sky130_fd_sc_hd__nand2_1 _20357_ (.A(\cs_registers_i.csr_mepc_o[14] ),
    .B(net269),
    .Y(_12783_));
 sky130_fd_sc_hd__o21ai_0 _20358_ (.A1(net269),
    .A2(_12782_),
    .B1(_12783_),
    .Y(_00263_));
 sky130_fd_sc_hd__nand2_1 _20359_ (.A(_12520_),
    .B(net281),
    .Y(_12784_));
 sky130_fd_sc_hd__nand2_1 _20360_ (.A(_11488_),
    .B(_12688_),
    .Y(_12785_));
 sky130_fd_sc_hd__o211ai_1 _20361_ (.A1(\cs_registers_i.mstack_epc_q[15] ),
    .A2(_12690_),
    .B1(_12784_),
    .C1(_12785_),
    .Y(_12786_));
 sky130_fd_sc_hd__nand2_1 _20362_ (.A(\cs_registers_i.csr_mepc_o[15] ),
    .B(net269),
    .Y(_12787_));
 sky130_fd_sc_hd__o21ai_0 _20363_ (.A1(net269),
    .A2(_12786_),
    .B1(_12787_),
    .Y(_00264_));
 sky130_fd_sc_hd__nand2_1 _20364_ (.A(_12523_),
    .B(net278),
    .Y(_12788_));
 sky130_fd_sc_hd__nand2_1 _20365_ (.A(_11505_),
    .B(_12688_),
    .Y(_12789_));
 sky130_fd_sc_hd__o211ai_1 _20366_ (.A1(\cs_registers_i.mstack_epc_q[16] ),
    .A2(_12690_),
    .B1(_12788_),
    .C1(_12789_),
    .Y(_12790_));
 sky130_fd_sc_hd__nand2_1 _20367_ (.A(\cs_registers_i.csr_mepc_o[16] ),
    .B(net270),
    .Y(_12791_));
 sky130_fd_sc_hd__o21ai_0 _20368_ (.A1(net270),
    .A2(_12790_),
    .B1(_12791_),
    .Y(_00265_));
 sky130_fd_sc_hd__nand2_1 _20369_ (.A(_12526_),
    .B(net278),
    .Y(_12792_));
 sky130_fd_sc_hd__nand2_1 _20370_ (.A(_11523_),
    .B(_12688_),
    .Y(_12793_));
 sky130_fd_sc_hd__o211ai_1 _20371_ (.A1(\cs_registers_i.mstack_epc_q[17] ),
    .A2(_12690_),
    .B1(_12792_),
    .C1(_12793_),
    .Y(_12794_));
 sky130_fd_sc_hd__nand2_1 _20372_ (.A(\cs_registers_i.csr_mepc_o[17] ),
    .B(net270),
    .Y(_12795_));
 sky130_fd_sc_hd__o21ai_0 _20373_ (.A1(net270),
    .A2(_12794_),
    .B1(_12795_),
    .Y(_00266_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_585 ();
 sky130_fd_sc_hd__nand2_1 _20375_ (.A(_12529_),
    .B(net280),
    .Y(_12797_));
 sky130_fd_sc_hd__nand2_1 _20376_ (.A(_11546_),
    .B(_12688_),
    .Y(_12798_));
 sky130_fd_sc_hd__o211ai_1 _20377_ (.A1(\cs_registers_i.mstack_epc_q[18] ),
    .A2(_12690_),
    .B1(_12797_),
    .C1(_12798_),
    .Y(_12799_));
 sky130_fd_sc_hd__nand2_1 _20378_ (.A(\cs_registers_i.csr_mepc_o[18] ),
    .B(_12760_),
    .Y(_12800_));
 sky130_fd_sc_hd__o21ai_0 _20379_ (.A1(_12760_),
    .A2(_12799_),
    .B1(_12800_),
    .Y(_00267_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_584 ();
 sky130_fd_sc_hd__nand2_1 _20381_ (.A(_12532_),
    .B(net278),
    .Y(_12802_));
 sky130_fd_sc_hd__nand2_1 _20382_ (.A(_11563_),
    .B(_12688_),
    .Y(_12803_));
 sky130_fd_sc_hd__o211ai_1 _20383_ (.A1(\cs_registers_i.mstack_epc_q[19] ),
    .A2(_12690_),
    .B1(_12802_),
    .C1(_12803_),
    .Y(_12804_));
 sky130_fd_sc_hd__nand2_1 _20384_ (.A(\cs_registers_i.csr_mepc_o[19] ),
    .B(net270),
    .Y(_12805_));
 sky130_fd_sc_hd__o21ai_0 _20385_ (.A1(net270),
    .A2(_12804_),
    .B1(_12805_),
    .Y(_00268_));
 sky130_fd_sc_hd__nand2_1 _20386_ (.A(_12538_),
    .B(net283),
    .Y(_12806_));
 sky130_fd_sc_hd__o211ai_1 _20387_ (.A1(\cs_registers_i.mstack_epc_q[1] ),
    .A2(_12690_),
    .B1(_12721_),
    .C1(_12806_),
    .Y(_12807_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_583 ();
 sky130_fd_sc_hd__nand2_1 _20389_ (.A(\cs_registers_i.csr_mepc_o[1] ),
    .B(net269),
    .Y(_12809_));
 sky130_fd_sc_hd__o21ai_0 _20390_ (.A1(net269),
    .A2(_12807_),
    .B1(_12809_),
    .Y(_00269_));
 sky130_fd_sc_hd__nand2_1 _20391_ (.A(_12543_),
    .B(net280),
    .Y(_12810_));
 sky130_fd_sc_hd__nand2_1 _20392_ (.A(_11599_),
    .B(_12688_),
    .Y(_12811_));
 sky130_fd_sc_hd__o211ai_1 _20393_ (.A1(\cs_registers_i.mstack_epc_q[20] ),
    .A2(_12690_),
    .B1(_12810_),
    .C1(_12811_),
    .Y(_12812_));
 sky130_fd_sc_hd__nand2_1 _20394_ (.A(\cs_registers_i.csr_mepc_o[20] ),
    .B(_12760_),
    .Y(_12813_));
 sky130_fd_sc_hd__o21ai_0 _20395_ (.A1(_12760_),
    .A2(_12812_),
    .B1(_12813_),
    .Y(_00270_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_582 ();
 sky130_fd_sc_hd__nand2_1 _20397_ (.A(_12546_),
    .B(net279),
    .Y(_12815_));
 sky130_fd_sc_hd__nand2_1 _20398_ (.A(_11623_),
    .B(_12688_),
    .Y(_12816_));
 sky130_fd_sc_hd__o211ai_1 _20399_ (.A1(\cs_registers_i.mstack_epc_q[21] ),
    .A2(_12690_),
    .B1(_12815_),
    .C1(_12816_),
    .Y(_12817_));
 sky130_fd_sc_hd__nand2_1 _20400_ (.A(\cs_registers_i.csr_mepc_o[21] ),
    .B(_12760_),
    .Y(_12818_));
 sky130_fd_sc_hd__o21ai_0 _20401_ (.A1(_12760_),
    .A2(_12817_),
    .B1(_12818_),
    .Y(_00271_));
 sky130_fd_sc_hd__nand2_1 _20402_ (.A(_12549_),
    .B(net280),
    .Y(_12819_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_581 ();
 sky130_fd_sc_hd__nand2_1 _20404_ (.A(_11643_),
    .B(_12688_),
    .Y(_12821_));
 sky130_fd_sc_hd__o211ai_1 _20405_ (.A1(\cs_registers_i.mstack_epc_q[22] ),
    .A2(_12690_),
    .B1(_12819_),
    .C1(_12821_),
    .Y(_12822_));
 sky130_fd_sc_hd__nand2_1 _20406_ (.A(\cs_registers_i.csr_mepc_o[22] ),
    .B(_12760_),
    .Y(_12823_));
 sky130_fd_sc_hd__o21ai_0 _20407_ (.A1(_12760_),
    .A2(_12822_),
    .B1(_12823_),
    .Y(_00272_));
 sky130_fd_sc_hd__nand2_1 _20408_ (.A(_12553_),
    .B(net280),
    .Y(_12824_));
 sky130_fd_sc_hd__nand2_1 _20409_ (.A(_11664_),
    .B(_12688_),
    .Y(_12825_));
 sky130_fd_sc_hd__o211ai_1 _20410_ (.A1(\cs_registers_i.mstack_epc_q[23] ),
    .A2(_12690_),
    .B1(_12824_),
    .C1(_12825_),
    .Y(_12826_));
 sky130_fd_sc_hd__nand2_1 _20411_ (.A(\cs_registers_i.csr_mepc_o[23] ),
    .B(_12760_),
    .Y(_12827_));
 sky130_fd_sc_hd__o21ai_0 _20412_ (.A1(_12760_),
    .A2(_12826_),
    .B1(_12827_),
    .Y(_00273_));
 sky130_fd_sc_hd__nand2_1 _20413_ (.A(_12557_),
    .B(net278),
    .Y(_12828_));
 sky130_fd_sc_hd__nand2_1 _20414_ (.A(_11684_),
    .B(_12688_),
    .Y(_12829_));
 sky130_fd_sc_hd__o211ai_1 _20415_ (.A1(\cs_registers_i.mstack_epc_q[24] ),
    .A2(_12690_),
    .B1(_12828_),
    .C1(_12829_),
    .Y(_12830_));
 sky130_fd_sc_hd__nand2_1 _20416_ (.A(\cs_registers_i.csr_mepc_o[24] ),
    .B(net270),
    .Y(_12831_));
 sky130_fd_sc_hd__o21ai_0 _20417_ (.A1(net270),
    .A2(_12830_),
    .B1(_12831_),
    .Y(_00274_));
 sky130_fd_sc_hd__nand2_1 _20418_ (.A(_12560_),
    .B(net279),
    .Y(_12832_));
 sky130_fd_sc_hd__nand2_1 _20419_ (.A(_11706_),
    .B(_12688_),
    .Y(_12833_));
 sky130_fd_sc_hd__o211ai_1 _20420_ (.A1(\cs_registers_i.mstack_epc_q[25] ),
    .A2(_12690_),
    .B1(_12832_),
    .C1(_12833_),
    .Y(_12834_));
 sky130_fd_sc_hd__nand2_1 _20421_ (.A(\cs_registers_i.csr_mepc_o[25] ),
    .B(_12760_),
    .Y(_12835_));
 sky130_fd_sc_hd__o21ai_0 _20422_ (.A1(_12760_),
    .A2(_12834_),
    .B1(_12835_),
    .Y(_00275_));
 sky130_fd_sc_hd__nand2_1 _20423_ (.A(_12563_),
    .B(net278),
    .Y(_12836_));
 sky130_fd_sc_hd__nand2_1 _20424_ (.A(_11726_),
    .B(_12688_),
    .Y(_12837_));
 sky130_fd_sc_hd__o211ai_1 _20425_ (.A1(\cs_registers_i.mstack_epc_q[26] ),
    .A2(_12690_),
    .B1(_12836_),
    .C1(_12837_),
    .Y(_12838_));
 sky130_fd_sc_hd__nand2_1 _20426_ (.A(\cs_registers_i.csr_mepc_o[26] ),
    .B(net270),
    .Y(_12839_));
 sky130_fd_sc_hd__o21ai_0 _20427_ (.A1(net270),
    .A2(_12838_),
    .B1(_12839_),
    .Y(_00276_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_580 ();
 sky130_fd_sc_hd__nand2_1 _20429_ (.A(_12566_),
    .B(net278),
    .Y(_12841_));
 sky130_fd_sc_hd__nand2_1 _20430_ (.A(_11746_),
    .B(_12688_),
    .Y(_12842_));
 sky130_fd_sc_hd__o211ai_1 _20431_ (.A1(\cs_registers_i.mstack_epc_q[27] ),
    .A2(_12690_),
    .B1(_12841_),
    .C1(_12842_),
    .Y(_12843_));
 sky130_fd_sc_hd__nand2_1 _20432_ (.A(\cs_registers_i.csr_mepc_o[27] ),
    .B(net270),
    .Y(_12844_));
 sky130_fd_sc_hd__o21ai_0 _20433_ (.A1(net270),
    .A2(_12843_),
    .B1(_12844_),
    .Y(_00277_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_579 ();
 sky130_fd_sc_hd__nand2_1 _20435_ (.A(_12569_),
    .B(net278),
    .Y(_12846_));
 sky130_fd_sc_hd__nand2_1 _20436_ (.A(_11765_),
    .B(_12688_),
    .Y(_12847_));
 sky130_fd_sc_hd__o211ai_1 _20437_ (.A1(\cs_registers_i.mstack_epc_q[28] ),
    .A2(_12690_),
    .B1(_12846_),
    .C1(_12847_),
    .Y(_12848_));
 sky130_fd_sc_hd__nand2_1 _20438_ (.A(\cs_registers_i.csr_mepc_o[28] ),
    .B(net270),
    .Y(_12849_));
 sky130_fd_sc_hd__o21ai_0 _20439_ (.A1(net270),
    .A2(_12848_),
    .B1(_12849_),
    .Y(_00278_));
 sky130_fd_sc_hd__nand2_1 _20440_ (.A(_12573_),
    .B(net278),
    .Y(_12850_));
 sky130_fd_sc_hd__nand2_1 _20441_ (.A(_11785_),
    .B(_12688_),
    .Y(_12851_));
 sky130_fd_sc_hd__o211ai_1 _20442_ (.A1(\cs_registers_i.mstack_epc_q[29] ),
    .A2(_12690_),
    .B1(_12850_),
    .C1(_12851_),
    .Y(_12852_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_578 ();
 sky130_fd_sc_hd__nand2_1 _20444_ (.A(\cs_registers_i.csr_mepc_o[29] ),
    .B(net270),
    .Y(_12854_));
 sky130_fd_sc_hd__o21ai_0 _20445_ (.A1(net270),
    .A2(_12852_),
    .B1(_12854_),
    .Y(_00279_));
 sky130_fd_sc_hd__nand2_1 _20446_ (.A(_12578_),
    .B(net283),
    .Y(_12855_));
 sky130_fd_sc_hd__o211ai_1 _20447_ (.A1(\cs_registers_i.mstack_epc_q[2] ),
    .A2(_12690_),
    .B1(_12736_),
    .C1(_12855_),
    .Y(_12856_));
 sky130_fd_sc_hd__nand2_1 _20448_ (.A(\cs_registers_i.csr_mepc_o[2] ),
    .B(net269),
    .Y(_12857_));
 sky130_fd_sc_hd__o21ai_0 _20449_ (.A1(net269),
    .A2(_12856_),
    .B1(_12857_),
    .Y(_00280_));
 sky130_fd_sc_hd__nand2_1 _20450_ (.A(_12581_),
    .B(net279),
    .Y(_12858_));
 sky130_fd_sc_hd__nand2_1 _20451_ (.A(_11808_),
    .B(_12688_),
    .Y(_12859_));
 sky130_fd_sc_hd__o211ai_1 _20452_ (.A1(\cs_registers_i.mstack_epc_q[30] ),
    .A2(_12690_),
    .B1(_12858_),
    .C1(_12859_),
    .Y(_12860_));
 sky130_fd_sc_hd__nand2_1 _20453_ (.A(\cs_registers_i.csr_mepc_o[30] ),
    .B(net270),
    .Y(_12861_));
 sky130_fd_sc_hd__o21ai_0 _20454_ (.A1(net270),
    .A2(_12860_),
    .B1(_12861_),
    .Y(_00281_));
 sky130_fd_sc_hd__nand2_1 _20455_ (.A(_12584_),
    .B(net280),
    .Y(_12862_));
 sky130_fd_sc_hd__o221ai_1 _20456_ (.A1(\cs_registers_i.mstack_epc_q[31] ),
    .A2(_12690_),
    .B1(_12758_),
    .B2(_12106_),
    .C1(_12862_),
    .Y(_12863_));
 sky130_fd_sc_hd__nand2_1 _20457_ (.A(\cs_registers_i.csr_mepc_o[31] ),
    .B(net270),
    .Y(_12864_));
 sky130_fd_sc_hd__o21ai_0 _20458_ (.A1(net270),
    .A2(_12863_),
    .B1(_12864_),
    .Y(_00282_));
 sky130_fd_sc_hd__nand2_1 _20459_ (.A(_12587_),
    .B(net281),
    .Y(_12865_));
 sky130_fd_sc_hd__o211ai_1 _20460_ (.A1(\cs_registers_i.mstack_epc_q[3] ),
    .A2(_12690_),
    .B1(_12745_),
    .C1(_12865_),
    .Y(_12866_));
 sky130_fd_sc_hd__nand2_1 _20461_ (.A(\cs_registers_i.csr_mepc_o[3] ),
    .B(net269),
    .Y(_12867_));
 sky130_fd_sc_hd__o21ai_0 _20462_ (.A1(net269),
    .A2(_12866_),
    .B1(_12867_),
    .Y(_00283_));
 sky130_fd_sc_hd__nand2_1 _20463_ (.A(_12590_),
    .B(net277),
    .Y(_12868_));
 sky130_fd_sc_hd__o211ai_1 _20464_ (.A1(\cs_registers_i.mstack_epc_q[4] ),
    .A2(_12690_),
    .B1(_12752_),
    .C1(_12868_),
    .Y(_12869_));
 sky130_fd_sc_hd__nand2_1 _20465_ (.A(\cs_registers_i.csr_mepc_o[4] ),
    .B(net269),
    .Y(_12870_));
 sky130_fd_sc_hd__o21ai_0 _20466_ (.A1(net269),
    .A2(_12869_),
    .B1(_12870_),
    .Y(_00284_));
 sky130_fd_sc_hd__nand2_1 _20467_ (.A(_12593_),
    .B(net277),
    .Y(_12871_));
 sky130_fd_sc_hd__o221ai_1 _20468_ (.A1(\cs_registers_i.mstack_epc_q[5] ),
    .A2(_12690_),
    .B1(_12758_),
    .B2(_11902_),
    .C1(_12871_),
    .Y(_12872_));
 sky130_fd_sc_hd__nand2_1 _20469_ (.A(\cs_registers_i.csr_mepc_o[5] ),
    .B(net269),
    .Y(_12873_));
 sky130_fd_sc_hd__o21ai_0 _20470_ (.A1(net269),
    .A2(_12872_),
    .B1(_12873_),
    .Y(_00285_));
 sky130_fd_sc_hd__nand2_1 _20471_ (.A(_12597_),
    .B(net277),
    .Y(_12874_));
 sky130_fd_sc_hd__o221ai_1 _20472_ (.A1(\cs_registers_i.mstack_epc_q[6] ),
    .A2(_12690_),
    .B1(_12758_),
    .B2(_11917_),
    .C1(_12874_),
    .Y(_12875_));
 sky130_fd_sc_hd__nand2_1 _20473_ (.A(\cs_registers_i.csr_mepc_o[6] ),
    .B(net269),
    .Y(_12876_));
 sky130_fd_sc_hd__o21ai_0 _20474_ (.A1(net269),
    .A2(_12875_),
    .B1(_12876_),
    .Y(_00286_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_577 ();
 sky130_fd_sc_hd__nand2_1 _20476_ (.A(_12600_),
    .B(net277),
    .Y(_12878_));
 sky130_fd_sc_hd__nand2_1 _20477_ (.A(_11935_),
    .B(_12688_),
    .Y(_12879_));
 sky130_fd_sc_hd__o211ai_1 _20478_ (.A1(\cs_registers_i.mstack_epc_q[7] ),
    .A2(_12690_),
    .B1(_12878_),
    .C1(_12879_),
    .Y(_12880_));
 sky130_fd_sc_hd__nand2_1 _20479_ (.A(\cs_registers_i.csr_mepc_o[7] ),
    .B(net269),
    .Y(_12881_));
 sky130_fd_sc_hd__o21ai_0 _20480_ (.A1(net269),
    .A2(_12880_),
    .B1(_12881_),
    .Y(_00287_));
 sky130_fd_sc_hd__nand2_1 _20481_ (.A(_12603_),
    .B(net277),
    .Y(_12882_));
 sky130_fd_sc_hd__nand2_1 _20482_ (.A(_11957_),
    .B(_12688_),
    .Y(_12883_));
 sky130_fd_sc_hd__o211ai_1 _20483_ (.A1(\cs_registers_i.mstack_epc_q[8] ),
    .A2(_12690_),
    .B1(_12882_),
    .C1(_12883_),
    .Y(_12884_));
 sky130_fd_sc_hd__nand2_1 _20484_ (.A(\cs_registers_i.csr_mepc_o[8] ),
    .B(net269),
    .Y(_12885_));
 sky130_fd_sc_hd__o21ai_0 _20485_ (.A1(net269),
    .A2(_12884_),
    .B1(_12885_),
    .Y(_00288_));
 sky130_fd_sc_hd__nand2_1 _20486_ (.A(_12606_),
    .B(net277),
    .Y(_12886_));
 sky130_fd_sc_hd__nand2_1 _20487_ (.A(_11973_),
    .B(_12688_),
    .Y(_12887_));
 sky130_fd_sc_hd__o211ai_1 _20488_ (.A1(\cs_registers_i.mstack_epc_q[9] ),
    .A2(_12690_),
    .B1(_12886_),
    .C1(_12887_),
    .Y(_12888_));
 sky130_fd_sc_hd__nand2_1 _20489_ (.A(\cs_registers_i.csr_mepc_o[9] ),
    .B(net269),
    .Y(_12889_));
 sky130_fd_sc_hd__o21ai_0 _20490_ (.A1(net269),
    .A2(_12888_),
    .B1(_12889_),
    .Y(_00289_));
 sky130_fd_sc_hd__nand2_8 _20491_ (.A(net271),
    .B(_11373_),
    .Y(_12890_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_575 ();
 sky130_fd_sc_hd__nand2_1 _20494_ (.A(\cs_registers_i.mie_q[0] ),
    .B(_12890_),
    .Y(_12893_));
 sky130_fd_sc_hd__o21ai_0 _20495_ (.A1(_11505_),
    .A2(_12890_),
    .B1(_12893_),
    .Y(_00290_));
 sky130_fd_sc_hd__nand2_1 _20496_ (.A(\cs_registers_i.mie_q[10] ),
    .B(_12890_),
    .Y(_12894_));
 sky130_fd_sc_hd__o21ai_0 _20497_ (.A1(_11726_),
    .A2(_12890_),
    .B1(_12894_),
    .Y(_00291_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_574 ();
 sky130_fd_sc_hd__nand2_1 _20499_ (.A(\cs_registers_i.mie_q[11] ),
    .B(_12890_),
    .Y(_12896_));
 sky130_fd_sc_hd__o21ai_0 _20500_ (.A1(_11746_),
    .A2(_12890_),
    .B1(_12896_),
    .Y(_00292_));
 sky130_fd_sc_hd__nand2_1 _20501_ (.A(\cs_registers_i.mie_q[12] ),
    .B(_12890_),
    .Y(_12897_));
 sky130_fd_sc_hd__o21ai_0 _20502_ (.A1(_11765_),
    .A2(_12890_),
    .B1(_12897_),
    .Y(_00293_));
 sky130_fd_sc_hd__nand2_1 _20503_ (.A(\cs_registers_i.mie_q[13] ),
    .B(_12890_),
    .Y(_12898_));
 sky130_fd_sc_hd__o21ai_0 _20504_ (.A1(_11785_),
    .A2(_12890_),
    .B1(_12898_),
    .Y(_00294_));
 sky130_fd_sc_hd__nand2_1 _20505_ (.A(\cs_registers_i.mie_q[14] ),
    .B(_12890_),
    .Y(_12899_));
 sky130_fd_sc_hd__o21ai_0 _20506_ (.A1(_11808_),
    .A2(_12890_),
    .B1(_12899_),
    .Y(_00295_));
 sky130_fd_sc_hd__nand2_1 _20507_ (.A(\cs_registers_i.mie_q[15] ),
    .B(_12890_),
    .Y(_12900_));
 sky130_fd_sc_hd__o21ai_0 _20508_ (.A1(_12481_),
    .A2(_12890_),
    .B1(_12900_),
    .Y(_00296_));
 sky130_fd_sc_hd__nand2_1 _20509_ (.A(\cs_registers_i.mie_q[16] ),
    .B(_12890_),
    .Y(_12901_));
 sky130_fd_sc_hd__o21ai_0 _20510_ (.A1(_11935_),
    .A2(_12890_),
    .B1(_12901_),
    .Y(_00297_));
 sky130_fd_sc_hd__nand2_1 _20511_ (.A(\cs_registers_i.mie_q[17] ),
    .B(_12890_),
    .Y(_12902_));
 sky130_fd_sc_hd__o21ai_0 _20512_ (.A1(_11867_),
    .A2(_12890_),
    .B1(_12902_),
    .Y(_00298_));
 sky130_fd_sc_hd__nand2_1 _20513_ (.A(\cs_registers_i.mie_q[1] ),
    .B(_12890_),
    .Y(_12903_));
 sky130_fd_sc_hd__o21ai_0 _20514_ (.A1(_11523_),
    .A2(_12890_),
    .B1(_12903_),
    .Y(_00299_));
 sky130_fd_sc_hd__nand2_1 _20515_ (.A(\cs_registers_i.mie_q[2] ),
    .B(_12890_),
    .Y(_12904_));
 sky130_fd_sc_hd__o21ai_0 _20516_ (.A1(_11546_),
    .A2(_12890_),
    .B1(_12904_),
    .Y(_00300_));
 sky130_fd_sc_hd__nand2_1 _20517_ (.A(\cs_registers_i.mie_q[3] ),
    .B(_12890_),
    .Y(_12905_));
 sky130_fd_sc_hd__o21ai_0 _20518_ (.A1(_11563_),
    .A2(_12890_),
    .B1(_12905_),
    .Y(_00301_));
 sky130_fd_sc_hd__nand2_1 _20519_ (.A(\cs_registers_i.mie_q[4] ),
    .B(_12890_),
    .Y(_12906_));
 sky130_fd_sc_hd__o21ai_0 _20520_ (.A1(_11599_),
    .A2(_12890_),
    .B1(_12906_),
    .Y(_00302_));
 sky130_fd_sc_hd__nand2_1 _20521_ (.A(\cs_registers_i.mie_q[5] ),
    .B(_12890_),
    .Y(_12907_));
 sky130_fd_sc_hd__o21ai_0 _20522_ (.A1(_11623_),
    .A2(_12890_),
    .B1(_12907_),
    .Y(_00303_));
 sky130_fd_sc_hd__nand2_1 _20523_ (.A(\cs_registers_i.mie_q[6] ),
    .B(_12890_),
    .Y(_12908_));
 sky130_fd_sc_hd__o21ai_0 _20524_ (.A1(_11643_),
    .A2(_12890_),
    .B1(_12908_),
    .Y(_00304_));
 sky130_fd_sc_hd__nand2_1 _20525_ (.A(\cs_registers_i.mie_q[7] ),
    .B(_12890_),
    .Y(_12909_));
 sky130_fd_sc_hd__o21ai_0 _20526_ (.A1(_11664_),
    .A2(_12890_),
    .B1(_12909_),
    .Y(_00305_));
 sky130_fd_sc_hd__nand2_1 _20527_ (.A(\cs_registers_i.mie_q[8] ),
    .B(_12890_),
    .Y(_12910_));
 sky130_fd_sc_hd__o21ai_0 _20528_ (.A1(_11684_),
    .A2(_12890_),
    .B1(_12910_),
    .Y(_00306_));
 sky130_fd_sc_hd__nand2_1 _20529_ (.A(\cs_registers_i.mie_q[9] ),
    .B(_12890_),
    .Y(_12911_));
 sky130_fd_sc_hd__o21ai_0 _20530_ (.A1(_11706_),
    .A2(_12890_),
    .B1(_12911_),
    .Y(_00307_));
 sky130_fd_sc_hd__nand2_8 _20531_ (.A(net271),
    .B(_11255_),
    .Y(_12912_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_572 ();
 sky130_fd_sc_hd__nand2_1 _20534_ (.A(\cs_registers_i.mscratch_q[0] ),
    .B(_12912_),
    .Y(_12915_));
 sky130_fd_sc_hd__o21ai_0 _20535_ (.A1(_11280_),
    .A2(_12912_),
    .B1(_12915_),
    .Y(_00308_));
 sky130_fd_sc_hd__mux2_1 _20536_ (.A0(_11357_),
    .A1(\cs_registers_i.mscratch_q[10] ),
    .S(_12912_),
    .X(_00309_));
 sky130_fd_sc_hd__nand2_1 _20537_ (.A(\cs_registers_i.mscratch_q[11] ),
    .B(_12912_),
    .Y(_12916_));
 sky130_fd_sc_hd__o21ai_0 _20538_ (.A1(_12481_),
    .A2(_12912_),
    .B1(_12916_),
    .Y(_00310_));
 sky130_fd_sc_hd__nand2_1 _20539_ (.A(\cs_registers_i.mscratch_q[12] ),
    .B(_12912_),
    .Y(_12917_));
 sky130_fd_sc_hd__o21ai_0 _20540_ (.A1(_11428_),
    .A2(_12912_),
    .B1(_12917_),
    .Y(_00311_));
 sky130_fd_sc_hd__nand2_1 _20541_ (.A(\cs_registers_i.mscratch_q[13] ),
    .B(_12912_),
    .Y(_12918_));
 sky130_fd_sc_hd__o21ai_0 _20542_ (.A1(_11448_),
    .A2(_12912_),
    .B1(_12918_),
    .Y(_00312_));
 sky130_fd_sc_hd__nand2_1 _20543_ (.A(\cs_registers_i.mscratch_q[14] ),
    .B(_12912_),
    .Y(_12919_));
 sky130_fd_sc_hd__o21ai_0 _20544_ (.A1(_11465_),
    .A2(_12912_),
    .B1(_12919_),
    .Y(_00313_));
 sky130_fd_sc_hd__nand2_1 _20545_ (.A(\cs_registers_i.mscratch_q[15] ),
    .B(_12912_),
    .Y(_12920_));
 sky130_fd_sc_hd__o21ai_0 _20546_ (.A1(_11488_),
    .A2(_12912_),
    .B1(_12920_),
    .Y(_00314_));
 sky130_fd_sc_hd__nand2_1 _20547_ (.A(\cs_registers_i.mscratch_q[16] ),
    .B(_12912_),
    .Y(_12921_));
 sky130_fd_sc_hd__o21ai_0 _20548_ (.A1(_11505_),
    .A2(_12912_),
    .B1(_12921_),
    .Y(_00315_));
 sky130_fd_sc_hd__nand2_1 _20549_ (.A(\cs_registers_i.mscratch_q[17] ),
    .B(_12912_),
    .Y(_12922_));
 sky130_fd_sc_hd__o21ai_0 _20550_ (.A1(_11523_),
    .A2(_12912_),
    .B1(_12922_),
    .Y(_00316_));
 sky130_fd_sc_hd__nand2_1 _20551_ (.A(\cs_registers_i.mscratch_q[18] ),
    .B(_12912_),
    .Y(_12923_));
 sky130_fd_sc_hd__o21ai_0 _20552_ (.A1(_11546_),
    .A2(_12912_),
    .B1(_12923_),
    .Y(_00317_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_571 ();
 sky130_fd_sc_hd__nand2_1 _20554_ (.A(\cs_registers_i.mscratch_q[19] ),
    .B(_12912_),
    .Y(_12925_));
 sky130_fd_sc_hd__o21ai_0 _20555_ (.A1(_11563_),
    .A2(_12912_),
    .B1(_12925_),
    .Y(_00318_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_570 ();
 sky130_fd_sc_hd__nand2_1 _20557_ (.A(\cs_registers_i.mscratch_q[1] ),
    .B(_12912_),
    .Y(_12927_));
 sky130_fd_sc_hd__o21ai_0 _20558_ (.A1(_11582_),
    .A2(_12912_),
    .B1(_12927_),
    .Y(_00319_));
 sky130_fd_sc_hd__nand2_1 _20559_ (.A(\cs_registers_i.mscratch_q[20] ),
    .B(_12912_),
    .Y(_12928_));
 sky130_fd_sc_hd__o21ai_0 _20560_ (.A1(_11599_),
    .A2(_12912_),
    .B1(_12928_),
    .Y(_00320_));
 sky130_fd_sc_hd__nand2_1 _20561_ (.A(\cs_registers_i.mscratch_q[21] ),
    .B(_12912_),
    .Y(_12929_));
 sky130_fd_sc_hd__o21ai_0 _20562_ (.A1(_11623_),
    .A2(_12912_),
    .B1(_12929_),
    .Y(_00321_));
 sky130_fd_sc_hd__nand2_1 _20563_ (.A(\cs_registers_i.mscratch_q[22] ),
    .B(_12912_),
    .Y(_12930_));
 sky130_fd_sc_hd__o21ai_0 _20564_ (.A1(_11643_),
    .A2(_12912_),
    .B1(_12930_),
    .Y(_00322_));
 sky130_fd_sc_hd__nand2_1 _20565_ (.A(\cs_registers_i.mscratch_q[23] ),
    .B(_12912_),
    .Y(_12931_));
 sky130_fd_sc_hd__o21ai_0 _20566_ (.A1(_11664_),
    .A2(_12912_),
    .B1(_12931_),
    .Y(_00323_));
 sky130_fd_sc_hd__nand2_1 _20567_ (.A(\cs_registers_i.mscratch_q[24] ),
    .B(_12912_),
    .Y(_12932_));
 sky130_fd_sc_hd__o21ai_0 _20568_ (.A1(_11684_),
    .A2(_12912_),
    .B1(_12932_),
    .Y(_00324_));
 sky130_fd_sc_hd__nand2_1 _20569_ (.A(\cs_registers_i.mscratch_q[25] ),
    .B(_12912_),
    .Y(_12933_));
 sky130_fd_sc_hd__o21ai_0 _20570_ (.A1(_11706_),
    .A2(_12912_),
    .B1(_12933_),
    .Y(_00325_));
 sky130_fd_sc_hd__nand2_1 _20571_ (.A(\cs_registers_i.mscratch_q[26] ),
    .B(_12912_),
    .Y(_12934_));
 sky130_fd_sc_hd__o21ai_0 _20572_ (.A1(_11726_),
    .A2(_12912_),
    .B1(_12934_),
    .Y(_00326_));
 sky130_fd_sc_hd__nand2_1 _20573_ (.A(\cs_registers_i.mscratch_q[27] ),
    .B(_12912_),
    .Y(_12935_));
 sky130_fd_sc_hd__o21ai_0 _20574_ (.A1(_11746_),
    .A2(_12912_),
    .B1(_12935_),
    .Y(_00327_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_569 ();
 sky130_fd_sc_hd__nand2_1 _20576_ (.A(\cs_registers_i.mscratch_q[28] ),
    .B(_12912_),
    .Y(_12937_));
 sky130_fd_sc_hd__o21ai_0 _20577_ (.A1(_11765_),
    .A2(_12912_),
    .B1(_12937_),
    .Y(_00328_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_568 ();
 sky130_fd_sc_hd__nand2_1 _20579_ (.A(\cs_registers_i.mscratch_q[29] ),
    .B(_12912_),
    .Y(_12939_));
 sky130_fd_sc_hd__o21ai_0 _20580_ (.A1(_11785_),
    .A2(_12912_),
    .B1(_12939_),
    .Y(_00329_));
 sky130_fd_sc_hd__nand2_1 _20581_ (.A(\cs_registers_i.mscratch_q[2] ),
    .B(_12912_),
    .Y(_12940_));
 sky130_fd_sc_hd__o21ai_0 _20582_ (.A1(_11309_),
    .A2(_12912_),
    .B1(_12940_),
    .Y(_00330_));
 sky130_fd_sc_hd__nand2_1 _20583_ (.A(\cs_registers_i.mscratch_q[30] ),
    .B(_12912_),
    .Y(_12941_));
 sky130_fd_sc_hd__o21ai_0 _20584_ (.A1(_11808_),
    .A2(_12912_),
    .B1(_12941_),
    .Y(_00331_));
 sky130_fd_sc_hd__nand2_1 _20585_ (.A(\cs_registers_i.mscratch_q[31] ),
    .B(_12912_),
    .Y(_12942_));
 sky130_fd_sc_hd__o21ai_0 _20586_ (.A1(_11826_),
    .A2(_12912_),
    .B1(_12942_),
    .Y(_00332_));
 sky130_fd_sc_hd__nand2_1 _20587_ (.A(\cs_registers_i.mscratch_q[3] ),
    .B(_12912_),
    .Y(_12943_));
 sky130_fd_sc_hd__o21ai_0 _20588_ (.A1(_11867_),
    .A2(_12912_),
    .B1(_12943_),
    .Y(_00333_));
 sky130_fd_sc_hd__nand2_1 _20589_ (.A(\cs_registers_i.mscratch_q[4] ),
    .B(_12912_),
    .Y(_12944_));
 sky130_fd_sc_hd__o21ai_0 _20590_ (.A1(_11887_),
    .A2(_12912_),
    .B1(_12944_),
    .Y(_00334_));
 sky130_fd_sc_hd__nand2_1 _20591_ (.A(\cs_registers_i.mscratch_q[5] ),
    .B(_12912_),
    .Y(_12945_));
 sky130_fd_sc_hd__o21ai_0 _20592_ (.A1(_12594_),
    .A2(_12912_),
    .B1(_12945_),
    .Y(_00335_));
 sky130_fd_sc_hd__nand2_1 _20593_ (.A(\cs_registers_i.mscratch_q[6] ),
    .B(_12912_),
    .Y(_12946_));
 sky130_fd_sc_hd__o21ai_0 _20594_ (.A1(_12113_),
    .A2(_12912_),
    .B1(_12946_),
    .Y(_00336_));
 sky130_fd_sc_hd__nand2_1 _20595_ (.A(\cs_registers_i.mscratch_q[7] ),
    .B(_12912_),
    .Y(_12947_));
 sky130_fd_sc_hd__o21ai_0 _20596_ (.A1(_11935_),
    .A2(_12912_),
    .B1(_12947_),
    .Y(_00337_));
 sky130_fd_sc_hd__nand2_1 _20597_ (.A(\cs_registers_i.mscratch_q[8] ),
    .B(_12912_),
    .Y(_12948_));
 sky130_fd_sc_hd__o21ai_0 _20598_ (.A1(_11957_),
    .A2(_12912_),
    .B1(_12948_),
    .Y(_00338_));
 sky130_fd_sc_hd__nand2_1 _20599_ (.A(\cs_registers_i.mscratch_q[9] ),
    .B(_12912_),
    .Y(_12949_));
 sky130_fd_sc_hd__o21ai_0 _20600_ (.A1(_11973_),
    .A2(_12912_),
    .B1(_12949_),
    .Y(_00339_));
 sky130_fd_sc_hd__mux2_1 _20601_ (.A0(\cs_registers_i.mstack_cause_q[0] ),
    .A1(\cs_registers_i.mcause_q[0] ),
    .S(net283),
    .X(_00340_));
 sky130_fd_sc_hd__mux2_1 _20602_ (.A0(\cs_registers_i.mstack_cause_q[1] ),
    .A1(\cs_registers_i.mcause_q[1] ),
    .S(net283),
    .X(_00341_));
 sky130_fd_sc_hd__mux2_1 _20603_ (.A0(\cs_registers_i.mstack_cause_q[2] ),
    .A1(\cs_registers_i.mcause_q[2] ),
    .S(net283),
    .X(_00342_));
 sky130_fd_sc_hd__mux2_1 _20604_ (.A0(\cs_registers_i.mstack_cause_q[3] ),
    .A1(\cs_registers_i.mcause_q[3] ),
    .S(net282),
    .X(_00343_));
 sky130_fd_sc_hd__mux2_1 _20605_ (.A0(\cs_registers_i.mstack_cause_q[4] ),
    .A1(\cs_registers_i.mcause_q[4] ),
    .S(net277),
    .X(_00344_));
 sky130_fd_sc_hd__mux2_1 _20606_ (.A0(\cs_registers_i.mstack_cause_q[5] ),
    .A1(\cs_registers_i.mcause_q[5] ),
    .S(net280),
    .X(_00345_));
 sky130_fd_sc_hd__mux2_1 _20607_ (.A0(\cs_registers_i.mstack_q[0] ),
    .A1(\cs_registers_i.mstack_d[0] ),
    .S(net282),
    .X(_00346_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_567 ();
 sky130_fd_sc_hd__mux2_1 _20609_ (.A0(\cs_registers_i.mstack_q[1] ),
    .A1(\cs_registers_i.mstack_d[1] ),
    .S(net280),
    .X(_00347_));
 sky130_fd_sc_hd__mux2_1 _20610_ (.A0(\cs_registers_i.mstack_q[2] ),
    .A1(\cs_registers_i.mstack_d[2] ),
    .S(net281),
    .X(_00348_));
 sky130_fd_sc_hd__mux2_1 _20611_ (.A0(\cs_registers_i.mstack_epc_q[0] ),
    .A1(\cs_registers_i.csr_mepc_o[0] ),
    .S(net282),
    .X(_00349_));
 sky130_fd_sc_hd__mux2_1 _20612_ (.A0(\cs_registers_i.mstack_epc_q[10] ),
    .A1(\cs_registers_i.csr_mepc_o[10] ),
    .S(net277),
    .X(_00350_));
 sky130_fd_sc_hd__mux2_1 _20613_ (.A0(\cs_registers_i.mstack_epc_q[11] ),
    .A1(\cs_registers_i.csr_mepc_o[11] ),
    .S(net281),
    .X(_00351_));
 sky130_fd_sc_hd__mux2_1 _20614_ (.A0(\cs_registers_i.mstack_epc_q[12] ),
    .A1(\cs_registers_i.csr_mepc_o[12] ),
    .S(net281),
    .X(_00352_));
 sky130_fd_sc_hd__mux2_1 _20615_ (.A0(\cs_registers_i.mstack_epc_q[13] ),
    .A1(\cs_registers_i.csr_mepc_o[13] ),
    .S(net281),
    .X(_00353_));
 sky130_fd_sc_hd__mux2_1 _20616_ (.A0(\cs_registers_i.mstack_epc_q[14] ),
    .A1(\cs_registers_i.csr_mepc_o[14] ),
    .S(net281),
    .X(_00354_));
 sky130_fd_sc_hd__mux2_1 _20617_ (.A0(\cs_registers_i.mstack_epc_q[15] ),
    .A1(\cs_registers_i.csr_mepc_o[15] ),
    .S(net281),
    .X(_00355_));
 sky130_fd_sc_hd__mux2_1 _20618_ (.A0(\cs_registers_i.mstack_epc_q[16] ),
    .A1(\cs_registers_i.csr_mepc_o[16] ),
    .S(net278),
    .X(_00356_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_566 ();
 sky130_fd_sc_hd__mux2_1 _20620_ (.A0(\cs_registers_i.mstack_epc_q[17] ),
    .A1(\cs_registers_i.csr_mepc_o[17] ),
    .S(net278),
    .X(_00357_));
 sky130_fd_sc_hd__mux2_1 _20621_ (.A0(\cs_registers_i.mstack_epc_q[18] ),
    .A1(\cs_registers_i.csr_mepc_o[18] ),
    .S(net280),
    .X(_00358_));
 sky130_fd_sc_hd__mux2_1 _20622_ (.A0(\cs_registers_i.mstack_epc_q[19] ),
    .A1(\cs_registers_i.csr_mepc_o[19] ),
    .S(net278),
    .X(_00359_));
 sky130_fd_sc_hd__mux2_1 _20623_ (.A0(\cs_registers_i.mstack_epc_q[1] ),
    .A1(\cs_registers_i.csr_mepc_o[1] ),
    .S(net283),
    .X(_00360_));
 sky130_fd_sc_hd__mux2_1 _20624_ (.A0(\cs_registers_i.mstack_epc_q[20] ),
    .A1(\cs_registers_i.csr_mepc_o[20] ),
    .S(net280),
    .X(_00361_));
 sky130_fd_sc_hd__mux2_1 _20625_ (.A0(\cs_registers_i.mstack_epc_q[21] ),
    .A1(\cs_registers_i.csr_mepc_o[21] ),
    .S(net279),
    .X(_00362_));
 sky130_fd_sc_hd__mux2_1 _20626_ (.A0(\cs_registers_i.mstack_epc_q[22] ),
    .A1(\cs_registers_i.csr_mepc_o[22] ),
    .S(net280),
    .X(_00363_));
 sky130_fd_sc_hd__mux2_1 _20627_ (.A0(\cs_registers_i.mstack_epc_q[23] ),
    .A1(\cs_registers_i.csr_mepc_o[23] ),
    .S(net280),
    .X(_00364_));
 sky130_fd_sc_hd__mux2_1 _20628_ (.A0(\cs_registers_i.mstack_epc_q[24] ),
    .A1(\cs_registers_i.csr_mepc_o[24] ),
    .S(net278),
    .X(_00365_));
 sky130_fd_sc_hd__mux2_1 _20629_ (.A0(\cs_registers_i.mstack_epc_q[25] ),
    .A1(\cs_registers_i.csr_mepc_o[25] ),
    .S(net279),
    .X(_00366_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_565 ();
 sky130_fd_sc_hd__mux2_1 _20631_ (.A0(\cs_registers_i.mstack_epc_q[26] ),
    .A1(\cs_registers_i.csr_mepc_o[26] ),
    .S(net278),
    .X(_00367_));
 sky130_fd_sc_hd__mux2_1 _20632_ (.A0(\cs_registers_i.mstack_epc_q[27] ),
    .A1(\cs_registers_i.csr_mepc_o[27] ),
    .S(net278),
    .X(_00368_));
 sky130_fd_sc_hd__mux2_1 _20633_ (.A0(\cs_registers_i.mstack_epc_q[28] ),
    .A1(\cs_registers_i.csr_mepc_o[28] ),
    .S(net278),
    .X(_00369_));
 sky130_fd_sc_hd__mux2_1 _20634_ (.A0(\cs_registers_i.mstack_epc_q[29] ),
    .A1(\cs_registers_i.csr_mepc_o[29] ),
    .S(net278),
    .X(_00370_));
 sky130_fd_sc_hd__mux2_1 _20635_ (.A0(\cs_registers_i.mstack_epc_q[2] ),
    .A1(\cs_registers_i.csr_mepc_o[2] ),
    .S(net283),
    .X(_00371_));
 sky130_fd_sc_hd__mux2_1 _20636_ (.A0(\cs_registers_i.mstack_epc_q[30] ),
    .A1(\cs_registers_i.csr_mepc_o[30] ),
    .S(net279),
    .X(_00372_));
 sky130_fd_sc_hd__mux2_1 _20637_ (.A0(\cs_registers_i.mstack_epc_q[31] ),
    .A1(\cs_registers_i.csr_mepc_o[31] ),
    .S(net280),
    .X(_00373_));
 sky130_fd_sc_hd__mux2_1 _20638_ (.A0(\cs_registers_i.mstack_epc_q[3] ),
    .A1(\cs_registers_i.csr_mepc_o[3] ),
    .S(net281),
    .X(_00374_));
 sky130_fd_sc_hd__mux2_1 _20639_ (.A0(\cs_registers_i.mstack_epc_q[4] ),
    .A1(\cs_registers_i.csr_mepc_o[4] ),
    .S(net277),
    .X(_00375_));
 sky130_fd_sc_hd__mux2_1 _20640_ (.A0(\cs_registers_i.mstack_epc_q[5] ),
    .A1(\cs_registers_i.csr_mepc_o[5] ),
    .S(net277),
    .X(_00376_));
 sky130_fd_sc_hd__mux2_1 _20641_ (.A0(\cs_registers_i.mstack_epc_q[6] ),
    .A1(\cs_registers_i.csr_mepc_o[6] ),
    .S(net277),
    .X(_00377_));
 sky130_fd_sc_hd__mux2_1 _20642_ (.A0(\cs_registers_i.mstack_epc_q[7] ),
    .A1(\cs_registers_i.csr_mepc_o[7] ),
    .S(net277),
    .X(_00378_));
 sky130_fd_sc_hd__mux2_1 _20643_ (.A0(\cs_registers_i.mstack_epc_q[8] ),
    .A1(\cs_registers_i.csr_mepc_o[8] ),
    .S(net277),
    .X(_00379_));
 sky130_fd_sc_hd__mux2_1 _20644_ (.A0(\cs_registers_i.mstack_epc_q[9] ),
    .A1(\cs_registers_i.csr_mepc_o[9] ),
    .S(net277),
    .X(_00380_));
 sky130_fd_sc_hd__nand2_4 _20645_ (.A(_11243_),
    .B(_11375_),
    .Y(_12953_));
 sky130_fd_sc_hd__nand2_1 _20646_ (.A(\cs_registers_i.csr_mstatus_tw_o ),
    .B(_12953_),
    .Y(_12954_));
 sky130_fd_sc_hd__o21ai_0 _20647_ (.A1(_11623_),
    .A2(_12953_),
    .B1(_12954_),
    .Y(_00381_));
 sky130_fd_sc_hd__nand2_1 _20648_ (.A(\cs_registers_i.mstatus_q[1] ),
    .B(_12953_),
    .Y(_12955_));
 sky130_fd_sc_hd__o21ai_0 _20649_ (.A1(_11523_),
    .A2(_12953_),
    .B1(_12955_),
    .Y(_00382_));
 sky130_fd_sc_hd__and2_0 _20650_ (.A(_12481_),
    .B(_11428_),
    .X(_12956_));
 sky130_fd_sc_hd__a22oi_1 _20651_ (.A1(\cs_registers_i.priv_lvl_q[0] ),
    .A2(net282),
    .B1(_12687_),
    .B2(\cs_registers_i.mstack_q[0] ),
    .Y(_12957_));
 sky130_fd_sc_hd__o21ai_0 _20652_ (.A1(_12953_),
    .A2(_12956_),
    .B1(_12957_),
    .Y(_12958_));
 sky130_fd_sc_hd__nand4_1 _20653_ (.A(net1137),
    .B(net1146),
    .C(_10858_),
    .D(_10875_),
    .Y(_12959_));
 sky130_fd_sc_hd__nor3_1 _20654_ (.A(_10896_),
    .B(_10886_),
    .C(_12959_),
    .Y(_12960_));
 sky130_fd_sc_hd__a211oi_2 _20655_ (.A1(_10931_),
    .A2(_12960_),
    .B1(net280),
    .C1(_12455_),
    .Y(_12961_));
 sky130_fd_sc_hd__mux2_1 _20656_ (.A0(_12958_),
    .A1(\cs_registers_i.mstack_d[0] ),
    .S(_12961_),
    .X(_00383_));
 sky130_fd_sc_hd__a22oi_1 _20657_ (.A1(\cs_registers_i.priv_lvl_q[1] ),
    .A2(net280),
    .B1(_12687_),
    .B2(\cs_registers_i.mstack_q[1] ),
    .Y(_12962_));
 sky130_fd_sc_hd__o21ai_0 _20658_ (.A1(_12953_),
    .A2(_12956_),
    .B1(_12962_),
    .Y(_12963_));
 sky130_fd_sc_hd__mux2_1 _20659_ (.A0(_12963_),
    .A1(\cs_registers_i.mstack_d[1] ),
    .S(_12961_),
    .X(_00384_));
 sky130_fd_sc_hd__nand2_1 _20660_ (.A(\cs_registers_i.csr_mstatus_mie_o ),
    .B(net281),
    .Y(_12964_));
 sky130_fd_sc_hd__o21ai_0 _20661_ (.A1(_11032_),
    .A2(\cs_registers_i.mstack_q[2] ),
    .B1(_12455_),
    .Y(_12965_));
 sky130_fd_sc_hd__nor2_1 _20662_ (.A(_11935_),
    .B(_12953_),
    .Y(_12966_));
 sky130_fd_sc_hd__a21oi_1 _20663_ (.A1(\cs_registers_i.mstack_d[2] ),
    .A2(_12953_),
    .B1(_12966_),
    .Y(_12967_));
 sky130_fd_sc_hd__or3_1 _20664_ (.A(_12455_),
    .B(net281),
    .C(_12967_),
    .X(_12968_));
 sky130_fd_sc_hd__nand3_1 _20665_ (.A(_12964_),
    .B(_12965_),
    .C(_12968_),
    .Y(_00385_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_564 ();
 sky130_fd_sc_hd__nor2_1 _20667_ (.A(_11867_),
    .B(_12953_),
    .Y(_12970_));
 sky130_fd_sc_hd__a21oi_1 _20668_ (.A1(\cs_registers_i.csr_mstatus_mie_o ),
    .A2(_12953_),
    .B1(_12970_),
    .Y(_12971_));
 sky130_fd_sc_hd__nor2_1 _20669_ (.A(_12452_),
    .B(_12971_),
    .Y(_12972_));
 sky130_fd_sc_hd__a21oi_1 _20670_ (.A1(\cs_registers_i.mstack_d[2] ),
    .A2(_12452_),
    .B1(_12972_),
    .Y(_12973_));
 sky130_fd_sc_hd__nor2_1 _20671_ (.A(net281),
    .B(_12973_),
    .Y(_00386_));
 sky130_fd_sc_hd__nand2_8 _20672_ (.A(_11243_),
    .B(_11270_),
    .Y(_12974_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_563 ();
 sky130_fd_sc_hd__nor2_1 _20674_ (.A(_11280_),
    .B(_12974_),
    .Y(_12976_));
 sky130_fd_sc_hd__a21oi_1 _20675_ (.A1(\cs_registers_i.mtval_q[0] ),
    .A2(_12974_),
    .B1(_12976_),
    .Y(_12977_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_562 ();
 sky130_fd_sc_hd__mux2_1 _20677_ (.A0(\id_stage_i.controller_i.instr_i[0] ),
    .A1(\id_stage_i.controller_i.instr_compressed_i[0] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .X(_12979_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_561 ();
 sky130_fd_sc_hd__a22o_1 _20679_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[0] ),
    .A2(net298),
    .B1(_12979_),
    .B2(\id_stage_i.controller_i.illegal_insn_q ),
    .X(_12981_));
 sky130_fd_sc_hd__nand4_1 _20680_ (.A(_12731_),
    .B(_12469_),
    .C(_12685_),
    .D(_12981_),
    .Y(_12982_));
 sky130_fd_sc_hd__o21ai_0 _20681_ (.A1(_12685_),
    .A2(_12977_),
    .B1(_12982_),
    .Y(_00387_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_560 ();
 sky130_fd_sc_hd__inv_1 _20683_ (.A(\cs_registers_i.pc_id_i[3] ),
    .Y(_12984_));
 sky130_fd_sc_hd__nand3_1 _20684_ (.A(\cs_registers_i.pc_id_i[1] ),
    .B(\cs_registers_i.pc_id_i[2] ),
    .C(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .Y(_12985_));
 sky130_fd_sc_hd__nor2_1 _20685_ (.A(_12984_),
    .B(_12985_),
    .Y(_12986_));
 sky130_fd_sc_hd__and3_1 _20686_ (.A(\cs_registers_i.pc_id_i[4] ),
    .B(\cs_registers_i.pc_id_i[5] ),
    .C(_12986_),
    .X(_12987_));
 sky130_fd_sc_hd__nand3_1 _20687_ (.A(\cs_registers_i.pc_id_i[6] ),
    .B(\cs_registers_i.pc_id_i[7] ),
    .C(_12987_),
    .Y(_12988_));
 sky130_fd_sc_hd__nor2_1 _20688_ (.A(_09185_),
    .B(_12988_),
    .Y(_12989_));
 sky130_fd_sc_hd__nand2_1 _20689_ (.A(\cs_registers_i.pc_id_i[9] ),
    .B(_12989_),
    .Y(_12990_));
 sky130_fd_sc_hd__xnor2_1 _20690_ (.A(\cs_registers_i.pc_id_i[10] ),
    .B(_12990_),
    .Y(_12991_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_558 ();
 sky130_fd_sc_hd__mux2_1 _20693_ (.A0(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .A1(\id_stage_i.controller_i.instr_compressed_i[10] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .X(_12994_));
 sky130_fd_sc_hd__a22oi_1 _20694_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[10] ),
    .A2(_12694_),
    .B1(_12994_),
    .B2(\id_stage_i.controller_i.illegal_insn_q ),
    .Y(_12995_));
 sky130_fd_sc_hd__nor2_1 _20695_ (.A(_11040_),
    .B(_12995_),
    .Y(_12996_));
 sky130_fd_sc_hd__a21oi_1 _20696_ (.A1(_11040_),
    .A2(_12991_),
    .B1(_12996_),
    .Y(_12997_));
 sky130_fd_sc_hd__nand2_8 _20697_ (.A(_12469_),
    .B(_12685_),
    .Y(_12998_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_557 ();
 sky130_fd_sc_hd__mux2i_1 _20699_ (.A0(_11357_),
    .A1(\cs_registers_i.mtval_q[10] ),
    .S(_12974_),
    .Y(_13000_));
 sky130_fd_sc_hd__o22ai_1 _20700_ (.A1(_12997_),
    .A2(_12998_),
    .B1(_13000_),
    .B2(net283),
    .Y(_00388_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_556 ();
 sky130_fd_sc_hd__nand3_1 _20702_ (.A(\cs_registers_i.pc_id_i[9] ),
    .B(\cs_registers_i.pc_id_i[10] ),
    .C(_12989_),
    .Y(_13002_));
 sky130_fd_sc_hd__xnor2_1 _20703_ (.A(\cs_registers_i.pc_id_i[11] ),
    .B(_13002_),
    .Y(_13003_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_553 ();
 sky130_fd_sc_hd__mux2_1 _20707_ (.A0(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .A1(\id_stage_i.controller_i.instr_compressed_i[11] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .X(_13007_));
 sky130_fd_sc_hd__a22oi_1 _20708_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[11] ),
    .A2(net298),
    .B1(_13007_),
    .B2(\id_stage_i.controller_i.illegal_insn_q ),
    .Y(_13008_));
 sky130_fd_sc_hd__nor2_1 _20709_ (.A(_11040_),
    .B(_13008_),
    .Y(_13009_));
 sky130_fd_sc_hd__a21oi_2 _20710_ (.A1(_11040_),
    .A2(_13003_),
    .B1(_13009_),
    .Y(_13010_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_552 ();
 sky130_fd_sc_hd__nor2_1 _20712_ (.A(_12481_),
    .B(_12974_),
    .Y(_13012_));
 sky130_fd_sc_hd__a21oi_1 _20713_ (.A1(\cs_registers_i.mtval_q[11] ),
    .A2(_12974_),
    .B1(_13012_),
    .Y(_13013_));
 sky130_fd_sc_hd__o22ai_1 _20714_ (.A1(_12998_),
    .A2(_13010_),
    .B1(_13013_),
    .B2(net281),
    .Y(_00389_));
 sky130_fd_sc_hd__nand4_1 _20715_ (.A(\cs_registers_i.pc_id_i[11] ),
    .B(\cs_registers_i.pc_id_i[9] ),
    .C(\cs_registers_i.pc_id_i[10] ),
    .D(_12989_),
    .Y(_13014_));
 sky130_fd_sc_hd__xnor2_1 _20716_ (.A(\cs_registers_i.pc_id_i[12] ),
    .B(_13014_),
    .Y(_13015_));
 sky130_fd_sc_hd__nand2_1 _20717_ (.A(\id_stage_i.controller_i.instr_is_compressed_i ),
    .B(\id_stage_i.controller_i.instr_compressed_i[12] ),
    .Y(_13016_));
 sky130_fd_sc_hd__o21ai_0 _20718_ (.A1(_08254_),
    .A2(\id_stage_i.controller_i.instr_is_compressed_i ),
    .B1(_13016_),
    .Y(_13017_));
 sky130_fd_sc_hd__a22oi_1 _20719_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[12] ),
    .A2(net298),
    .B1(_13017_),
    .B2(\id_stage_i.controller_i.illegal_insn_q ),
    .Y(_13018_));
 sky130_fd_sc_hd__nor2_1 _20720_ (.A(_11040_),
    .B(_13018_),
    .Y(_13019_));
 sky130_fd_sc_hd__a21oi_1 _20721_ (.A1(_11040_),
    .A2(_13015_),
    .B1(_13019_),
    .Y(_13020_));
 sky130_fd_sc_hd__nor2_1 _20722_ (.A(_11428_),
    .B(_12974_),
    .Y(_13021_));
 sky130_fd_sc_hd__a21oi_1 _20723_ (.A1(\cs_registers_i.mtval_q[12] ),
    .A2(_12974_),
    .B1(_13021_),
    .Y(_13022_));
 sky130_fd_sc_hd__o22ai_1 _20724_ (.A1(_12998_),
    .A2(_13020_),
    .B1(_13022_),
    .B2(_12685_),
    .Y(_00390_));
 sky130_fd_sc_hd__inv_1 _20725_ (.A(\cs_registers_i.pc_id_i[12] ),
    .Y(_13023_));
 sky130_fd_sc_hd__nor2_1 _20726_ (.A(_13023_),
    .B(_13014_),
    .Y(_13024_));
 sky130_fd_sc_hd__xor2_1 _20727_ (.A(\cs_registers_i.pc_id_i[13] ),
    .B(_13024_),
    .X(_13025_));
 sky130_fd_sc_hd__mux2_1 _20728_ (.A0(net676),
    .A1(\id_stage_i.controller_i.instr_compressed_i[13] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .X(_13026_));
 sky130_fd_sc_hd__a22oi_1 _20729_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[13] ),
    .A2(net298),
    .B1(_13026_),
    .B2(\id_stage_i.controller_i.illegal_insn_q ),
    .Y(_13027_));
 sky130_fd_sc_hd__nor2_1 _20730_ (.A(_11040_),
    .B(_13027_),
    .Y(_13028_));
 sky130_fd_sc_hd__a21oi_1 _20731_ (.A1(_11040_),
    .A2(_13025_),
    .B1(_13028_),
    .Y(_13029_));
 sky130_fd_sc_hd__nor2_1 _20732_ (.A(_11448_),
    .B(_12974_),
    .Y(_13030_));
 sky130_fd_sc_hd__a21oi_1 _20733_ (.A1(\cs_registers_i.mtval_q[13] ),
    .A2(_12974_),
    .B1(_13030_),
    .Y(_13031_));
 sky130_fd_sc_hd__o22ai_1 _20734_ (.A1(_12998_),
    .A2(_13029_),
    .B1(_13031_),
    .B2(_12685_),
    .Y(_00391_));
 sky130_fd_sc_hd__and2_1 _20735_ (.A(\cs_registers_i.pc_id_i[13] ),
    .B(_13024_),
    .X(_13032_));
 sky130_fd_sc_hd__xor2_1 _20736_ (.A(\cs_registers_i.pc_id_i[14] ),
    .B(_13032_),
    .X(_13033_));
 sky130_fd_sc_hd__nand2_1 _20737_ (.A(\id_stage_i.controller_i.instr_is_compressed_i ),
    .B(\id_stage_i.controller_i.instr_compressed_i[14] ),
    .Y(_13034_));
 sky130_fd_sc_hd__o21ai_0 _20738_ (.A1(_08100_),
    .A2(\id_stage_i.controller_i.instr_is_compressed_i ),
    .B1(_13034_),
    .Y(_13035_));
 sky130_fd_sc_hd__a22oi_1 _20739_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[14] ),
    .A2(net298),
    .B1(_13035_),
    .B2(\id_stage_i.controller_i.illegal_insn_q ),
    .Y(_13036_));
 sky130_fd_sc_hd__nor2_1 _20740_ (.A(_11040_),
    .B(_13036_),
    .Y(_13037_));
 sky130_fd_sc_hd__a21oi_1 _20741_ (.A1(_11040_),
    .A2(_13033_),
    .B1(_13037_),
    .Y(_13038_));
 sky130_fd_sc_hd__nor2_1 _20742_ (.A(_11465_),
    .B(_12974_),
    .Y(_13039_));
 sky130_fd_sc_hd__a21oi_1 _20743_ (.A1(\cs_registers_i.mtval_q[14] ),
    .A2(_12974_),
    .B1(_13039_),
    .Y(_13040_));
 sky130_fd_sc_hd__o22ai_1 _20744_ (.A1(_12998_),
    .A2(_13038_),
    .B1(_13040_),
    .B2(_12685_),
    .Y(_00392_));
 sky130_fd_sc_hd__nand2_1 _20745_ (.A(\cs_registers_i.pc_id_i[14] ),
    .B(_13032_),
    .Y(_13041_));
 sky130_fd_sc_hd__xnor2_1 _20746_ (.A(\cs_registers_i.pc_id_i[15] ),
    .B(_13041_),
    .Y(_13042_));
 sky130_fd_sc_hd__mux2_2 _20747_ (.A0(net571),
    .A1(\id_stage_i.controller_i.instr_compressed_i[15] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .X(_13043_));
 sky130_fd_sc_hd__a22oi_1 _20748_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[15] ),
    .A2(net298),
    .B1(_13043_),
    .B2(\id_stage_i.controller_i.illegal_insn_q ),
    .Y(_13044_));
 sky130_fd_sc_hd__nor2_1 _20749_ (.A(_11040_),
    .B(_13044_),
    .Y(_13045_));
 sky130_fd_sc_hd__a21oi_1 _20750_ (.A1(_11040_),
    .A2(_13042_),
    .B1(_13045_),
    .Y(_13046_));
 sky130_fd_sc_hd__nor2_1 _20751_ (.A(_11488_),
    .B(_12974_),
    .Y(_13047_));
 sky130_fd_sc_hd__a21oi_1 _20752_ (.A1(\cs_registers_i.mtval_q[15] ),
    .A2(_12974_),
    .B1(_13047_),
    .Y(_13048_));
 sky130_fd_sc_hd__o22ai_1 _20753_ (.A1(_12998_),
    .A2(_13046_),
    .B1(_13048_),
    .B2(_12685_),
    .Y(_00393_));
 sky130_fd_sc_hd__nand3_4 _20754_ (.A(\cs_registers_i.pc_id_i[14] ),
    .B(\cs_registers_i.pc_id_i[15] ),
    .C(_13032_),
    .Y(_13049_));
 sky130_fd_sc_hd__xnor2_1 _20755_ (.A(\cs_registers_i.pc_id_i[16] ),
    .B(_13049_),
    .Y(_13050_));
 sky130_fd_sc_hd__nor2b_4 _20756_ (.A(\id_stage_i.controller_i.instr_is_compressed_i ),
    .B_N(\id_stage_i.controller_i.illegal_insn_q ),
    .Y(_13051_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_550 ();
 sky130_fd_sc_hd__a22oi_1 _20759_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[16] ),
    .A2(net298),
    .B1(_13051_),
    .B2(net627),
    .Y(_13054_));
 sky130_fd_sc_hd__nor2_1 _20760_ (.A(_11040_),
    .B(_13054_),
    .Y(_13055_));
 sky130_fd_sc_hd__a21oi_1 _20761_ (.A1(_11040_),
    .A2(_13050_),
    .B1(_13055_),
    .Y(_13056_));
 sky130_fd_sc_hd__nor2_1 _20762_ (.A(_11505_),
    .B(_12974_),
    .Y(_13057_));
 sky130_fd_sc_hd__a21oi_1 _20763_ (.A1(\cs_registers_i.mtval_q[16] ),
    .A2(_12974_),
    .B1(_13057_),
    .Y(_13058_));
 sky130_fd_sc_hd__o22ai_1 _20764_ (.A1(_12998_),
    .A2(_13056_),
    .B1(_13058_),
    .B2(net278),
    .Y(_00394_));
 sky130_fd_sc_hd__inv_1 _20765_ (.A(\cs_registers_i.pc_id_i[16] ),
    .Y(_13059_));
 sky130_fd_sc_hd__nor2_1 _20766_ (.A(_13059_),
    .B(_13049_),
    .Y(_13060_));
 sky130_fd_sc_hd__xor2_1 _20767_ (.A(\cs_registers_i.pc_id_i[17] ),
    .B(_13060_),
    .X(_13061_));
 sky130_fd_sc_hd__a22oi_1 _20768_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[17] ),
    .A2(net298),
    .B1(_13051_),
    .B2(net662),
    .Y(_13062_));
 sky130_fd_sc_hd__nor2_1 _20769_ (.A(_11040_),
    .B(_13062_),
    .Y(_13063_));
 sky130_fd_sc_hd__a21oi_1 _20770_ (.A1(_11040_),
    .A2(_13061_),
    .B1(_13063_),
    .Y(_13064_));
 sky130_fd_sc_hd__nor2_1 _20771_ (.A(_11523_),
    .B(_12974_),
    .Y(_13065_));
 sky130_fd_sc_hd__a21oi_1 _20772_ (.A1(\cs_registers_i.mtval_q[17] ),
    .A2(_12974_),
    .B1(_13065_),
    .Y(_13066_));
 sky130_fd_sc_hd__o22ai_1 _20773_ (.A1(_12998_),
    .A2(_13064_),
    .B1(_13066_),
    .B2(net278),
    .Y(_00395_));
 sky130_fd_sc_hd__nand2_1 _20774_ (.A(\cs_registers_i.pc_id_i[17] ),
    .B(_13060_),
    .Y(_13067_));
 sky130_fd_sc_hd__xnor2_1 _20775_ (.A(\cs_registers_i.pc_id_i[18] ),
    .B(_13067_),
    .Y(_13068_));
 sky130_fd_sc_hd__a22oi_1 _20776_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[18] ),
    .A2(net298),
    .B1(_13051_),
    .B2(net588),
    .Y(_13069_));
 sky130_fd_sc_hd__nor2_1 _20777_ (.A(_11040_),
    .B(_13069_),
    .Y(_13070_));
 sky130_fd_sc_hd__a21oi_1 _20778_ (.A1(_11040_),
    .A2(_13068_),
    .B1(_13070_),
    .Y(_13071_));
 sky130_fd_sc_hd__nor2_1 _20779_ (.A(_11546_),
    .B(_12974_),
    .Y(_13072_));
 sky130_fd_sc_hd__a21oi_1 _20780_ (.A1(\cs_registers_i.mtval_q[18] ),
    .A2(_12974_),
    .B1(_13072_),
    .Y(_13073_));
 sky130_fd_sc_hd__o22ai_1 _20781_ (.A1(_12998_),
    .A2(_13071_),
    .B1(_13073_),
    .B2(net278),
    .Y(_00396_));
 sky130_fd_sc_hd__nand3_1 _20782_ (.A(\cs_registers_i.pc_id_i[17] ),
    .B(\cs_registers_i.pc_id_i[18] ),
    .C(_13060_),
    .Y(_13074_));
 sky130_fd_sc_hd__xnor2_1 _20783_ (.A(\cs_registers_i.pc_id_i[19] ),
    .B(_13074_),
    .Y(_13075_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_549 ();
 sky130_fd_sc_hd__a22oi_1 _20785_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[19] ),
    .A2(net298),
    .B1(_13051_),
    .B2(net385),
    .Y(_13077_));
 sky130_fd_sc_hd__nor2_1 _20786_ (.A(_11040_),
    .B(_13077_),
    .Y(_13078_));
 sky130_fd_sc_hd__a21oi_1 _20787_ (.A1(_11040_),
    .A2(_13075_),
    .B1(_13078_),
    .Y(_13079_));
 sky130_fd_sc_hd__nor2_1 _20788_ (.A(_11563_),
    .B(_12974_),
    .Y(_13080_));
 sky130_fd_sc_hd__a21oi_1 _20789_ (.A1(\cs_registers_i.mtval_q[19] ),
    .A2(_12974_),
    .B1(_13080_),
    .Y(_13081_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_548 ();
 sky130_fd_sc_hd__o22ai_1 _20791_ (.A1(_12998_),
    .A2(_13079_),
    .B1(_13081_),
    .B2(net278),
    .Y(_00397_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_547 ();
 sky130_fd_sc_hd__xor2_1 _20793_ (.A(\cs_registers_i.pc_id_i[1] ),
    .B(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .X(_13084_));
 sky130_fd_sc_hd__mux2_1 _20794_ (.A0(\id_stage_i.controller_i.instr_i[1] ),
    .A1(\id_stage_i.controller_i.instr_compressed_i[1] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .X(_13085_));
 sky130_fd_sc_hd__a22oi_1 _20795_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[1] ),
    .A2(_12694_),
    .B1(_13085_),
    .B2(\id_stage_i.controller_i.illegal_insn_q ),
    .Y(_13086_));
 sky130_fd_sc_hd__nor2_1 _20796_ (.A(_11040_),
    .B(_13086_),
    .Y(_13087_));
 sky130_fd_sc_hd__a21oi_1 _20797_ (.A1(_11040_),
    .A2(_13084_),
    .B1(_13087_),
    .Y(_13088_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_546 ();
 sky130_fd_sc_hd__nor2_1 _20799_ (.A(_11582_),
    .B(_12974_),
    .Y(_13090_));
 sky130_fd_sc_hd__a21oi_1 _20800_ (.A1(\cs_registers_i.mtval_q[1] ),
    .A2(_12974_),
    .B1(_13090_),
    .Y(_13091_));
 sky130_fd_sc_hd__o22ai_1 _20801_ (.A1(_12998_),
    .A2(_13088_),
    .B1(_13091_),
    .B2(net283),
    .Y(_00398_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_545 ();
 sky130_fd_sc_hd__inv_1 _20803_ (.A(\cs_registers_i.pc_id_i[19] ),
    .Y(_13093_));
 sky130_fd_sc_hd__nor2_1 _20804_ (.A(_13093_),
    .B(_13074_),
    .Y(_13094_));
 sky130_fd_sc_hd__xor2_1 _20805_ (.A(\cs_registers_i.pc_id_i[20] ),
    .B(_13094_),
    .X(_13095_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_544 ();
 sky130_fd_sc_hd__a22oi_1 _20807_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[20] ),
    .A2(net298),
    .B1(_13051_),
    .B2(net382),
    .Y(_13097_));
 sky130_fd_sc_hd__nor2_1 _20808_ (.A(_11040_),
    .B(_13097_),
    .Y(_13098_));
 sky130_fd_sc_hd__a21oi_1 _20809_ (.A1(_11040_),
    .A2(_13095_),
    .B1(_13098_),
    .Y(_13099_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_543 ();
 sky130_fd_sc_hd__nor2_1 _20811_ (.A(_11599_),
    .B(_12974_),
    .Y(_13101_));
 sky130_fd_sc_hd__a21oi_1 _20812_ (.A1(\cs_registers_i.mtval_q[20] ),
    .A2(_12974_),
    .B1(_13101_),
    .Y(_13102_));
 sky130_fd_sc_hd__o22ai_1 _20813_ (.A1(_12998_),
    .A2(_13099_),
    .B1(_13102_),
    .B2(net279),
    .Y(_00399_));
 sky130_fd_sc_hd__nand2_1 _20814_ (.A(\cs_registers_i.pc_id_i[20] ),
    .B(_13094_),
    .Y(_13103_));
 sky130_fd_sc_hd__xnor2_1 _20815_ (.A(\cs_registers_i.pc_id_i[21] ),
    .B(_13103_),
    .Y(_13104_));
 sky130_fd_sc_hd__a22oi_1 _20816_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[21] ),
    .A2(net298),
    .B1(_13051_),
    .B2(net372),
    .Y(_13105_));
 sky130_fd_sc_hd__nor2_1 _20817_ (.A(_11040_),
    .B(_13105_),
    .Y(_13106_));
 sky130_fd_sc_hd__a21oi_1 _20818_ (.A1(_11040_),
    .A2(_13104_),
    .B1(_13106_),
    .Y(_13107_));
 sky130_fd_sc_hd__nor2_1 _20819_ (.A(_11623_),
    .B(_12974_),
    .Y(_13108_));
 sky130_fd_sc_hd__a21oi_1 _20820_ (.A1(\cs_registers_i.mtval_q[21] ),
    .A2(_12974_),
    .B1(_13108_),
    .Y(_13109_));
 sky130_fd_sc_hd__o22ai_1 _20821_ (.A1(_12998_),
    .A2(_13107_),
    .B1(_13109_),
    .B2(net279),
    .Y(_00400_));
 sky130_fd_sc_hd__nand3_1 _20822_ (.A(\cs_registers_i.pc_id_i[20] ),
    .B(\cs_registers_i.pc_id_i[21] ),
    .C(_13094_),
    .Y(_13110_));
 sky130_fd_sc_hd__xnor2_1 _20823_ (.A(\cs_registers_i.pc_id_i[22] ),
    .B(_13110_),
    .Y(_13111_));
 sky130_fd_sc_hd__a22oi_1 _20824_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[22] ),
    .A2(net298),
    .B1(_13051_),
    .B2(net555),
    .Y(_13112_));
 sky130_fd_sc_hd__nor2_1 _20825_ (.A(_11040_),
    .B(_13112_),
    .Y(_13113_));
 sky130_fd_sc_hd__a21oi_1 _20826_ (.A1(_11040_),
    .A2(_13111_),
    .B1(_13113_),
    .Y(_13114_));
 sky130_fd_sc_hd__nor2_1 _20827_ (.A(_11643_),
    .B(_12974_),
    .Y(_13115_));
 sky130_fd_sc_hd__a21oi_1 _20828_ (.A1(\cs_registers_i.mtval_q[22] ),
    .A2(_12974_),
    .B1(_13115_),
    .Y(_13116_));
 sky130_fd_sc_hd__o22ai_1 _20829_ (.A1(_12998_),
    .A2(_13114_),
    .B1(_13116_),
    .B2(net279),
    .Y(_00401_));
 sky130_fd_sc_hd__inv_1 _20830_ (.A(\cs_registers_i.pc_id_i[22] ),
    .Y(_13117_));
 sky130_fd_sc_hd__nor2_1 _20831_ (.A(_13117_),
    .B(_13110_),
    .Y(_13118_));
 sky130_fd_sc_hd__xor2_1 _20832_ (.A(\cs_registers_i.pc_id_i[23] ),
    .B(_13118_),
    .X(_13119_));
 sky130_fd_sc_hd__a22oi_1 _20833_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[23] ),
    .A2(net298),
    .B1(_13051_),
    .B2(net547),
    .Y(_13120_));
 sky130_fd_sc_hd__nor2_1 _20834_ (.A(_11040_),
    .B(_13120_),
    .Y(_13121_));
 sky130_fd_sc_hd__a21oi_1 _20835_ (.A1(_11040_),
    .A2(_13119_),
    .B1(_13121_),
    .Y(_13122_));
 sky130_fd_sc_hd__nor2_1 _20836_ (.A(_11664_),
    .B(_12974_),
    .Y(_13123_));
 sky130_fd_sc_hd__a21oi_1 _20837_ (.A1(\cs_registers_i.mtval_q[23] ),
    .A2(_12974_),
    .B1(_13123_),
    .Y(_13124_));
 sky130_fd_sc_hd__o22ai_1 _20838_ (.A1(_12998_),
    .A2(_13122_),
    .B1(_13124_),
    .B2(net279),
    .Y(_00402_));
 sky130_fd_sc_hd__nand2_1 _20839_ (.A(\cs_registers_i.pc_id_i[23] ),
    .B(_13118_),
    .Y(_13125_));
 sky130_fd_sc_hd__xnor2_1 _20840_ (.A(\cs_registers_i.pc_id_i[24] ),
    .B(_13125_),
    .Y(_13126_));
 sky130_fd_sc_hd__a22oi_1 _20841_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[24] ),
    .A2(net298),
    .B1(_13051_),
    .B2(net755),
    .Y(_13127_));
 sky130_fd_sc_hd__nor2_1 _20842_ (.A(_11040_),
    .B(_13127_),
    .Y(_13128_));
 sky130_fd_sc_hd__a21oi_2 _20843_ (.A1(_11040_),
    .A2(_13126_),
    .B1(_13128_),
    .Y(_13129_));
 sky130_fd_sc_hd__nor2_1 _20844_ (.A(_11684_),
    .B(_12974_),
    .Y(_13130_));
 sky130_fd_sc_hd__a21oi_1 _20845_ (.A1(\cs_registers_i.mtval_q[24] ),
    .A2(_12974_),
    .B1(_13130_),
    .Y(_13131_));
 sky130_fd_sc_hd__o22ai_1 _20846_ (.A1(_12998_),
    .A2(_13129_),
    .B1(_13131_),
    .B2(net278),
    .Y(_00403_));
 sky130_fd_sc_hd__nand3_1 _20847_ (.A(\cs_registers_i.pc_id_i[23] ),
    .B(\cs_registers_i.pc_id_i[24] ),
    .C(_13118_),
    .Y(_13132_));
 sky130_fd_sc_hd__xnor2_1 _20848_ (.A(\cs_registers_i.pc_id_i[25] ),
    .B(_13132_),
    .Y(_13133_));
 sky130_fd_sc_hd__a22oi_1 _20849_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[25] ),
    .A2(net298),
    .B1(_13051_),
    .B2(net584),
    .Y(_13134_));
 sky130_fd_sc_hd__nor2_1 _20850_ (.A(_11040_),
    .B(_13134_),
    .Y(_13135_));
 sky130_fd_sc_hd__a21oi_1 _20851_ (.A1(_11040_),
    .A2(_13133_),
    .B1(_13135_),
    .Y(_13136_));
 sky130_fd_sc_hd__nor2_1 _20852_ (.A(_11706_),
    .B(_12974_),
    .Y(_13137_));
 sky130_fd_sc_hd__a21oi_1 _20853_ (.A1(\cs_registers_i.mtval_q[25] ),
    .A2(_12974_),
    .B1(_13137_),
    .Y(_13138_));
 sky130_fd_sc_hd__o22ai_1 _20854_ (.A1(_12998_),
    .A2(_13136_),
    .B1(_13138_),
    .B2(net279),
    .Y(_00404_));
 sky130_fd_sc_hd__inv_1 _20855_ (.A(\cs_registers_i.pc_id_i[25] ),
    .Y(_13139_));
 sky130_fd_sc_hd__nor2_1 _20856_ (.A(_13139_),
    .B(_13132_),
    .Y(_13140_));
 sky130_fd_sc_hd__xor2_1 _20857_ (.A(\cs_registers_i.pc_id_i[26] ),
    .B(_13140_),
    .X(_13141_));
 sky130_fd_sc_hd__a22oi_1 _20858_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[26] ),
    .A2(net298),
    .B1(_13051_),
    .B2(net668),
    .Y(_13142_));
 sky130_fd_sc_hd__nor2_1 _20859_ (.A(_11040_),
    .B(_13142_),
    .Y(_13143_));
 sky130_fd_sc_hd__a21oi_1 _20860_ (.A1(_11040_),
    .A2(_13141_),
    .B1(_13143_),
    .Y(_13144_));
 sky130_fd_sc_hd__nor2_1 _20861_ (.A(_11726_),
    .B(_12974_),
    .Y(_13145_));
 sky130_fd_sc_hd__a21oi_1 _20862_ (.A1(\cs_registers_i.mtval_q[26] ),
    .A2(_12974_),
    .B1(_13145_),
    .Y(_13146_));
 sky130_fd_sc_hd__o22ai_1 _20863_ (.A1(_12998_),
    .A2(_13144_),
    .B1(_13146_),
    .B2(net278),
    .Y(_00405_));
 sky130_fd_sc_hd__nand2_1 _20864_ (.A(\cs_registers_i.pc_id_i[26] ),
    .B(_13140_),
    .Y(_13147_));
 sky130_fd_sc_hd__xnor2_1 _20865_ (.A(\cs_registers_i.pc_id_i[27] ),
    .B(_13147_),
    .Y(_13148_));
 sky130_fd_sc_hd__a22oi_1 _20866_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[27] ),
    .A2(net298),
    .B1(_13051_),
    .B2(net806),
    .Y(_13149_));
 sky130_fd_sc_hd__nor2_1 _20867_ (.A(_11040_),
    .B(_13149_),
    .Y(_13150_));
 sky130_fd_sc_hd__a21oi_1 _20868_ (.A1(_11040_),
    .A2(_13148_),
    .B1(_13150_),
    .Y(_13151_));
 sky130_fd_sc_hd__nor2_1 _20869_ (.A(_11746_),
    .B(_12974_),
    .Y(_13152_));
 sky130_fd_sc_hd__a21oi_1 _20870_ (.A1(\cs_registers_i.mtval_q[27] ),
    .A2(_12974_),
    .B1(_13152_),
    .Y(_13153_));
 sky130_fd_sc_hd__o22ai_1 _20871_ (.A1(_12998_),
    .A2(_13151_),
    .B1(_13153_),
    .B2(net278),
    .Y(_00406_));
 sky130_fd_sc_hd__nand3_1 _20872_ (.A(\cs_registers_i.pc_id_i[26] ),
    .B(\cs_registers_i.pc_id_i[27] ),
    .C(_13140_),
    .Y(_13154_));
 sky130_fd_sc_hd__xnor2_1 _20873_ (.A(\cs_registers_i.pc_id_i[28] ),
    .B(_13154_),
    .Y(_13155_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_542 ();
 sky130_fd_sc_hd__a22oi_1 _20875_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[28] ),
    .A2(net298),
    .B1(_13051_),
    .B2(net816),
    .Y(_13157_));
 sky130_fd_sc_hd__nor2_1 _20876_ (.A(_11040_),
    .B(_13157_),
    .Y(_13158_));
 sky130_fd_sc_hd__a21oi_2 _20877_ (.A1(_11040_),
    .A2(_13155_),
    .B1(_13158_),
    .Y(_13159_));
 sky130_fd_sc_hd__nor2_1 _20878_ (.A(_11765_),
    .B(_12974_),
    .Y(_13160_));
 sky130_fd_sc_hd__a21oi_1 _20879_ (.A1(\cs_registers_i.mtval_q[28] ),
    .A2(_12974_),
    .B1(_13160_),
    .Y(_13161_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_541 ();
 sky130_fd_sc_hd__o22ai_1 _20881_ (.A1(_12998_),
    .A2(_13159_),
    .B1(_13161_),
    .B2(net278),
    .Y(_00407_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_540 ();
 sky130_fd_sc_hd__inv_1 _20883_ (.A(\cs_registers_i.pc_id_i[28] ),
    .Y(_13164_));
 sky130_fd_sc_hd__nor2_1 _20884_ (.A(_13164_),
    .B(_13154_),
    .Y(_13165_));
 sky130_fd_sc_hd__xor2_1 _20885_ (.A(\cs_registers_i.pc_id_i[29] ),
    .B(_13165_),
    .X(_13166_));
 sky130_fd_sc_hd__a22oi_1 _20886_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[29] ),
    .A2(net298),
    .B1(_13051_),
    .B2(net671),
    .Y(_13167_));
 sky130_fd_sc_hd__nor2_1 _20887_ (.A(_11040_),
    .B(_13167_),
    .Y(_13168_));
 sky130_fd_sc_hd__a21oi_1 _20888_ (.A1(_11040_),
    .A2(_13166_),
    .B1(_13168_),
    .Y(_13169_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_539 ();
 sky130_fd_sc_hd__nor2_1 _20890_ (.A(_11785_),
    .B(_12974_),
    .Y(_13171_));
 sky130_fd_sc_hd__a21oi_1 _20891_ (.A1(\cs_registers_i.mtval_q[29] ),
    .A2(_12974_),
    .B1(_13171_),
    .Y(_13172_));
 sky130_fd_sc_hd__o22ai_1 _20892_ (.A1(_12998_),
    .A2(_13169_),
    .B1(_13172_),
    .B2(net278),
    .Y(_00408_));
 sky130_fd_sc_hd__nand2_1 _20893_ (.A(\cs_registers_i.pc_id_i[1] ),
    .B(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .Y(_13173_));
 sky130_fd_sc_hd__xnor2_1 _20894_ (.A(\cs_registers_i.pc_id_i[2] ),
    .B(_13173_),
    .Y(_13174_));
 sky130_fd_sc_hd__nand2_1 _20895_ (.A(\id_stage_i.controller_i.instr_is_compressed_i ),
    .B(\id_stage_i.controller_i.instr_compressed_i[2] ),
    .Y(_13175_));
 sky130_fd_sc_hd__o21ai_0 _20896_ (.A1(_08239_),
    .A2(\id_stage_i.controller_i.instr_is_compressed_i ),
    .B1(_13175_),
    .Y(_13176_));
 sky130_fd_sc_hd__a22oi_1 _20897_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[2] ),
    .A2(_12694_),
    .B1(_13176_),
    .B2(\id_stage_i.controller_i.illegal_insn_q ),
    .Y(_13177_));
 sky130_fd_sc_hd__nor2_1 _20898_ (.A(_11040_),
    .B(_13177_),
    .Y(_13178_));
 sky130_fd_sc_hd__a21oi_1 _20899_ (.A1(_11040_),
    .A2(_13174_),
    .B1(_13178_),
    .Y(_13179_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_538 ();
 sky130_fd_sc_hd__nor2_1 _20901_ (.A(_11309_),
    .B(_12974_),
    .Y(_13181_));
 sky130_fd_sc_hd__a21oi_1 _20902_ (.A1(\cs_registers_i.mtval_q[2] ),
    .A2(_12974_),
    .B1(_13181_),
    .Y(_13182_));
 sky130_fd_sc_hd__o22ai_1 _20903_ (.A1(_12998_),
    .A2(_13179_),
    .B1(_13182_),
    .B2(_12685_),
    .Y(_00409_));
 sky130_fd_sc_hd__nand2_1 _20904_ (.A(\cs_registers_i.pc_id_i[29] ),
    .B(_13165_),
    .Y(_13183_));
 sky130_fd_sc_hd__xnor2_1 _20905_ (.A(\cs_registers_i.pc_id_i[30] ),
    .B(_13183_),
    .Y(_13184_));
 sky130_fd_sc_hd__a22oi_1 _20906_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[30] ),
    .A2(net298),
    .B1(_13051_),
    .B2(net924),
    .Y(_13185_));
 sky130_fd_sc_hd__nor2_1 _20907_ (.A(_11040_),
    .B(_13185_),
    .Y(_13186_));
 sky130_fd_sc_hd__a21oi_1 _20908_ (.A1(_11040_),
    .A2(_13184_),
    .B1(_13186_),
    .Y(_13187_));
 sky130_fd_sc_hd__nor2_1 _20909_ (.A(_11808_),
    .B(_12974_),
    .Y(_13188_));
 sky130_fd_sc_hd__a21oi_1 _20910_ (.A1(\cs_registers_i.mtval_q[30] ),
    .A2(_12974_),
    .B1(_13188_),
    .Y(_13189_));
 sky130_fd_sc_hd__o22ai_1 _20911_ (.A1(_12998_),
    .A2(_13187_),
    .B1(_13189_),
    .B2(net279),
    .Y(_00410_));
 sky130_fd_sc_hd__nand3_1 _20912_ (.A(\cs_registers_i.pc_id_i[29] ),
    .B(\cs_registers_i.pc_id_i[30] ),
    .C(_13165_),
    .Y(_13190_));
 sky130_fd_sc_hd__xnor2_1 _20913_ (.A(\cs_registers_i.pc_id_i[31] ),
    .B(_13190_),
    .Y(_13191_));
 sky130_fd_sc_hd__a221o_1 _20914_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[31] ),
    .A2(net298),
    .B1(_13051_),
    .B2(net832),
    .C1(_11040_),
    .X(_13192_));
 sky130_fd_sc_hd__o21ai_0 _20915_ (.A1(_12731_),
    .A2(_13191_),
    .B1(_13192_),
    .Y(_13193_));
 sky130_fd_sc_hd__nor2_1 _20916_ (.A(_11826_),
    .B(_12974_),
    .Y(_13194_));
 sky130_fd_sc_hd__a21oi_1 _20917_ (.A1(\cs_registers_i.mtval_q[31] ),
    .A2(_12974_),
    .B1(_13194_),
    .Y(_13195_));
 sky130_fd_sc_hd__o22ai_1 _20918_ (.A1(_12998_),
    .A2(_13193_),
    .B1(_13195_),
    .B2(net279),
    .Y(_00411_));
 sky130_fd_sc_hd__xnor2_1 _20919_ (.A(\cs_registers_i.pc_id_i[3] ),
    .B(_12985_),
    .Y(_13196_));
 sky130_fd_sc_hd__nand2_1 _20920_ (.A(\id_stage_i.controller_i.instr_is_compressed_i ),
    .B(\id_stage_i.controller_i.instr_compressed_i[3] ),
    .Y(_13197_));
 sky130_fd_sc_hd__o21ai_0 _20921_ (.A1(_08234_),
    .A2(\id_stage_i.controller_i.instr_is_compressed_i ),
    .B1(_13197_),
    .Y(_13198_));
 sky130_fd_sc_hd__a22oi_1 _20922_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[3] ),
    .A2(_12694_),
    .B1(_13198_),
    .B2(\id_stage_i.controller_i.illegal_insn_q ),
    .Y(_13199_));
 sky130_fd_sc_hd__nor2_1 _20923_ (.A(_11040_),
    .B(_13199_),
    .Y(_13200_));
 sky130_fd_sc_hd__a21oi_2 _20924_ (.A1(_11040_),
    .A2(_13196_),
    .B1(_13200_),
    .Y(_13201_));
 sky130_fd_sc_hd__nor2_1 _20925_ (.A(_11867_),
    .B(_12974_),
    .Y(_13202_));
 sky130_fd_sc_hd__a21oi_1 _20926_ (.A1(\cs_registers_i.mtval_q[3] ),
    .A2(_12974_),
    .B1(_13202_),
    .Y(_13203_));
 sky130_fd_sc_hd__o22ai_1 _20927_ (.A1(_12998_),
    .A2(_13201_),
    .B1(_13203_),
    .B2(_12685_),
    .Y(_00412_));
 sky130_fd_sc_hd__xor2_1 _20928_ (.A(\cs_registers_i.pc_id_i[4] ),
    .B(_12986_),
    .X(_13204_));
 sky130_fd_sc_hd__mux2_1 _20929_ (.A0(\id_stage_i.controller_i.instr_i[4] ),
    .A1(\id_stage_i.controller_i.instr_compressed_i[4] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .X(_13205_));
 sky130_fd_sc_hd__a22oi_1 _20930_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[4] ),
    .A2(_12694_),
    .B1(_13205_),
    .B2(\id_stage_i.controller_i.illegal_insn_q ),
    .Y(_13206_));
 sky130_fd_sc_hd__nor2_1 _20931_ (.A(_11040_),
    .B(_13206_),
    .Y(_13207_));
 sky130_fd_sc_hd__a21oi_1 _20932_ (.A1(_11040_),
    .A2(_13204_),
    .B1(_13207_),
    .Y(_13208_));
 sky130_fd_sc_hd__nor2_1 _20933_ (.A(_11887_),
    .B(_12974_),
    .Y(_13209_));
 sky130_fd_sc_hd__a21oi_1 _20934_ (.A1(\cs_registers_i.mtval_q[4] ),
    .A2(_12974_),
    .B1(_13209_),
    .Y(_13210_));
 sky130_fd_sc_hd__o22ai_1 _20935_ (.A1(_12998_),
    .A2(_13208_),
    .B1(_13210_),
    .B2(_12685_),
    .Y(_00413_));
 sky130_fd_sc_hd__nand2_1 _20936_ (.A(\cs_registers_i.pc_id_i[4] ),
    .B(_12986_),
    .Y(_13211_));
 sky130_fd_sc_hd__xnor2_1 _20937_ (.A(\cs_registers_i.pc_id_i[5] ),
    .B(_13211_),
    .Y(_13212_));
 sky130_fd_sc_hd__mux2_1 _20938_ (.A0(net564),
    .A1(\id_stage_i.controller_i.instr_compressed_i[5] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .X(_13213_));
 sky130_fd_sc_hd__a22oi_1 _20939_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[5] ),
    .A2(_12694_),
    .B1(_13213_),
    .B2(\id_stage_i.controller_i.illegal_insn_q ),
    .Y(_13214_));
 sky130_fd_sc_hd__nor2_1 _20940_ (.A(_11040_),
    .B(_13214_),
    .Y(_13215_));
 sky130_fd_sc_hd__a21oi_2 _20941_ (.A1(_11040_),
    .A2(_13212_),
    .B1(_13215_),
    .Y(_13216_));
 sky130_fd_sc_hd__nor2_1 _20942_ (.A(_12594_),
    .B(_12974_),
    .Y(_13217_));
 sky130_fd_sc_hd__a21oi_1 _20943_ (.A1(\cs_registers_i.mtval_q[5] ),
    .A2(_12974_),
    .B1(_13217_),
    .Y(_13218_));
 sky130_fd_sc_hd__o22ai_1 _20944_ (.A1(_12998_),
    .A2(_13216_),
    .B1(_13218_),
    .B2(net277),
    .Y(_00414_));
 sky130_fd_sc_hd__xnor2_1 _20945_ (.A(_08545_),
    .B(_12987_),
    .Y(_13219_));
 sky130_fd_sc_hd__mux2_1 _20946_ (.A0(\id_stage_i.controller_i.instr_i[6] ),
    .A1(\id_stage_i.controller_i.instr_compressed_i[6] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .X(_13220_));
 sky130_fd_sc_hd__a22oi_1 _20947_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[6] ),
    .A2(_12694_),
    .B1(_13220_),
    .B2(\id_stage_i.controller_i.illegal_insn_q ),
    .Y(_13221_));
 sky130_fd_sc_hd__nor2_1 _20948_ (.A(_11040_),
    .B(_13221_),
    .Y(_13222_));
 sky130_fd_sc_hd__a21oi_1 _20949_ (.A1(_11040_),
    .A2(_13219_),
    .B1(_13222_),
    .Y(_13223_));
 sky130_fd_sc_hd__nor2_1 _20950_ (.A(_12113_),
    .B(_12974_),
    .Y(_13224_));
 sky130_fd_sc_hd__a21oi_1 _20951_ (.A1(\cs_registers_i.mtval_q[6] ),
    .A2(_12974_),
    .B1(_13224_),
    .Y(_13225_));
 sky130_fd_sc_hd__o22ai_1 _20952_ (.A1(_12998_),
    .A2(_13223_),
    .B1(_13225_),
    .B2(net277),
    .Y(_00415_));
 sky130_fd_sc_hd__nand2_1 _20953_ (.A(\cs_registers_i.pc_id_i[6] ),
    .B(_12987_),
    .Y(_13226_));
 sky130_fd_sc_hd__xnor2_1 _20954_ (.A(\cs_registers_i.pc_id_i[7] ),
    .B(_13226_),
    .Y(_13227_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_537 ();
 sky130_fd_sc_hd__mux2_1 _20956_ (.A0(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .A1(\id_stage_i.controller_i.instr_compressed_i[7] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .X(_13229_));
 sky130_fd_sc_hd__a22oi_1 _20957_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[7] ),
    .A2(_12694_),
    .B1(_13229_),
    .B2(\id_stage_i.controller_i.illegal_insn_q ),
    .Y(_13230_));
 sky130_fd_sc_hd__nor2_1 _20958_ (.A(_11040_),
    .B(_13230_),
    .Y(_13231_));
 sky130_fd_sc_hd__a21oi_1 _20959_ (.A1(_11040_),
    .A2(_13227_),
    .B1(_13231_),
    .Y(_13232_));
 sky130_fd_sc_hd__nor2_1 _20960_ (.A(_11935_),
    .B(_12974_),
    .Y(_13233_));
 sky130_fd_sc_hd__a21oi_1 _20961_ (.A1(\cs_registers_i.mtval_q[7] ),
    .A2(_12974_),
    .B1(_13233_),
    .Y(_13234_));
 sky130_fd_sc_hd__o22ai_1 _20962_ (.A1(_12998_),
    .A2(_13232_),
    .B1(_13234_),
    .B2(_12685_),
    .Y(_00416_));
 sky130_fd_sc_hd__xnor2_1 _20963_ (.A(\cs_registers_i.pc_id_i[8] ),
    .B(_12988_),
    .Y(_13235_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_536 ();
 sky130_fd_sc_hd__mux2_1 _20965_ (.A0(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .A1(\id_stage_i.controller_i.instr_compressed_i[8] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .X(_13237_));
 sky130_fd_sc_hd__a22oi_1 _20966_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[8] ),
    .A2(_12694_),
    .B1(_13237_),
    .B2(\id_stage_i.controller_i.illegal_insn_q ),
    .Y(_13238_));
 sky130_fd_sc_hd__nor2_1 _20967_ (.A(_11040_),
    .B(_13238_),
    .Y(_13239_));
 sky130_fd_sc_hd__a21oi_1 _20968_ (.A1(_11040_),
    .A2(_13235_),
    .B1(_13239_),
    .Y(_13240_));
 sky130_fd_sc_hd__nor2_1 _20969_ (.A(_11957_),
    .B(_12974_),
    .Y(_13241_));
 sky130_fd_sc_hd__a21oi_1 _20970_ (.A1(\cs_registers_i.mtval_q[8] ),
    .A2(_12974_),
    .B1(_13241_),
    .Y(_13242_));
 sky130_fd_sc_hd__o22ai_1 _20971_ (.A1(_12998_),
    .A2(_13240_),
    .B1(_13242_),
    .B2(net277),
    .Y(_00417_));
 sky130_fd_sc_hd__xnor2_1 _20972_ (.A(_09288_),
    .B(_12989_),
    .Y(_13243_));
 sky130_fd_sc_hd__mux2_1 _20973_ (.A0(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .A1(\id_stage_i.controller_i.instr_compressed_i[9] ),
    .S(\id_stage_i.controller_i.instr_is_compressed_i ),
    .X(_13244_));
 sky130_fd_sc_hd__a22oi_1 _20974_ (.A1(\id_stage_i.controller_i.lsu_addr_last_i[9] ),
    .A2(_12694_),
    .B1(_13244_),
    .B2(\id_stage_i.controller_i.illegal_insn_q ),
    .Y(_13245_));
 sky130_fd_sc_hd__nor2_1 _20975_ (.A(_11040_),
    .B(_13245_),
    .Y(_13246_));
 sky130_fd_sc_hd__a21oi_1 _20976_ (.A1(_11040_),
    .A2(_13243_),
    .B1(_13246_),
    .Y(_13247_));
 sky130_fd_sc_hd__nor2_1 _20977_ (.A(_11973_),
    .B(_12974_),
    .Y(_13248_));
 sky130_fd_sc_hd__a21oi_1 _20978_ (.A1(\cs_registers_i.mtval_q[9] ),
    .A2(_12974_),
    .B1(_13248_),
    .Y(_13249_));
 sky130_fd_sc_hd__o22ai_1 _20979_ (.A1(_12998_),
    .A2(_13247_),
    .B1(_13249_),
    .B2(_12685_),
    .Y(_00418_));
 sky130_fd_sc_hd__inv_1 _20980_ (.A(_10918_),
    .Y(_13250_));
 sky130_fd_sc_hd__o21ai_4 _20981_ (.A1(_13250_),
    .A2(_11313_),
    .B1(_11006_),
    .Y(_13251_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_533 ();
 sky130_fd_sc_hd__mux2i_1 _20985_ (.A0(net1),
    .A1(_11357_),
    .S(_11006_),
    .Y(_13255_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_532 ();
 sky130_fd_sc_hd__nor2_1 _20987_ (.A(\cs_registers_i.csr_mtvec_o[10] ),
    .B(net1018),
    .Y(_13257_));
 sky130_fd_sc_hd__a21oi_1 _20988_ (.A1(net1018),
    .A2(_13255_),
    .B1(_13257_),
    .Y(_00419_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_530 ();
 sky130_fd_sc_hd__nand2_1 _20991_ (.A(_11006_),
    .B(_12481_),
    .Y(_13260_));
 sky130_fd_sc_hd__o21ai_0 _20992_ (.A1(net2),
    .A2(_11006_),
    .B1(_13260_),
    .Y(_13261_));
 sky130_fd_sc_hd__nor2_1 _20993_ (.A(\cs_registers_i.csr_mtvec_o[11] ),
    .B(net1018),
    .Y(_13262_));
 sky130_fd_sc_hd__a21oi_1 _20994_ (.A1(net1018),
    .A2(_13261_),
    .B1(_13262_),
    .Y(_00420_));
 sky130_fd_sc_hd__nand2_1 _20995_ (.A(_11006_),
    .B(_11428_),
    .Y(_13263_));
 sky130_fd_sc_hd__o21ai_0 _20996_ (.A1(net3),
    .A2(_11006_),
    .B1(_13263_),
    .Y(_13264_));
 sky130_fd_sc_hd__nor2_1 _20997_ (.A(\cs_registers_i.csr_mtvec_o[12] ),
    .B(net1018),
    .Y(_13265_));
 sky130_fd_sc_hd__a21oi_1 _20998_ (.A1(net1018),
    .A2(_13264_),
    .B1(_13265_),
    .Y(_00421_));
 sky130_fd_sc_hd__nand2_1 _20999_ (.A(_11006_),
    .B(_11448_),
    .Y(_13266_));
 sky130_fd_sc_hd__o21ai_0 _21000_ (.A1(net4),
    .A2(_11006_),
    .B1(_13266_),
    .Y(_13267_));
 sky130_fd_sc_hd__nor2_1 _21001_ (.A(\cs_registers_i.csr_mtvec_o[13] ),
    .B(net1018),
    .Y(_13268_));
 sky130_fd_sc_hd__a21oi_1 _21002_ (.A1(net1018),
    .A2(_13267_),
    .B1(_13268_),
    .Y(_00422_));
 sky130_fd_sc_hd__nand2_1 _21003_ (.A(_11006_),
    .B(_11465_),
    .Y(_13269_));
 sky130_fd_sc_hd__o21ai_0 _21004_ (.A1(net5),
    .A2(_11006_),
    .B1(_13269_),
    .Y(_13270_));
 sky130_fd_sc_hd__nor2_1 _21005_ (.A(\cs_registers_i.csr_mtvec_o[14] ),
    .B(net1018),
    .Y(_13271_));
 sky130_fd_sc_hd__a21oi_1 _21006_ (.A1(net1018),
    .A2(_13270_),
    .B1(_13271_),
    .Y(_00423_));
 sky130_fd_sc_hd__nand2_1 _21007_ (.A(_11006_),
    .B(_11488_),
    .Y(_13272_));
 sky130_fd_sc_hd__o21ai_0 _21008_ (.A1(net6),
    .A2(_11006_),
    .B1(_13272_),
    .Y(_13273_));
 sky130_fd_sc_hd__nor2_1 _21009_ (.A(\cs_registers_i.csr_mtvec_o[15] ),
    .B(net1018),
    .Y(_13274_));
 sky130_fd_sc_hd__a21oi_1 _21010_ (.A1(net1018),
    .A2(_13273_),
    .B1(_13274_),
    .Y(_00424_));
 sky130_fd_sc_hd__nand2_1 _21011_ (.A(_11006_),
    .B(_11505_),
    .Y(_13275_));
 sky130_fd_sc_hd__o21ai_0 _21012_ (.A1(net7),
    .A2(_11006_),
    .B1(_13275_),
    .Y(_13276_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_529 ();
 sky130_fd_sc_hd__nor2_1 _21014_ (.A(\cs_registers_i.csr_mtvec_o[16] ),
    .B(_13251_),
    .Y(_13278_));
 sky130_fd_sc_hd__a21oi_1 _21015_ (.A1(_13251_),
    .A2(_13276_),
    .B1(_13278_),
    .Y(_00425_));
 sky130_fd_sc_hd__nand2_1 _21016_ (.A(_11006_),
    .B(_11523_),
    .Y(_13279_));
 sky130_fd_sc_hd__o21ai_0 _21017_ (.A1(net8),
    .A2(_11006_),
    .B1(_13279_),
    .Y(_13280_));
 sky130_fd_sc_hd__nor2_1 _21018_ (.A(\cs_registers_i.csr_mtvec_o[17] ),
    .B(_13251_),
    .Y(_13281_));
 sky130_fd_sc_hd__a21oi_1 _21019_ (.A1(_13251_),
    .A2(_13280_),
    .B1(_13281_),
    .Y(_00426_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_528 ();
 sky130_fd_sc_hd__nand2_1 _21021_ (.A(_11006_),
    .B(_11546_),
    .Y(_13283_));
 sky130_fd_sc_hd__o21ai_0 _21022_ (.A1(net9),
    .A2(_11006_),
    .B1(_13283_),
    .Y(_13284_));
 sky130_fd_sc_hd__nor2_1 _21023_ (.A(\cs_registers_i.csr_mtvec_o[18] ),
    .B(_13251_),
    .Y(_13285_));
 sky130_fd_sc_hd__a21oi_1 _21024_ (.A1(_13251_),
    .A2(_13284_),
    .B1(_13285_),
    .Y(_00427_));
 sky130_fd_sc_hd__nand2_1 _21025_ (.A(_11006_),
    .B(_11563_),
    .Y(_13286_));
 sky130_fd_sc_hd__o21ai_0 _21026_ (.A1(net10),
    .A2(_11006_),
    .B1(_13286_),
    .Y(_13287_));
 sky130_fd_sc_hd__nor2_1 _21027_ (.A(\cs_registers_i.csr_mtvec_o[19] ),
    .B(_13251_),
    .Y(_13288_));
 sky130_fd_sc_hd__a21oi_1 _21028_ (.A1(_13251_),
    .A2(_13287_),
    .B1(_13288_),
    .Y(_00428_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_527 ();
 sky130_fd_sc_hd__nand2_1 _21030_ (.A(_11006_),
    .B(_11599_),
    .Y(_13290_));
 sky130_fd_sc_hd__o21ai_0 _21031_ (.A1(net11),
    .A2(_11006_),
    .B1(_13290_),
    .Y(_13291_));
 sky130_fd_sc_hd__nor2_1 _21032_ (.A(\cs_registers_i.csr_mtvec_o[20] ),
    .B(net1018),
    .Y(_13292_));
 sky130_fd_sc_hd__a21oi_1 _21033_ (.A1(net1018),
    .A2(_13291_),
    .B1(_13292_),
    .Y(_00429_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_526 ();
 sky130_fd_sc_hd__nand2_1 _21035_ (.A(_11006_),
    .B(_11623_),
    .Y(_13294_));
 sky130_fd_sc_hd__o21ai_0 _21036_ (.A1(net12),
    .A2(_11006_),
    .B1(_13294_),
    .Y(_13295_));
 sky130_fd_sc_hd__nor2_1 _21037_ (.A(\cs_registers_i.csr_mtvec_o[21] ),
    .B(net1018),
    .Y(_13296_));
 sky130_fd_sc_hd__a21oi_1 _21038_ (.A1(net1018),
    .A2(_13295_),
    .B1(_13296_),
    .Y(_00430_));
 sky130_fd_sc_hd__nand2_1 _21039_ (.A(_11006_),
    .B(_11643_),
    .Y(_13297_));
 sky130_fd_sc_hd__o21ai_0 _21040_ (.A1(net13),
    .A2(_11006_),
    .B1(_13297_),
    .Y(_13298_));
 sky130_fd_sc_hd__nor2_1 _21041_ (.A(\cs_registers_i.csr_mtvec_o[22] ),
    .B(net1018),
    .Y(_13299_));
 sky130_fd_sc_hd__a21oi_1 _21042_ (.A1(net1018),
    .A2(_13298_),
    .B1(_13299_),
    .Y(_00431_));
 sky130_fd_sc_hd__nand2_1 _21043_ (.A(_11006_),
    .B(_11664_),
    .Y(_13300_));
 sky130_fd_sc_hd__o21ai_0 _21044_ (.A1(net14),
    .A2(_11006_),
    .B1(_13300_),
    .Y(_13301_));
 sky130_fd_sc_hd__nor2_1 _21045_ (.A(\cs_registers_i.csr_mtvec_o[23] ),
    .B(net1018),
    .Y(_13302_));
 sky130_fd_sc_hd__a21oi_1 _21046_ (.A1(net1018),
    .A2(_13301_),
    .B1(_13302_),
    .Y(_00432_));
 sky130_fd_sc_hd__nand2_1 _21047_ (.A(_11006_),
    .B(_11684_),
    .Y(_13303_));
 sky130_fd_sc_hd__o21ai_0 _21048_ (.A1(net15),
    .A2(_11006_),
    .B1(_13303_),
    .Y(_13304_));
 sky130_fd_sc_hd__nor2_1 _21049_ (.A(\cs_registers_i.csr_mtvec_o[24] ),
    .B(_13251_),
    .Y(_13305_));
 sky130_fd_sc_hd__a21oi_1 _21050_ (.A1(_13251_),
    .A2(_13304_),
    .B1(_13305_),
    .Y(_00433_));
 sky130_fd_sc_hd__nand2_1 _21051_ (.A(_11006_),
    .B(_11706_),
    .Y(_13306_));
 sky130_fd_sc_hd__o21ai_0 _21052_ (.A1(net16),
    .A2(_11006_),
    .B1(_13306_),
    .Y(_13307_));
 sky130_fd_sc_hd__nor2_1 _21053_ (.A(\cs_registers_i.csr_mtvec_o[25] ),
    .B(net1018),
    .Y(_13308_));
 sky130_fd_sc_hd__a21oi_1 _21054_ (.A1(net1018),
    .A2(_13307_),
    .B1(_13308_),
    .Y(_00434_));
 sky130_fd_sc_hd__nand2_1 _21055_ (.A(_11006_),
    .B(_11726_),
    .Y(_13309_));
 sky130_fd_sc_hd__o21ai_0 _21056_ (.A1(net17),
    .A2(_11006_),
    .B1(_13309_),
    .Y(_13310_));
 sky130_fd_sc_hd__nor2_1 _21057_ (.A(\cs_registers_i.csr_mtvec_o[26] ),
    .B(_13251_),
    .Y(_13311_));
 sky130_fd_sc_hd__a21oi_1 _21058_ (.A1(_13251_),
    .A2(_13310_),
    .B1(_13311_),
    .Y(_00435_));
 sky130_fd_sc_hd__nand2_1 _21059_ (.A(_11006_),
    .B(_11746_),
    .Y(_13312_));
 sky130_fd_sc_hd__o21ai_0 _21060_ (.A1(net18),
    .A2(_11006_),
    .B1(_13312_),
    .Y(_13313_));
 sky130_fd_sc_hd__nor2_1 _21061_ (.A(\cs_registers_i.csr_mtvec_o[27] ),
    .B(_13251_),
    .Y(_13314_));
 sky130_fd_sc_hd__a21oi_1 _21062_ (.A1(net1018),
    .A2(_13313_),
    .B1(_13314_),
    .Y(_00436_));
 sky130_fd_sc_hd__nand2_1 _21063_ (.A(_11006_),
    .B(_11765_),
    .Y(_13315_));
 sky130_fd_sc_hd__o21ai_0 _21064_ (.A1(net19),
    .A2(_11006_),
    .B1(_13315_),
    .Y(_13316_));
 sky130_fd_sc_hd__nor2_1 _21065_ (.A(\cs_registers_i.csr_mtvec_o[28] ),
    .B(_13251_),
    .Y(_13317_));
 sky130_fd_sc_hd__a21oi_1 _21066_ (.A1(_13251_),
    .A2(_13316_),
    .B1(_13317_),
    .Y(_00437_));
 sky130_fd_sc_hd__nand2_1 _21067_ (.A(_11006_),
    .B(_11785_),
    .Y(_13318_));
 sky130_fd_sc_hd__o21ai_0 _21068_ (.A1(net20),
    .A2(_11006_),
    .B1(_13318_),
    .Y(_13319_));
 sky130_fd_sc_hd__nor2_1 _21069_ (.A(\cs_registers_i.csr_mtvec_o[29] ),
    .B(_13251_),
    .Y(_13320_));
 sky130_fd_sc_hd__a21oi_1 _21070_ (.A1(_13251_),
    .A2(_13319_),
    .B1(_13320_),
    .Y(_00438_));
 sky130_fd_sc_hd__nand2_1 _21071_ (.A(_11006_),
    .B(_11808_),
    .Y(_13321_));
 sky130_fd_sc_hd__o21ai_0 _21072_ (.A1(net21),
    .A2(_11006_),
    .B1(_13321_),
    .Y(_13322_));
 sky130_fd_sc_hd__nor2_1 _21073_ (.A(\cs_registers_i.csr_mtvec_o[30] ),
    .B(net1018),
    .Y(_13323_));
 sky130_fd_sc_hd__a21oi_1 _21074_ (.A1(net1018),
    .A2(_13322_),
    .B1(_13323_),
    .Y(_00439_));
 sky130_fd_sc_hd__nand2_1 _21075_ (.A(_11006_),
    .B(_11826_),
    .Y(_13324_));
 sky130_fd_sc_hd__o21ai_0 _21076_ (.A1(net22),
    .A2(_11006_),
    .B1(_13324_),
    .Y(_13325_));
 sky130_fd_sc_hd__nor2_1 _21077_ (.A(\cs_registers_i.csr_mtvec_o[31] ),
    .B(_13251_),
    .Y(_13326_));
 sky130_fd_sc_hd__a21oi_1 _21078_ (.A1(_13251_),
    .A2(_13325_),
    .B1(_13326_),
    .Y(_00440_));
 sky130_fd_sc_hd__nand2_1 _21079_ (.A(_11006_),
    .B(_11957_),
    .Y(_13327_));
 sky130_fd_sc_hd__o21ai_0 _21080_ (.A1(net23),
    .A2(_11006_),
    .B1(_13327_),
    .Y(_13328_));
 sky130_fd_sc_hd__nor2_1 _21081_ (.A(\cs_registers_i.csr_mtvec_o[8] ),
    .B(net1018),
    .Y(_13329_));
 sky130_fd_sc_hd__a21oi_1 _21082_ (.A1(net1018),
    .A2(_13328_),
    .B1(_13329_),
    .Y(_00441_));
 sky130_fd_sc_hd__nand2_1 _21083_ (.A(_11006_),
    .B(_11973_),
    .Y(_13330_));
 sky130_fd_sc_hd__o21ai_0 _21084_ (.A1(net24),
    .A2(_11006_),
    .B1(_13330_),
    .Y(_13331_));
 sky130_fd_sc_hd__nor2_1 _21085_ (.A(\cs_registers_i.csr_mtvec_o[9] ),
    .B(net1018),
    .Y(_13332_));
 sky130_fd_sc_hd__a21oi_1 _21086_ (.A1(net1018),
    .A2(_13331_),
    .B1(_13332_),
    .Y(_00442_));
 sky130_fd_sc_hd__nor2_4 _21087_ (.A(net445),
    .B(_10950_),
    .Y(_13333_));
 sky130_fd_sc_hd__nand3_1 _21088_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .B(_10951_),
    .C(_13333_),
    .Y(_13334_));
 sky130_fd_sc_hd__mux2_1 _21089_ (.A0(_10988_),
    .A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_by_zero_q ),
    .S(_13334_),
    .X(_00443_));
 sky130_fd_sc_hd__nor2_8 _21090_ (.A(_08100_),
    .B(net739),
    .Y(_13335_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_525 ();
 sky130_fd_sc_hd__nor3_2 _21092_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .C(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .Y(_13337_));
 sky130_fd_sc_hd__and3_1 _21093_ (.A(net1524),
    .B(_13335_),
    .C(_13337_),
    .X(_13338_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_524 ();
 sky130_fd_sc_hd__a21oi_1 _21095_ (.A1(net1524),
    .A2(_13335_),
    .B1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_13340_));
 sky130_fd_sc_hd__a21oi_1 _21096_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .A2(_13338_),
    .B1(_13340_),
    .Y(_00444_));
 sky130_fd_sc_hd__nor2b_1 _21097_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B_N(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .Y(_13341_));
 sky130_fd_sc_hd__nand2_1 _21098_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B(_13337_),
    .Y(_13342_));
 sky130_fd_sc_hd__a21oi_1 _21099_ (.A1(_10951_),
    .A2(_13342_),
    .B1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .Y(_13343_));
 sky130_fd_sc_hd__a21oi_1 _21100_ (.A1(_13338_),
    .A2(_13341_),
    .B1(_13343_),
    .Y(_00445_));
 sky130_fd_sc_hd__nor2_2 _21101_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_13344_));
 sky130_fd_sc_hd__or2_4 _21102_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .X(_13345_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_523 ();
 sky130_fd_sc_hd__nand2_1 _21104_ (.A(_13337_),
    .B(_13345_),
    .Y(_13347_));
 sky130_fd_sc_hd__a21oi_1 _21105_ (.A1(_10951_),
    .A2(_13347_),
    .B1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .Y(_13348_));
 sky130_fd_sc_hd__a31oi_1 _21106_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .A2(_13338_),
    .A3(_13344_),
    .B1(_13348_),
    .Y(_00446_));
 sky130_fd_sc_hd__o21a_1 _21107_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .A2(_13345_),
    .B1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .X(_13349_));
 sky130_fd_sc_hd__nor3_4 _21108_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .C(_13345_),
    .Y(_13350_));
 sky130_fd_sc_hd__nor2_2 _21109_ (.A(_13349_),
    .B(_13350_),
    .Y(_13351_));
 sky130_fd_sc_hd__nor2_1 _21110_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .B(_10951_),
    .Y(_13352_));
 sky130_fd_sc_hd__a31oi_1 _21111_ (.A1(_10951_),
    .A2(_13337_),
    .A3(_13351_),
    .B1(_13352_),
    .Y(_00447_));
 sky130_fd_sc_hd__nand2b_1 _21112_ (.A_N(_13350_),
    .B(_13337_),
    .Y(_13353_));
 sky130_fd_sc_hd__a21oi_1 _21113_ (.A1(_10951_),
    .A2(_13353_),
    .B1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .Y(_13354_));
 sky130_fd_sc_hd__a31oi_1 _21114_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .A2(_13338_),
    .A3(_13350_),
    .B1(_13354_),
    .Y(_00448_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_521 ();
 sky130_fd_sc_hd__o21ai_4 _21117_ (.A1(net665),
    .A2(_08231_),
    .B1(net491),
    .Y(_13357_));
 sky130_fd_sc_hd__and3_4 _21118_ (.A(net316),
    .B(_10691_),
    .C(_13357_),
    .X(_13358_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_519 ();
 sky130_fd_sc_hd__mux2i_1 _21121_ (.A0(net497),
    .A1(net288),
    .S(_13358_),
    .Y(_13361_));
 sky130_fd_sc_hd__nand2_1 _21122_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[0] ),
    .B(_11214_),
    .Y(_13362_));
 sky130_fd_sc_hd__o21ai_0 _21123_ (.A1(_11214_),
    .A2(_13361_),
    .B1(_13362_),
    .Y(_00449_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_517 ();
 sky130_fd_sc_hd__nor2_1 _21126_ (.A(_09380_),
    .B(_13358_),
    .Y(_13365_));
 sky130_fd_sc_hd__a21oi_1 _21127_ (.A1(net1578),
    .A2(_13358_),
    .B1(_13365_),
    .Y(_13366_));
 sky130_fd_sc_hd__nand2_1 _21128_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[10] ),
    .B(_11214_),
    .Y(_13367_));
 sky130_fd_sc_hd__o21ai_0 _21129_ (.A1(_11214_),
    .A2(_13366_),
    .B1(_13367_),
    .Y(_00450_));
 sky130_fd_sc_hd__mux2i_1 _21130_ (.A0(net1189),
    .A1(net152),
    .S(_13358_),
    .Y(_13368_));
 sky130_fd_sc_hd__nand2_1 _21131_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[11] ),
    .B(_11214_),
    .Y(_13369_));
 sky130_fd_sc_hd__o21ai_0 _21132_ (.A1(_11214_),
    .A2(_13368_),
    .B1(_13369_),
    .Y(_00451_));
 sky130_fd_sc_hd__nor2_1 _21133_ (.A(_09553_),
    .B(_13358_),
    .Y(_13370_));
 sky130_fd_sc_hd__a21oi_1 _21134_ (.A1(net153),
    .A2(_13358_),
    .B1(_13370_),
    .Y(_13371_));
 sky130_fd_sc_hd__nand2_1 _21135_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[12] ),
    .B(_11214_),
    .Y(_13372_));
 sky130_fd_sc_hd__o21ai_0 _21136_ (.A1(_11214_),
    .A2(_13371_),
    .B1(_13372_),
    .Y(_00452_));
 sky130_fd_sc_hd__nor2_1 _21137_ (.A(net648),
    .B(_13358_),
    .Y(_13373_));
 sky130_fd_sc_hd__a21oi_1 _21138_ (.A1(net154),
    .A2(_13358_),
    .B1(_13373_),
    .Y(_13374_));
 sky130_fd_sc_hd__nand2_1 _21139_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[13] ),
    .B(_11214_),
    .Y(_13375_));
 sky130_fd_sc_hd__o21ai_0 _21140_ (.A1(_11214_),
    .A2(_13374_),
    .B1(_13375_),
    .Y(_00453_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_516 ();
 sky130_fd_sc_hd__nor2_1 _21142_ (.A(_09632_),
    .B(_13358_),
    .Y(_13377_));
 sky130_fd_sc_hd__a21oi_1 _21143_ (.A1(net1583),
    .A2(_13358_),
    .B1(_13377_),
    .Y(_13378_));
 sky130_fd_sc_hd__nand2_1 _21144_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[14] ),
    .B(_11214_),
    .Y(_13379_));
 sky130_fd_sc_hd__o21ai_0 _21145_ (.A1(_11214_),
    .A2(_13378_),
    .B1(_13379_),
    .Y(_00454_));
 sky130_fd_sc_hd__mux2i_1 _21146_ (.A0(net838),
    .A1(net721),
    .S(_13358_),
    .Y(_13380_));
 sky130_fd_sc_hd__nand2_1 _21147_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[15] ),
    .B(_11214_),
    .Y(_13381_));
 sky130_fd_sc_hd__o21ai_0 _21148_ (.A1(_11214_),
    .A2(_13380_),
    .B1(_13381_),
    .Y(_00455_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_515 ();
 sky130_fd_sc_hd__nor2_1 _21150_ (.A(_09821_),
    .B(_13358_),
    .Y(_13383_));
 sky130_fd_sc_hd__a21oi_1 _21151_ (.A1(net1581),
    .A2(_13358_),
    .B1(_13383_),
    .Y(_13384_));
 sky130_fd_sc_hd__nand2_1 _21152_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[16] ),
    .B(_11214_),
    .Y(_13385_));
 sky130_fd_sc_hd__o21ai_0 _21153_ (.A1(_11214_),
    .A2(_13384_),
    .B1(_13385_),
    .Y(_00456_));
 sky130_fd_sc_hd__mux2i_1 _21154_ (.A0(net776),
    .A1(net1560),
    .S(_13358_),
    .Y(_13386_));
 sky130_fd_sc_hd__nand2_1 _21155_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[17] ),
    .B(_11214_),
    .Y(_13387_));
 sky130_fd_sc_hd__o21ai_0 _21156_ (.A1(_11214_),
    .A2(_13386_),
    .B1(_13387_),
    .Y(_00457_));
 sky130_fd_sc_hd__mux2i_1 _21157_ (.A0(net961),
    .A1(net1241),
    .S(_13358_),
    .Y(_13388_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_514 ();
 sky130_fd_sc_hd__nand2_1 _21159_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[18] ),
    .B(_11214_),
    .Y(_13390_));
 sky130_fd_sc_hd__o21ai_0 _21160_ (.A1(_11214_),
    .A2(_13388_),
    .B1(_13390_),
    .Y(_00458_));
 sky130_fd_sc_hd__nor2_1 _21161_ (.A(_09969_),
    .B(_13358_),
    .Y(_13391_));
 sky130_fd_sc_hd__a21oi_1 _21162_ (.A1(net1260),
    .A2(_13358_),
    .B1(_13391_),
    .Y(_13392_));
 sky130_fd_sc_hd__nand2_1 _21163_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[19] ),
    .B(_11214_),
    .Y(_13393_));
 sky130_fd_sc_hd__o21ai_0 _21164_ (.A1(_11214_),
    .A2(_13392_),
    .B1(_13393_),
    .Y(_00459_));
 sky130_fd_sc_hd__xor2_4 _21165_ (.A(net987),
    .B(_10969_),
    .X(_13394_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_513 ();
 sky130_fd_sc_hd__nand2_1 _21167_ (.A(net276),
    .B(_13358_),
    .Y(_13396_));
 sky130_fd_sc_hd__o21ai_0 _21168_ (.A1(net561),
    .A2(_13358_),
    .B1(_13396_),
    .Y(_13397_));
 sky130_fd_sc_hd__nand2_1 _21169_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[1] ),
    .B(_11214_),
    .Y(_13398_));
 sky130_fd_sc_hd__o21ai_0 _21170_ (.A1(_11214_),
    .A2(_13397_),
    .B1(_13398_),
    .Y(_00460_));
 sky130_fd_sc_hd__nor2_1 _21171_ (.A(_10061_),
    .B(_13358_),
    .Y(_13399_));
 sky130_fd_sc_hd__a21oi_1 _21172_ (.A1(net691),
    .A2(_13358_),
    .B1(_13399_),
    .Y(_13400_));
 sky130_fd_sc_hd__nand2_1 _21173_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[20] ),
    .B(_11214_),
    .Y(_13401_));
 sky130_fd_sc_hd__o21ai_0 _21174_ (.A1(_11214_),
    .A2(_13400_),
    .B1(_13401_),
    .Y(_00461_));
 sky130_fd_sc_hd__nor2_1 _21175_ (.A(_10130_),
    .B(_13358_),
    .Y(_13402_));
 sky130_fd_sc_hd__a21oi_1 _21176_ (.A1(net1257),
    .A2(_13358_),
    .B1(_13402_),
    .Y(_13403_));
 sky130_fd_sc_hd__nand2_1 _21177_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[21] ),
    .B(_11214_),
    .Y(_13404_));
 sky130_fd_sc_hd__o21ai_0 _21178_ (.A1(_11214_),
    .A2(_13403_),
    .B1(_13404_),
    .Y(_00462_));
 sky130_fd_sc_hd__nor2_1 _21179_ (.A(_10168_),
    .B(_13358_),
    .Y(_13405_));
 sky130_fd_sc_hd__a21oi_1 _21180_ (.A1(net993),
    .A2(_13358_),
    .B1(_13405_),
    .Y(_13406_));
 sky130_fd_sc_hd__nand2_1 _21181_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[22] ),
    .B(_11214_),
    .Y(_13407_));
 sky130_fd_sc_hd__o21ai_0 _21182_ (.A1(_11214_),
    .A2(_13406_),
    .B1(_13407_),
    .Y(_00463_));
 sky130_fd_sc_hd__nor2_1 _21183_ (.A(_10232_),
    .B(_13358_),
    .Y(_13408_));
 sky130_fd_sc_hd__a21oi_1 _21184_ (.A1(net164),
    .A2(_13358_),
    .B1(_13408_),
    .Y(_13409_));
 sky130_fd_sc_hd__nand2_1 _21185_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[23] ),
    .B(_11214_),
    .Y(_13410_));
 sky130_fd_sc_hd__o21ai_0 _21186_ (.A1(_11214_),
    .A2(_13409_),
    .B1(_13410_),
    .Y(_00464_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_512 ();
 sky130_fd_sc_hd__nor2_1 _21188_ (.A(_10365_),
    .B(_13358_),
    .Y(_13412_));
 sky130_fd_sc_hd__a21oi_1 _21189_ (.A1(net165),
    .A2(_13358_),
    .B1(_13412_),
    .Y(_13413_));
 sky130_fd_sc_hd__nand2_1 _21190_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[24] ),
    .B(_11214_),
    .Y(_13414_));
 sky130_fd_sc_hd__o21ai_0 _21191_ (.A1(_11214_),
    .A2(_13413_),
    .B1(_13414_),
    .Y(_00465_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_511 ();
 sky130_fd_sc_hd__nor2_1 _21193_ (.A(_10299_),
    .B(_13358_),
    .Y(_13416_));
 sky130_fd_sc_hd__a21oi_1 _21194_ (.A1(net166),
    .A2(_13358_),
    .B1(_13416_),
    .Y(_13417_));
 sky130_fd_sc_hd__nand2_1 _21195_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[25] ),
    .B(_11214_),
    .Y(_13418_));
 sky130_fd_sc_hd__o21ai_0 _21196_ (.A1(_11214_),
    .A2(_13417_),
    .B1(_13418_),
    .Y(_00466_));
 sky130_fd_sc_hd__nor2_1 _21197_ (.A(_10457_),
    .B(_13358_),
    .Y(_13419_));
 sky130_fd_sc_hd__a21oi_1 _21198_ (.A1(net167),
    .A2(_13358_),
    .B1(_13419_),
    .Y(_13420_));
 sky130_fd_sc_hd__nand2_1 _21199_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[26] ),
    .B(_11214_),
    .Y(_13421_));
 sky130_fd_sc_hd__o21ai_0 _21200_ (.A1(_11214_),
    .A2(_13420_),
    .B1(_13421_),
    .Y(_00467_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_510 ();
 sky130_fd_sc_hd__nor2_1 _21202_ (.A(_10493_),
    .B(_13358_),
    .Y(_13423_));
 sky130_fd_sc_hd__a21oi_1 _21203_ (.A1(net688),
    .A2(_13358_),
    .B1(_13423_),
    .Y(_13424_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_509 ();
 sky130_fd_sc_hd__nand2_1 _21205_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[27] ),
    .B(_11214_),
    .Y(_13426_));
 sky130_fd_sc_hd__o21ai_0 _21206_ (.A1(_11214_),
    .A2(_13424_),
    .B1(_13426_),
    .Y(_00468_));
 sky130_fd_sc_hd__nor2_1 _21207_ (.A(_10644_),
    .B(_13358_),
    .Y(_13427_));
 sky130_fd_sc_hd__a21oi_1 _21208_ (.A1(net494),
    .A2(_13358_),
    .B1(_13427_),
    .Y(_13428_));
 sky130_fd_sc_hd__nand2_1 _21209_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[28] ),
    .B(_11214_),
    .Y(_13429_));
 sky130_fd_sc_hd__o21ai_0 _21210_ (.A1(_11214_),
    .A2(_13428_),
    .B1(_13429_),
    .Y(_00469_));
 sky130_fd_sc_hd__nor2_1 _21211_ (.A(_10557_),
    .B(_13358_),
    .Y(_13430_));
 sky130_fd_sc_hd__a21oi_1 _21212_ (.A1(net170),
    .A2(_13358_),
    .B1(_13430_),
    .Y(_13431_));
 sky130_fd_sc_hd__nand2_1 _21213_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[29] ),
    .B(_11214_),
    .Y(_13432_));
 sky130_fd_sc_hd__o21ai_0 _21214_ (.A1(_11214_),
    .A2(_13431_),
    .B1(_13432_),
    .Y(_00470_));
 sky130_fd_sc_hd__nor2_1 _21215_ (.A(net751),
    .B(_13358_),
    .Y(_13433_));
 sky130_fd_sc_hd__a21oi_1 _21216_ (.A1(net171),
    .A2(_13358_),
    .B1(_13433_),
    .Y(_13434_));
 sky130_fd_sc_hd__nand2_1 _21217_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[2] ),
    .B(_11214_),
    .Y(_13435_));
 sky130_fd_sc_hd__o21ai_0 _21218_ (.A1(_11214_),
    .A2(_13434_),
    .B1(_13435_),
    .Y(_00471_));
 sky130_fd_sc_hd__nor2_1 _21219_ (.A(_10789_),
    .B(_13358_),
    .Y(_13436_));
 sky130_fd_sc_hd__a21oi_1 _21220_ (.A1(net172),
    .A2(_13358_),
    .B1(_13436_),
    .Y(_13437_));
 sky130_fd_sc_hd__nand2_1 _21221_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[30] ),
    .B(_11214_),
    .Y(_13438_));
 sky130_fd_sc_hd__o21ai_0 _21222_ (.A1(_11214_),
    .A2(_13437_),
    .B1(_13438_),
    .Y(_00472_));
 sky130_fd_sc_hd__nand3_4 _21223_ (.A(net564),
    .B(_08262_),
    .C(net600),
    .Y(_13439_));
 sky130_fd_sc_hd__nand4_4 _21224_ (.A(net580),
    .B(_08235_),
    .C(_08216_),
    .D(net527),
    .Y(_13440_));
 sky130_fd_sc_hd__nor2_2 _21225_ (.A(_13439_),
    .B(_13440_),
    .Y(_13441_));
 sky130_fd_sc_hd__nand2_4 _21226_ (.A(_13441_),
    .B(_13357_),
    .Y(_13442_));
 sky130_fd_sc_hd__o21ai_0 _21227_ (.A1(net483),
    .A2(_13442_),
    .B1(_10691_),
    .Y(_13443_));
 sky130_fd_sc_hd__nand2_1 _21228_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ),
    .B(_11214_),
    .Y(_13444_));
 sky130_fd_sc_hd__o21ai_0 _21229_ (.A1(_11214_),
    .A2(_13443_),
    .B1(_13444_),
    .Y(_00473_));
 sky130_fd_sc_hd__nor2_1 _21230_ (.A(net839),
    .B(_13358_),
    .Y(_13445_));
 sky130_fd_sc_hd__a21oi_1 _21231_ (.A1(net174),
    .A2(_13358_),
    .B1(_13445_),
    .Y(_13446_));
 sky130_fd_sc_hd__nand2_1 _21232_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[3] ),
    .B(_11214_),
    .Y(_13447_));
 sky130_fd_sc_hd__o21ai_0 _21233_ (.A1(_11214_),
    .A2(_13446_),
    .B1(_13447_),
    .Y(_00474_));
 sky130_fd_sc_hd__nor2_1 _21234_ (.A(net1459),
    .B(_13358_),
    .Y(_13448_));
 sky130_fd_sc_hd__a21oi_1 _21235_ (.A1(net175),
    .A2(_13358_),
    .B1(_13448_),
    .Y(_13449_));
 sky130_fd_sc_hd__nand2_1 _21236_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[4] ),
    .B(_11214_),
    .Y(_13450_));
 sky130_fd_sc_hd__o21ai_0 _21237_ (.A1(_11214_),
    .A2(_13449_),
    .B1(_13450_),
    .Y(_00475_));
 sky130_fd_sc_hd__nor2_1 _21238_ (.A(net798),
    .B(_13358_),
    .Y(_13451_));
 sky130_fd_sc_hd__a21oi_1 _21239_ (.A1(net1062),
    .A2(_13358_),
    .B1(_13451_),
    .Y(_13452_));
 sky130_fd_sc_hd__nand2_1 _21240_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[5] ),
    .B(_11214_),
    .Y(_13453_));
 sky130_fd_sc_hd__o21ai_0 _21241_ (.A1(_11214_),
    .A2(_13452_),
    .B1(_13453_),
    .Y(_00476_));
 sky130_fd_sc_hd__nor2_1 _21242_ (.A(net574),
    .B(_13358_),
    .Y(_13454_));
 sky130_fd_sc_hd__a21oi_1 _21243_ (.A1(net177),
    .A2(_13358_),
    .B1(_13454_),
    .Y(_13455_));
 sky130_fd_sc_hd__nand2_1 _21244_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[6] ),
    .B(_11214_),
    .Y(_13456_));
 sky130_fd_sc_hd__o21ai_0 _21245_ (.A1(_11214_),
    .A2(_13455_),
    .B1(_13456_),
    .Y(_00477_));
 sky130_fd_sc_hd__nor2_1 _21246_ (.A(net768),
    .B(_13358_),
    .Y(_13457_));
 sky130_fd_sc_hd__a21oi_1 _21247_ (.A1(net178),
    .A2(_13358_),
    .B1(_13457_),
    .Y(_13458_));
 sky130_fd_sc_hd__nand2_1 _21248_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[7] ),
    .B(_11214_),
    .Y(_13459_));
 sky130_fd_sc_hd__o21ai_0 _21249_ (.A1(_11214_),
    .A2(_13458_),
    .B1(_13459_),
    .Y(_00478_));
 sky130_fd_sc_hd__nor2_1 _21250_ (.A(_09184_),
    .B(_13358_),
    .Y(_13460_));
 sky130_fd_sc_hd__a21oi_1 _21251_ (.A1(net179),
    .A2(_13358_),
    .B1(_13460_),
    .Y(_13461_));
 sky130_fd_sc_hd__nand2_1 _21252_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[8] ),
    .B(_11214_),
    .Y(_13462_));
 sky130_fd_sc_hd__o21ai_0 _21253_ (.A1(_11214_),
    .A2(_13461_),
    .B1(_13462_),
    .Y(_00479_));
 sky130_fd_sc_hd__nor2_1 _21254_ (.A(net1121),
    .B(_13358_),
    .Y(_13463_));
 sky130_fd_sc_hd__a21oi_1 _21255_ (.A1(net180),
    .A2(_13358_),
    .B1(_13463_),
    .Y(_13464_));
 sky130_fd_sc_hd__nand2_1 _21256_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[9] ),
    .B(_11214_),
    .Y(_13465_));
 sky130_fd_sc_hd__o21ai_0 _21257_ (.A1(_11214_),
    .A2(_13464_),
    .B1(_13465_),
    .Y(_00480_));
 sky130_fd_sc_hd__clkinv_4 _21258_ (.A(net173),
    .Y(_13466_));
 sky130_fd_sc_hd__a21oi_2 _21259_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[31] ),
    .A2(net481),
    .B1(_10727_),
    .Y(_13467_));
 sky130_fd_sc_hd__a21oi_4 _21260_ (.A1(_10728_),
    .A2(net793),
    .B1(_13467_),
    .Y(_13468_));
 sky130_fd_sc_hd__nor2_4 _21261_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .B(_13468_),
    .Y(_13469_));
 sky130_fd_sc_hd__nor2_4 _21262_ (.A(_10810_),
    .B(_10815_),
    .Y(_13470_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_508 ();
 sky130_fd_sc_hd__nand3_4 _21264_ (.A(_10810_),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .C(_10951_),
    .Y(_13472_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_507 ();
 sky130_fd_sc_hd__a32o_1 _21266_ (.A1(_13350_),
    .A2(_13469_),
    .A3(_13470_),
    .B1(_13472_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[0] ),
    .X(_00481_));
 sky130_fd_sc_hd__nor2b_1 _21267_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .B_N(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .Y(_13474_));
 sky130_fd_sc_hd__nand2_2 _21268_ (.A(_13469_),
    .B(_13474_),
    .Y(_13475_));
 sky130_fd_sc_hd__nand2_2 _21269_ (.A(_13341_),
    .B(_13470_),
    .Y(_13476_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_506 ();
 sky130_fd_sc_hd__nand2_1 _21271_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[10] ),
    .B(_13472_),
    .Y(_13478_));
 sky130_fd_sc_hd__o21ai_0 _21272_ (.A1(_13475_),
    .A2(_13476_),
    .B1(_13478_),
    .Y(_00482_));
 sky130_fd_sc_hd__nand3_4 _21273_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .C(_13470_),
    .Y(_13479_));
 sky130_fd_sc_hd__nand2_1 _21274_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[11] ),
    .B(_13472_),
    .Y(_13480_));
 sky130_fd_sc_hd__o21ai_0 _21275_ (.A1(_13475_),
    .A2(_13479_),
    .B1(_13480_),
    .Y(_00483_));
 sky130_fd_sc_hd__nand3_4 _21276_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .C(_13469_),
    .Y(_13481_));
 sky130_fd_sc_hd__nand2_2 _21277_ (.A(_13344_),
    .B(_13470_),
    .Y(_13482_));
 sky130_fd_sc_hd__nand2_1 _21278_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[12] ),
    .B(_13472_),
    .Y(_13483_));
 sky130_fd_sc_hd__o21ai_0 _21279_ (.A1(_13481_),
    .A2(_13482_),
    .B1(_13483_),
    .Y(_00484_));
 sky130_fd_sc_hd__nand2_2 _21280_ (.A(_10820_),
    .B(_13470_),
    .Y(_13484_));
 sky130_fd_sc_hd__nand2_1 _21281_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[13] ),
    .B(_13472_),
    .Y(_13485_));
 sky130_fd_sc_hd__o21ai_0 _21282_ (.A1(_13481_),
    .A2(_13484_),
    .B1(_13485_),
    .Y(_00485_));
 sky130_fd_sc_hd__nand2_1 _21283_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[14] ),
    .B(_13472_),
    .Y(_13486_));
 sky130_fd_sc_hd__o21ai_0 _21284_ (.A1(_13476_),
    .A2(_13481_),
    .B1(_13486_),
    .Y(_00486_));
 sky130_fd_sc_hd__nand2_1 _21285_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[15] ),
    .B(_13472_),
    .Y(_13487_));
 sky130_fd_sc_hd__o21ai_0 _21286_ (.A1(_13479_),
    .A2(_13481_),
    .B1(_13487_),
    .Y(_00487_));
 sky130_fd_sc_hd__a21o_4 _21287_ (.A1(_10728_),
    .A2(net793),
    .B1(_13467_),
    .X(_13488_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_505 ();
 sky130_fd_sc_hd__and2_4 _21289_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .B(_13488_),
    .X(_13490_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_504 ();
 sky130_fd_sc_hd__a32o_1 _21291_ (.A1(_13350_),
    .A2(_13470_),
    .A3(_13490_),
    .B1(_13472_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[16] ),
    .X(_00488_));
 sky130_fd_sc_hd__nor3_1 _21292_ (.A(_10810_),
    .B(_10815_),
    .C(_10824_),
    .Y(_13492_));
 sky130_fd_sc_hd__a22o_1 _21293_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[17] ),
    .A2(_13472_),
    .B1(_13490_),
    .B2(_13492_),
    .X(_00489_));
 sky130_fd_sc_hd__nand2_1 _21294_ (.A(_10823_),
    .B(_13490_),
    .Y(_13493_));
 sky130_fd_sc_hd__nand2_1 _21295_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[18] ),
    .B(_13472_),
    .Y(_13494_));
 sky130_fd_sc_hd__o21ai_0 _21296_ (.A1(_13476_),
    .A2(_13493_),
    .B1(_13494_),
    .Y(_00490_));
 sky130_fd_sc_hd__nand2_1 _21297_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[19] ),
    .B(_13472_),
    .Y(_13495_));
 sky130_fd_sc_hd__o21ai_0 _21298_ (.A1(_13479_),
    .A2(_13493_),
    .B1(_13495_),
    .Y(_00491_));
 sky130_fd_sc_hd__a22o_1 _21299_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[1] ),
    .A2(_13472_),
    .B1(_13492_),
    .B2(_13469_),
    .X(_00492_));
 sky130_fd_sc_hd__nor2b_1 _21300_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .B_N(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .Y(_13496_));
 sky130_fd_sc_hd__nand2_4 _21301_ (.A(_13490_),
    .B(_13496_),
    .Y(_13497_));
 sky130_fd_sc_hd__nand2_1 _21302_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[20] ),
    .B(_13472_),
    .Y(_13498_));
 sky130_fd_sc_hd__o21ai_0 _21303_ (.A1(_13482_),
    .A2(_13497_),
    .B1(_13498_),
    .Y(_00493_));
 sky130_fd_sc_hd__nand2_1 _21304_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[21] ),
    .B(_13472_),
    .Y(_13499_));
 sky130_fd_sc_hd__o21ai_0 _21305_ (.A1(_13484_),
    .A2(_13497_),
    .B1(_13499_),
    .Y(_00494_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_503 ();
 sky130_fd_sc_hd__nand2_1 _21307_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[22] ),
    .B(_13472_),
    .Y(_13501_));
 sky130_fd_sc_hd__o21ai_0 _21308_ (.A1(_13476_),
    .A2(_13497_),
    .B1(_13501_),
    .Y(_00495_));
 sky130_fd_sc_hd__nand2_1 _21309_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[23] ),
    .B(_13472_),
    .Y(_13502_));
 sky130_fd_sc_hd__o21ai_0 _21310_ (.A1(_13479_),
    .A2(_13497_),
    .B1(_13502_),
    .Y(_00496_));
 sky130_fd_sc_hd__nand2_2 _21311_ (.A(_13474_),
    .B(_13490_),
    .Y(_13503_));
 sky130_fd_sc_hd__nand2_1 _21312_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[24] ),
    .B(_13472_),
    .Y(_01645_));
 sky130_fd_sc_hd__o21ai_0 _21313_ (.A1(_13482_),
    .A2(_13503_),
    .B1(_01645_),
    .Y(_00497_));
 sky130_fd_sc_hd__nand2_1 _21314_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[25] ),
    .B(_13472_),
    .Y(_01646_));
 sky130_fd_sc_hd__o21ai_0 _21315_ (.A1(_13484_),
    .A2(_13503_),
    .B1(_01646_),
    .Y(_00498_));
 sky130_fd_sc_hd__nand2_1 _21316_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[26] ),
    .B(_13472_),
    .Y(_01647_));
 sky130_fd_sc_hd__o21ai_0 _21317_ (.A1(_13476_),
    .A2(_13503_),
    .B1(_01647_),
    .Y(_00499_));
 sky130_fd_sc_hd__nand2_1 _21318_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[27] ),
    .B(_13472_),
    .Y(_01648_));
 sky130_fd_sc_hd__o21ai_0 _21319_ (.A1(_13479_),
    .A2(_13503_),
    .B1(_01648_),
    .Y(_00500_));
 sky130_fd_sc_hd__nand3_4 _21320_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .C(_13490_),
    .Y(_01649_));
 sky130_fd_sc_hd__nand2_1 _21321_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[28] ),
    .B(_13472_),
    .Y(_01650_));
 sky130_fd_sc_hd__o21ai_0 _21322_ (.A1(_13482_),
    .A2(_01649_),
    .B1(_01650_),
    .Y(_00501_));
 sky130_fd_sc_hd__nand2_1 _21323_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[29] ),
    .B(_13472_),
    .Y(_01651_));
 sky130_fd_sc_hd__o21ai_0 _21324_ (.A1(_13484_),
    .A2(_01649_),
    .B1(_01651_),
    .Y(_00502_));
 sky130_fd_sc_hd__nand2_1 _21325_ (.A(_10823_),
    .B(_13469_),
    .Y(_01652_));
 sky130_fd_sc_hd__nand2_1 _21326_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[2] ),
    .B(_13472_),
    .Y(_01653_));
 sky130_fd_sc_hd__o21ai_0 _21327_ (.A1(_13476_),
    .A2(_01652_),
    .B1(_01653_),
    .Y(_00503_));
 sky130_fd_sc_hd__nand2_1 _21328_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[30] ),
    .B(_13472_),
    .Y(_01654_));
 sky130_fd_sc_hd__o21ai_0 _21329_ (.A1(_13476_),
    .A2(_01649_),
    .B1(_01654_),
    .Y(_00504_));
 sky130_fd_sc_hd__nand2_1 _21330_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[31] ),
    .B(_13472_),
    .Y(_01655_));
 sky130_fd_sc_hd__o21ai_0 _21331_ (.A1(_13479_),
    .A2(_01649_),
    .B1(_01655_),
    .Y(_00505_));
 sky130_fd_sc_hd__nand2_1 _21332_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[3] ),
    .B(_13472_),
    .Y(_01656_));
 sky130_fd_sc_hd__o21ai_0 _21333_ (.A1(_13479_),
    .A2(_01652_),
    .B1(_01656_),
    .Y(_00506_));
 sky130_fd_sc_hd__nand2_2 _21334_ (.A(_13469_),
    .B(_13496_),
    .Y(_01657_));
 sky130_fd_sc_hd__nand2_1 _21335_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[4] ),
    .B(_13472_),
    .Y(_01658_));
 sky130_fd_sc_hd__o21ai_0 _21336_ (.A1(_13482_),
    .A2(_01657_),
    .B1(_01658_),
    .Y(_00507_));
 sky130_fd_sc_hd__nand2_1 _21337_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[5] ),
    .B(_13472_),
    .Y(_01659_));
 sky130_fd_sc_hd__o21ai_0 _21338_ (.A1(_13484_),
    .A2(_01657_),
    .B1(_01659_),
    .Y(_00508_));
 sky130_fd_sc_hd__nand2_1 _21339_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[6] ),
    .B(_13472_),
    .Y(_01660_));
 sky130_fd_sc_hd__o21ai_0 _21340_ (.A1(_13476_),
    .A2(_01657_),
    .B1(_01660_),
    .Y(_00509_));
 sky130_fd_sc_hd__nand2_1 _21341_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[7] ),
    .B(_13472_),
    .Y(_01661_));
 sky130_fd_sc_hd__o21ai_0 _21342_ (.A1(_13479_),
    .A2(_01657_),
    .B1(_01661_),
    .Y(_00510_));
 sky130_fd_sc_hd__nand2_1 _21343_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[8] ),
    .B(_13472_),
    .Y(_01662_));
 sky130_fd_sc_hd__o21ai_0 _21344_ (.A1(_13475_),
    .A2(_13482_),
    .B1(_01662_),
    .Y(_00511_));
 sky130_fd_sc_hd__nand2_1 _21345_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ),
    .B(_13472_),
    .Y(_01663_));
 sky130_fd_sc_hd__o21ai_0 _21346_ (.A1(_13475_),
    .A2(_13484_),
    .B1(_01663_),
    .Y(_00512_));
 sky130_fd_sc_hd__or2_0 _21347_ (.A(fetch_enable_q),
    .B(net61),
    .X(_00513_));
 sky130_fd_sc_hd__o311a_1 _21348_ (.A1(net846),
    .A2(_08227_),
    .A3(_08282_),
    .B1(_08446_),
    .C1(_08581_),
    .X(_01664_));
 sky130_fd_sc_hd__nor3_4 _21349_ (.A(_11197_),
    .B(_12128_),
    .C(_01664_),
    .Y(_01665_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_499 ();
 sky130_fd_sc_hd__clkinv_4 _21354_ (.A(\load_store_unit_i.rdata_offset_q[0] ),
    .Y(_01670_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_498 ();
 sky130_fd_sc_hd__nor2_8 _21356_ (.A(_01670_),
    .B(\load_store_unit_i.rdata_offset_q[1] ),
    .Y(_01672_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_497 ();
 sky130_fd_sc_hd__nor2_8 _21358_ (.A(\load_store_unit_i.data_type_q[2] ),
    .B(\load_store_unit_i.data_type_q[1] ),
    .Y(_01674_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_493 ();
 sky130_fd_sc_hd__and3_1 _21363_ (.A(_01670_),
    .B(\load_store_unit_i.rdata_offset_q[1] ),
    .C(net34),
    .X(_01679_));
 sky130_fd_sc_hd__a211oi_2 _21364_ (.A1(net57),
    .A2(_01672_),
    .B1(_01674_),
    .C1(_01679_),
    .Y(_01680_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_492 ();
 sky130_fd_sc_hd__clkinv_4 _21366_ (.A(\load_store_unit_i.rdata_offset_q[1] ),
    .Y(_01682_));
 sky130_fd_sc_hd__nor2_4 _21367_ (.A(\load_store_unit_i.rdata_offset_q[0] ),
    .B(_01682_),
    .Y(_01683_));
 sky130_fd_sc_hd__or2_4 _21368_ (.A(\load_store_unit_i.data_type_q[2] ),
    .B(\load_store_unit_i.data_type_q[1] ),
    .X(_01684_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_490 ();
 sky130_fd_sc_hd__a221oi_2 _21371_ (.A1(\load_store_unit_i.rdata_q[8] ),
    .A2(_01672_),
    .B1(_01683_),
    .B2(\load_store_unit_i.rdata_q[16] ),
    .C1(_01684_),
    .Y(_01687_));
 sky130_fd_sc_hd__nand2b_4 _21372_ (.A_N(\load_store_unit_i.data_type_q[2] ),
    .B(\load_store_unit_i.data_type_q[1] ),
    .Y(_01688_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_489 ();
 sky130_fd_sc_hd__a22oi_2 _21374_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(net43),
    .B1(_01688_),
    .B2(\load_store_unit_i.rdata_q[24] ),
    .Y(_01690_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_487 ();
 sky130_fd_sc_hd__nand2_4 _21377_ (.A(\load_store_unit_i.rdata_offset_q[0] ),
    .B(\load_store_unit_i.rdata_offset_q[1] ),
    .Y(_01693_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_486 ();
 sky130_fd_sc_hd__nand3_1 _21379_ (.A(_01670_),
    .B(_01682_),
    .C(net27),
    .Y(_01695_));
 sky130_fd_sc_hd__o221ai_4 _21380_ (.A1(_01680_),
    .A2(_01687_),
    .B1(_01690_),
    .B2(_01693_),
    .C1(_01695_),
    .Y(_01696_));
 sky130_fd_sc_hd__nand2_2 _21381_ (.A(_11277_),
    .B(net1484),
    .Y(_01697_));
 sky130_fd_sc_hd__nor3_4 _21382_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .C(net316),
    .Y(_01698_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_485 ();
 sky130_fd_sc_hd__nor2_4 _21384_ (.A(_13335_),
    .B(_01698_),
    .Y(_01700_));
 sky130_fd_sc_hd__mux2i_1 _21385_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[48] ),
    .A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[32] ),
    .S(net316),
    .Y(_01701_));
 sky130_fd_sc_hd__or2_4 _21386_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .X(_01702_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_479 ();
 sky130_fd_sc_hd__nand2_1 _21393_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[48] ),
    .B(net322),
    .Y(_01709_));
 sky130_fd_sc_hd__o21ai_2 _21394_ (.A1(_08280_),
    .A2(_01701_),
    .B1(_01709_),
    .Y(_01710_));
 sky130_fd_sc_hd__nand4_4 _21395_ (.A(_09834_),
    .B(_09848_),
    .C(_09841_),
    .D(_09855_),
    .Y(_01711_));
 sky130_fd_sc_hd__nor2_8 _21396_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .Y(_01712_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_477 ();
 sky130_fd_sc_hd__nand2_2 _21399_ (.A(_08916_),
    .B(net320),
    .Y(_01715_));
 sky130_fd_sc_hd__nand3_4 _21400_ (.A(_08926_),
    .B(_08947_),
    .C(_08940_),
    .Y(_01716_));
 sky130_fd_sc_hd__o22ai_4 _21401_ (.A1(net320),
    .A2(_01711_),
    .B1(_01715_),
    .B2(_01716_),
    .Y(_01717_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_476 ();
 sky130_fd_sc_hd__and3_2 _21403_ (.A(_09799_),
    .B(_09813_),
    .C(_09820_),
    .X(_01719_));
 sky130_fd_sc_hd__or2_4 _21404_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .X(_01720_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_473 ();
 sky130_fd_sc_hd__nor4_4 _21408_ (.A(_08873_),
    .B(_08886_),
    .C(_08894_),
    .D(_01720_),
    .Y(_01724_));
 sky130_fd_sc_hd__a21oi_4 _21409_ (.A1(_01719_),
    .A2(_01720_),
    .B1(_01724_),
    .Y(_01725_));
 sky130_fd_sc_hd__nor2_1 _21410_ (.A(net945),
    .B(net1279),
    .Y(_01726_));
 sky130_fd_sc_hd__xnor2_1 _21411_ (.A(_01710_),
    .B(_01726_),
    .Y(_01727_));
 sky130_fd_sc_hd__nand2_1 _21412_ (.A(_01700_),
    .B(_01727_),
    .Y(_01728_));
 sky130_fd_sc_hd__o21ai_2 _21413_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[32] ),
    .A2(_01700_),
    .B1(_01728_),
    .Y(_01729_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_472 ();
 sky130_fd_sc_hd__a21oi_1 _21415_ (.A1(_08272_),
    .A2(_01729_),
    .B1(_08632_),
    .Y(_01731_));
 sky130_fd_sc_hd__o22ai_4 _21416_ (.A1(net265),
    .A2(_01696_),
    .B1(_01697_),
    .B2(_01731_),
    .Y(_01732_));
 sky130_fd_sc_hd__nor2_8 _21417_ (.A(net1461),
    .B(_11171_),
    .Y(_01733_));
 sky130_fd_sc_hd__nor2_8 _21418_ (.A(_08382_),
    .B(_08428_),
    .Y(_01734_));
 sky130_fd_sc_hd__and3_2 _21419_ (.A(_10695_),
    .B(_11175_),
    .C(_01734_),
    .X(_01735_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_471 ();
 sky130_fd_sc_hd__a21oi_4 _21421_ (.A1(net711),
    .A2(_10891_),
    .B1(_08381_),
    .Y(_01737_));
 sky130_fd_sc_hd__xnor2_4 _21422_ (.A(net1131),
    .B(_01737_),
    .Y(_01738_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_468 ();
 sky130_fd_sc_hd__nor2_4 _21426_ (.A(_08381_),
    .B(_10895_),
    .Y(_01742_));
 sky130_fd_sc_hd__xnor2_4 _21427_ (.A(_11246_),
    .B(_01742_),
    .Y(_01743_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_466 ();
 sky130_fd_sc_hd__nand2_2 _21430_ (.A(_01738_),
    .B(_01743_),
    .Y(_01746_));
 sky130_fd_sc_hd__nand2_4 _21431_ (.A(_08362_),
    .B(_10894_),
    .Y(_01747_));
 sky130_fd_sc_hd__xor2_4 _21432_ (.A(net709),
    .B(_01747_),
    .X(_01748_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_465 ();
 sky130_fd_sc_hd__nand2_4 _21434_ (.A(_08362_),
    .B(net643),
    .Y(_01750_));
 sky130_fd_sc_hd__xnor2_4 _21435_ (.A(net729),
    .B(_01750_),
    .Y(_01751_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 ();
 sky130_fd_sc_hd__and2_1 _21439_ (.A(_11175_),
    .B(_01734_),
    .X(_01755_));
 sky130_fd_sc_hd__nand2_4 _21440_ (.A(_10695_),
    .B(_01755_),
    .Y(_01756_));
 sky130_fd_sc_hd__o21ai_0 _21441_ (.A1(_01748_),
    .A2(_01751_),
    .B1(_01756_),
    .Y(_01757_));
 sky130_fd_sc_hd__xnor2_4 _21442_ (.A(net710),
    .B(_01747_),
    .Y(_01758_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 ();
 sky130_fd_sc_hd__nand2b_4 _21445_ (.A_N(_08428_),
    .B(_08410_),
    .Y(_01761_));
 sky130_fd_sc_hd__nor3_4 _21446_ (.A(net1463),
    .B(_11171_),
    .C(_01761_),
    .Y(_01762_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_459 ();
 sky130_fd_sc_hd__nor2_1 _21448_ (.A(_10695_),
    .B(_01762_),
    .Y(_01764_));
 sky130_fd_sc_hd__a21oi_1 _21449_ (.A1(_08897_),
    .A2(_01762_),
    .B1(_01764_),
    .Y(_01765_));
 sky130_fd_sc_hd__o21ai_2 _21450_ (.A1(_10902_),
    .A2(_01755_),
    .B1(_01765_),
    .Y(_01766_));
 sky130_fd_sc_hd__nand2_1 _21451_ (.A(_01758_),
    .B(_01766_),
    .Y(_01767_));
 sky130_fd_sc_hd__nand2_1 _21452_ (.A(_01757_),
    .B(_01767_),
    .Y(_01768_));
 sky130_fd_sc_hd__nor2_1 _21453_ (.A(_01768_),
    .B(_01746_),
    .Y(_01769_));
 sky130_fd_sc_hd__a21oi_1 _21454_ (.A1(_01735_),
    .A2(_01746_),
    .B1(_01769_),
    .Y(_01770_));
 sky130_fd_sc_hd__xor2_4 _21455_ (.A(net730),
    .B(_01750_),
    .X(_01771_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_458 ();
 sky130_fd_sc_hd__nand2_8 _21457_ (.A(_01733_),
    .B(_01734_),
    .Y(_01773_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_457 ();
 sky130_fd_sc_hd__mux2i_1 _21459_ (.A0(net954),
    .A1(_10468_),
    .S(_01773_),
    .Y(_01775_));
 sky130_fd_sc_hd__nor2_1 _21460_ (.A(_10497_),
    .B(net295),
    .Y(_01776_));
 sky130_fd_sc_hd__a21oi_1 _21461_ (.A1(_08585_),
    .A2(net294),
    .B1(_01776_),
    .Y(_01777_));
 sky130_fd_sc_hd__nand2_1 _21462_ (.A(net300),
    .B(_01777_),
    .Y(_01778_));
 sky130_fd_sc_hd__o21ai_0 _21463_ (.A1(net300),
    .A2(_01775_),
    .B1(_01778_),
    .Y(_01779_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_456 ();
 sky130_fd_sc_hd__mux2i_1 _21465_ (.A0(_08375_),
    .A1(_10368_),
    .S(_01773_),
    .Y(_01781_));
 sky130_fd_sc_hd__nor2_1 _21466_ (.A(net300),
    .B(_01781_),
    .Y(_01782_));
 sky130_fd_sc_hd__nand2_1 _21467_ (.A(_10303_),
    .B(_01773_),
    .Y(_01783_));
 sky130_fd_sc_hd__o21ai_0 _21468_ (.A1(_08547_),
    .A2(_01773_),
    .B1(_01783_),
    .Y(_01784_));
 sky130_fd_sc_hd__nor2_1 _21469_ (.A(net1466),
    .B(_01784_),
    .Y(_01785_));
 sky130_fd_sc_hd__nor2_1 _21470_ (.A(_01782_),
    .B(_01785_),
    .Y(_01786_));
 sky130_fd_sc_hd__nand2_1 _21471_ (.A(_01771_),
    .B(_01786_),
    .Y(_01787_));
 sky130_fd_sc_hd__o21ai_1 _21472_ (.A1(_01771_),
    .A2(_01779_),
    .B1(_01787_),
    .Y(_01788_));
 sky130_fd_sc_hd__nor2_1 _21473_ (.A(_10655_),
    .B(net295),
    .Y(_01789_));
 sky130_fd_sc_hd__a21oi_1 _21474_ (.A1(_08636_),
    .A2(net294),
    .B1(_01789_),
    .Y(_01790_));
 sky130_fd_sc_hd__nand2_1 _21475_ (.A(_08850_),
    .B(net295),
    .Y(_01791_));
 sky130_fd_sc_hd__o21ai_0 _21476_ (.A1(_10561_),
    .A2(net295),
    .B1(_01791_),
    .Y(_01792_));
 sky130_fd_sc_hd__nor2_1 _21477_ (.A(net1466),
    .B(_01792_),
    .Y(_01793_));
 sky130_fd_sc_hd__a21oi_1 _21478_ (.A1(net1466),
    .A2(_01790_),
    .B1(_01793_),
    .Y(_01794_));
 sky130_fd_sc_hd__nand2_1 _21479_ (.A(_09044_),
    .B(net295),
    .Y(_01795_));
 sky130_fd_sc_hd__o21ai_0 _21480_ (.A1(_10799_),
    .A2(net295),
    .B1(_01795_),
    .Y(_01796_));
 sky130_fd_sc_hd__nand2_1 _21481_ (.A(net637),
    .B(_01765_),
    .Y(_01797_));
 sky130_fd_sc_hd__o21ai_0 _21482_ (.A1(net638),
    .A2(_01796_),
    .B1(_01797_),
    .Y(_01798_));
 sky130_fd_sc_hd__nor2_1 _21483_ (.A(_01771_),
    .B(_01798_),
    .Y(_01799_));
 sky130_fd_sc_hd__a21oi_1 _21484_ (.A1(_01771_),
    .A2(_01794_),
    .B1(_01799_),
    .Y(_01800_));
 sky130_fd_sc_hd__nand2_1 _21485_ (.A(_01748_),
    .B(_01800_),
    .Y(_01801_));
 sky130_fd_sc_hd__o21ai_1 _21486_ (.A1(_01748_),
    .A2(_01788_),
    .B1(_01801_),
    .Y(_01802_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_454 ();
 sky130_fd_sc_hd__mux2i_1 _21489_ (.A0(_09679_),
    .A1(_09825_),
    .S(_01773_),
    .Y(_01805_));
 sky130_fd_sc_hd__nor2_1 _21490_ (.A(_09640_),
    .B(_01773_),
    .Y(_01806_));
 sky130_fd_sc_hd__a21oi_1 _21491_ (.A1(_09754_),
    .A2(_01773_),
    .B1(_01806_),
    .Y(_01807_));
 sky130_fd_sc_hd__nand2_1 _21492_ (.A(net299),
    .B(_01807_),
    .Y(_01808_));
 sky130_fd_sc_hd__o21ai_1 _21493_ (.A1(net299),
    .A2(_01805_),
    .B1(_01808_),
    .Y(_01809_));
 sky130_fd_sc_hd__mux2i_1 _21494_ (.A0(_09450_),
    .A1(_09898_),
    .S(_01773_),
    .Y(_01810_));
 sky130_fd_sc_hd__mux2i_4 _21495_ (.A0(_09562_),
    .A1(_10008_),
    .S(_01773_),
    .Y(_01811_));
 sky130_fd_sc_hd__mux2i_2 _21496_ (.A0(_01810_),
    .A1(_01811_),
    .S(net299),
    .Y(_01812_));
 sky130_fd_sc_hd__mux2i_2 _21497_ (.A0(_01809_),
    .A1(_01812_),
    .S(_01751_),
    .Y(_01813_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_453 ();
 sky130_fd_sc_hd__nand2_1 _21499_ (.A(net879),
    .B(net294),
    .Y(_01815_));
 sky130_fd_sc_hd__o21ai_2 _21500_ (.A1(_10070_),
    .A2(net294),
    .B1(_01815_),
    .Y(_01816_));
 sky130_fd_sc_hd__mux2i_4 _21501_ (.A0(_09385_),
    .A1(_10145_),
    .S(_01773_),
    .Y(_01817_));
 sky130_fd_sc_hd__mux2i_2 _21502_ (.A0(_01816_),
    .A1(_01817_),
    .S(net299),
    .Y(_01818_));
 sky130_fd_sc_hd__mux2i_4 _21503_ (.A0(_09290_),
    .A1(_10172_),
    .S(_01773_),
    .Y(_01819_));
 sky130_fd_sc_hd__nand2_1 _21504_ (.A(_10272_),
    .B(_01773_),
    .Y(_01820_));
 sky130_fd_sc_hd__o21ai_1 _21505_ (.A1(_09187_),
    .A2(_01773_),
    .B1(_01820_),
    .Y(_01821_));
 sky130_fd_sc_hd__mux2i_2 _21506_ (.A0(_01819_),
    .A1(_01821_),
    .S(net299),
    .Y(_01822_));
 sky130_fd_sc_hd__mux2i_2 _21507_ (.A0(_01818_),
    .A1(_01822_),
    .S(_01751_),
    .Y(_01823_));
 sky130_fd_sc_hd__mux2i_2 _21508_ (.A0(_01813_),
    .A1(_01823_),
    .S(_01748_),
    .Y(_01824_));
 sky130_fd_sc_hd__mux2i_1 _21509_ (.A0(_01802_),
    .A1(_01824_),
    .S(_01738_),
    .Y(_01825_));
 sky130_fd_sc_hd__xor2_4 _21510_ (.A(net1132),
    .B(_01737_),
    .X(_01826_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 ();
 sky130_fd_sc_hd__mux2i_2 _21514_ (.A0(net954),
    .A1(_10468_),
    .S(net294),
    .Y(_01830_));
 sky130_fd_sc_hd__nand2_1 _21515_ (.A(_10497_),
    .B(net294),
    .Y(_01831_));
 sky130_fd_sc_hd__o21ai_0 _21516_ (.A1(_08585_),
    .A2(net294),
    .B1(_01831_),
    .Y(_01832_));
 sky130_fd_sc_hd__nand2_1 _21517_ (.A(net1468),
    .B(_01832_),
    .Y(_01833_));
 sky130_fd_sc_hd__o21ai_1 _21518_ (.A1(net1468),
    .A2(_01830_),
    .B1(_01833_),
    .Y(_01834_));
 sky130_fd_sc_hd__nor2_1 _21519_ (.A(_01751_),
    .B(_01834_),
    .Y(_01835_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 ();
 sky130_fd_sc_hd__nand2_1 _21521_ (.A(_10303_),
    .B(net294),
    .Y(_01837_));
 sky130_fd_sc_hd__o21ai_1 _21522_ (.A1(_08547_),
    .A2(net294),
    .B1(_01837_),
    .Y(_01838_));
 sky130_fd_sc_hd__nor2_1 _21523_ (.A(_10368_),
    .B(_01773_),
    .Y(_01839_));
 sky130_fd_sc_hd__nor2_1 _21524_ (.A(_08375_),
    .B(net294),
    .Y(_01840_));
 sky130_fd_sc_hd__nor2_1 _21525_ (.A(_01839_),
    .B(_01840_),
    .Y(_01841_));
 sky130_fd_sc_hd__nand2_1 _21526_ (.A(net300),
    .B(_01841_),
    .Y(_01842_));
 sky130_fd_sc_hd__o21ai_0 _21527_ (.A1(net300),
    .A2(_01838_),
    .B1(_01842_),
    .Y(_01843_));
 sky130_fd_sc_hd__nor2_1 _21528_ (.A(_01771_),
    .B(_01843_),
    .Y(_01844_));
 sky130_fd_sc_hd__nor3_1 _21529_ (.A(_01758_),
    .B(_01835_),
    .C(_01844_),
    .Y(_01845_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 ();
 sky130_fd_sc_hd__nor2_1 _21531_ (.A(_10799_),
    .B(_01773_),
    .Y(_01847_));
 sky130_fd_sc_hd__a21oi_1 _21532_ (.A1(_09044_),
    .A2(_01773_),
    .B1(_01847_),
    .Y(_01848_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 ();
 sky130_fd_sc_hd__nor2_1 _21534_ (.A(_10695_),
    .B(_01773_),
    .Y(_01850_));
 sky130_fd_sc_hd__a211oi_1 _21535_ (.A1(net731),
    .A2(_01773_),
    .B1(_01850_),
    .C1(net300),
    .Y(_01851_));
 sky130_fd_sc_hd__a211oi_1 _21536_ (.A1(net300),
    .A2(_01848_),
    .B1(_01851_),
    .C1(_01751_),
    .Y(_01852_));
 sky130_fd_sc_hd__nand2_1 _21537_ (.A(_08850_),
    .B(_01773_),
    .Y(_01853_));
 sky130_fd_sc_hd__o21ai_1 _21538_ (.A1(_10561_),
    .A2(_01773_),
    .B1(_01853_),
    .Y(_01854_));
 sky130_fd_sc_hd__nand2_1 _21539_ (.A(_08636_),
    .B(_01773_),
    .Y(_01855_));
 sky130_fd_sc_hd__o21ai_1 _21540_ (.A1(_10655_),
    .A2(_01773_),
    .B1(_01855_),
    .Y(_01856_));
 sky130_fd_sc_hd__mux2i_2 _21541_ (.A0(_01854_),
    .A1(_01856_),
    .S(net300),
    .Y(_01857_));
 sky130_fd_sc_hd__nor2_1 _21542_ (.A(_01771_),
    .B(_01857_),
    .Y(_01858_));
 sky130_fd_sc_hd__nor3_1 _21543_ (.A(_01748_),
    .B(_01852_),
    .C(_01858_),
    .Y(_01859_));
 sky130_fd_sc_hd__nand2_1 _21544_ (.A(_10272_),
    .B(net294),
    .Y(_01860_));
 sky130_fd_sc_hd__o21ai_1 _21545_ (.A1(_09187_),
    .A2(net294),
    .B1(_01860_),
    .Y(_01861_));
 sky130_fd_sc_hd__mux2i_2 _21546_ (.A0(_09290_),
    .A1(_10172_),
    .S(net294),
    .Y(_01862_));
 sky130_fd_sc_hd__mux2i_2 _21547_ (.A0(_01861_),
    .A1(_01862_),
    .S(net300),
    .Y(_01863_));
 sky130_fd_sc_hd__mux2i_2 _21548_ (.A0(_09385_),
    .A1(_10145_),
    .S(net294),
    .Y(_01864_));
 sky130_fd_sc_hd__nand2_1 _21549_ (.A(net879),
    .B(_01773_),
    .Y(_01865_));
 sky130_fd_sc_hd__o21ai_2 _21550_ (.A1(_10070_),
    .A2(_01773_),
    .B1(_01865_),
    .Y(_01866_));
 sky130_fd_sc_hd__mux2i_2 _21551_ (.A0(_01864_),
    .A1(_01866_),
    .S(net300),
    .Y(_01867_));
 sky130_fd_sc_hd__mux2i_2 _21552_ (.A0(_01863_),
    .A1(_01867_),
    .S(_01751_),
    .Y(_01868_));
 sky130_fd_sc_hd__mux2i_4 _21553_ (.A0(_09562_),
    .A1(_10008_),
    .S(net294),
    .Y(_01869_));
 sky130_fd_sc_hd__mux2i_4 _21554_ (.A0(net738),
    .A1(_09898_),
    .S(net294),
    .Y(_01870_));
 sky130_fd_sc_hd__mux2i_4 _21555_ (.A0(_01869_),
    .A1(_01870_),
    .S(net299),
    .Y(_01871_));
 sky130_fd_sc_hd__mux2i_1 _21556_ (.A0(_09679_),
    .A1(_09825_),
    .S(net294),
    .Y(_01872_));
 sky130_fd_sc_hd__nor2_1 _21557_ (.A(_09640_),
    .B(net294),
    .Y(_01873_));
 sky130_fd_sc_hd__a21oi_1 _21558_ (.A1(_09754_),
    .A2(net294),
    .B1(_01873_),
    .Y(_01874_));
 sky130_fd_sc_hd__nor2_1 _21559_ (.A(net299),
    .B(_01874_),
    .Y(_01875_));
 sky130_fd_sc_hd__a21oi_2 _21560_ (.A1(net299),
    .A2(_01872_),
    .B1(_01875_),
    .Y(_01876_));
 sky130_fd_sc_hd__mux2i_4 _21561_ (.A0(_01871_),
    .A1(_01876_),
    .S(_01751_),
    .Y(_01877_));
 sky130_fd_sc_hd__mux2i_4 _21562_ (.A0(_01868_),
    .A1(_01877_),
    .S(_01748_),
    .Y(_01878_));
 sky130_fd_sc_hd__or2_0 _21563_ (.A(_01738_),
    .B(_01878_),
    .X(_01879_));
 sky130_fd_sc_hd__o31ai_2 _21564_ (.A1(_01826_),
    .A2(_01845_),
    .A3(_01859_),
    .B1(_01879_),
    .Y(_01880_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 ();
 sky130_fd_sc_hd__mux2i_2 _21566_ (.A0(_01825_),
    .A1(_01880_),
    .S(_01743_),
    .Y(_01882_));
 sky130_fd_sc_hd__nor2_1 _21567_ (.A(_01733_),
    .B(_01882_),
    .Y(_01883_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_444 ();
 sky130_fd_sc_hd__a211oi_2 _21570_ (.A1(_01733_),
    .A2(_01770_),
    .B1(_01883_),
    .C1(_01761_),
    .Y(_01886_));
 sky130_fd_sc_hd__nand2_1 _21571_ (.A(_08414_),
    .B(_08428_),
    .Y(_01887_));
 sky130_fd_sc_hd__inv_2 _21572_ (.A(_01887_),
    .Y(_01888_));
 sky130_fd_sc_hd__nand2_8 _21573_ (.A(net1048),
    .B(_01888_),
    .Y(_01889_));
 sky130_fd_sc_hd__nor2_2 _21574_ (.A(_08429_),
    .B(_11171_),
    .Y(_01890_));
 sky130_fd_sc_hd__nand2_1 _21575_ (.A(net1462),
    .B(_01888_),
    .Y(_01891_));
 sky130_fd_sc_hd__o21ai_2 _21576_ (.A1(net646),
    .A2(net1463),
    .B1(_01891_),
    .Y(_01892_));
 sky130_fd_sc_hd__and2_4 _21577_ (.A(_01890_),
    .B(_01892_),
    .X(_01893_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_442 ();
 sky130_fd_sc_hd__nand2_8 _21580_ (.A(_01888_),
    .B(_01733_),
    .Y(_01896_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_441 ();
 sky130_fd_sc_hd__nor2_8 _21582_ (.A(_08429_),
    .B(net645),
    .Y(_01898_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_440 ();
 sky130_fd_sc_hd__nor3_1 _21584_ (.A(_08897_),
    .B(_10902_),
    .C(_01898_),
    .Y(_01900_));
 sky130_fd_sc_hd__a21oi_1 _21585_ (.A1(_08897_),
    .A2(_01896_),
    .B1(_01900_),
    .Y(_01901_));
 sky130_fd_sc_hd__nor3_4 _21586_ (.A(_08424_),
    .B(_01887_),
    .C(_11171_),
    .Y(_01902_));
 sky130_fd_sc_hd__nor2_4 _21587_ (.A(_01893_),
    .B(_01902_),
    .Y(_01903_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_439 ();
 sky130_fd_sc_hd__o21ai_0 _21589_ (.A1(_08897_),
    .A2(_01903_),
    .B1(_10902_),
    .Y(_01905_));
 sky130_fd_sc_hd__o21ai_1 _21590_ (.A1(_01893_),
    .A2(_01901_),
    .B1(_01905_),
    .Y(_01906_));
 sky130_fd_sc_hd__o211ai_4 _21591_ (.A1(_10967_),
    .A2(_01889_),
    .B1(_01906_),
    .C1(_08290_),
    .Y(_01907_));
 sky130_fd_sc_hd__a2111oi_4 _21592_ (.A1(_08429_),
    .A2(_11192_),
    .B1(_01697_),
    .C1(_01886_),
    .D1(_01907_),
    .Y(_01908_));
 sky130_fd_sc_hd__nor2_8 _21593_ (.A(_01732_),
    .B(_01908_),
    .Y(_01909_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_438 ();
 sky130_fd_sc_hd__nor4_2 _21595_ (.A(\load_store_unit_i.data_we_q ),
    .B(net25),
    .C(\load_store_unit_i.lsu_err_q ),
    .D(_10849_),
    .Y(_01911_));
 sky130_fd_sc_hd__nor2_4 _21596_ (.A(net267),
    .B(_01911_),
    .Y(_01912_));
 sky130_fd_sc_hd__or4_4 _21597_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .B(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .C(net448),
    .D(_01912_),
    .X(_01913_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 ();
 sky130_fd_sc_hd__nand2b_4 _21599_ (.A_N(net1021),
    .B(net331),
    .Y(_01915_));
 sky130_fd_sc_hd__nor2_8 _21600_ (.A(_01913_),
    .B(_01915_),
    .Y(_01916_));
 sky130_fd_sc_hd__nand2_1 _21601_ (.A(_01909_),
    .B(_01916_),
    .Y(_01917_));
 sky130_fd_sc_hd__nor4_4 _21602_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .B(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .C(net447),
    .D(_01912_),
    .Y(_01918_));
 sky130_fd_sc_hd__nor2b_4 _21603_ (.A(net1020),
    .B_N(net331),
    .Y(_01919_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 ();
 sky130_fd_sc_hd__nand2_8 _21605_ (.A(_01918_),
    .B(_01919_),
    .Y(_01921_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 ();
 sky130_fd_sc_hd__nand2_1 _21607_ (.A(\gen_regfile_ff.register_file_i.rf_reg[32] ),
    .B(_01921_),
    .Y(_01923_));
 sky130_fd_sc_hd__nand2_1 _21608_ (.A(_01917_),
    .B(_01923_),
    .Y(_00514_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_434 ();
 sky130_fd_sc_hd__nor3_1 _21610_ (.A(_08585_),
    .B(net974),
    .C(_01898_),
    .Y(_01925_));
 sky130_fd_sc_hd__a21oi_1 _21611_ (.A1(_08585_),
    .A2(_01896_),
    .B1(_01925_),
    .Y(_01926_));
 sky130_fd_sc_hd__o21ai_0 _21612_ (.A1(_08585_),
    .A2(_01903_),
    .B1(net974),
    .Y(_01927_));
 sky130_fd_sc_hd__o21ai_0 _21613_ (.A1(_01893_),
    .A2(_01926_),
    .B1(_01927_),
    .Y(_01928_));
 sky130_fd_sc_hd__and3_4 _21614_ (.A(net1048),
    .B(_08414_),
    .C(_08428_),
    .X(_01929_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_429 ();
 sky130_fd_sc_hd__mux2i_1 _21620_ (.A0(_01777_),
    .A1(_01790_),
    .S(net300),
    .Y(_01935_));
 sky130_fd_sc_hd__mux2i_1 _21621_ (.A0(_01792_),
    .A1(_01796_),
    .S(net638),
    .Y(_01936_));
 sky130_fd_sc_hd__nor2_1 _21622_ (.A(_01771_),
    .B(_01936_),
    .Y(_01937_));
 sky130_fd_sc_hd__a21oi_1 _21623_ (.A1(_01771_),
    .A2(_01935_),
    .B1(_01937_),
    .Y(_01938_));
 sky130_fd_sc_hd__a211oi_1 _21624_ (.A1(_01756_),
    .A2(_01751_),
    .B1(_01766_),
    .C1(_01758_),
    .Y(_01939_));
 sky130_fd_sc_hd__a21oi_1 _21625_ (.A1(_01758_),
    .A2(_01938_),
    .B1(_01939_),
    .Y(_01940_));
 sky130_fd_sc_hd__nor2_1 _21626_ (.A(_01735_),
    .B(_01738_),
    .Y(_01941_));
 sky130_fd_sc_hd__a21oi_1 _21627_ (.A1(_01738_),
    .A2(_01940_),
    .B1(_01941_),
    .Y(_01942_));
 sky130_fd_sc_hd__nor2_2 _21628_ (.A(_01756_),
    .B(_01743_),
    .Y(_01943_));
 sky130_fd_sc_hd__a21oi_1 _21629_ (.A1(_01743_),
    .A2(_01942_),
    .B1(_01943_),
    .Y(_01944_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_428 ();
 sky130_fd_sc_hd__mux2i_2 _21631_ (.A0(_01788_),
    .A1(_01823_),
    .S(_01758_),
    .Y(_01946_));
 sky130_fd_sc_hd__nor2_1 _21632_ (.A(_01756_),
    .B(_01758_),
    .Y(_01947_));
 sky130_fd_sc_hd__a21oi_1 _21633_ (.A1(_01758_),
    .A2(_01800_),
    .B1(_01947_),
    .Y(_01948_));
 sky130_fd_sc_hd__nand2_1 _21634_ (.A(_01826_),
    .B(_01948_),
    .Y(_01949_));
 sky130_fd_sc_hd__o21ai_1 _21635_ (.A1(_01826_),
    .A2(_01946_),
    .B1(_01949_),
    .Y(_01950_));
 sky130_fd_sc_hd__mux2i_1 _21636_ (.A0(_01813_),
    .A1(_01877_),
    .S(_01758_),
    .Y(_01951_));
 sky130_fd_sc_hd__or3_1 _21637_ (.A(_01748_),
    .B(_01835_),
    .C(_01844_),
    .X(_01952_));
 sky130_fd_sc_hd__o211ai_1 _21638_ (.A1(_01758_),
    .A2(_01868_),
    .B1(_01952_),
    .C1(_01738_),
    .Y(_01953_));
 sky130_fd_sc_hd__o211ai_1 _21639_ (.A1(_01738_),
    .A2(_01951_),
    .B1(_01953_),
    .C1(_01743_),
    .Y(_01954_));
 sky130_fd_sc_hd__o21ai_1 _21640_ (.A1(_01743_),
    .A2(_01950_),
    .B1(_01954_),
    .Y(_01955_));
 sky130_fd_sc_hd__nor2_1 _21641_ (.A(_01762_),
    .B(_01955_),
    .Y(_01956_));
 sky130_fd_sc_hd__a211oi_2 _21642_ (.A1(_01762_),
    .A2(_01944_),
    .B1(_01956_),
    .C1(_01761_),
    .Y(_01957_));
 sky130_fd_sc_hd__a21oi_1 _21643_ (.A1(net175),
    .A2(_01929_),
    .B1(_01957_),
    .Y(_01958_));
 sky130_fd_sc_hd__nand3_1 _21644_ (.A(net739),
    .B(_01928_),
    .C(_01958_),
    .Y(_01959_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_425 ();
 sky130_fd_sc_hd__mux2i_1 _21648_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[50] ),
    .A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[34] ),
    .S(net316),
    .Y(_01963_));
 sky130_fd_sc_hd__nand2_1 _21649_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[50] ),
    .B(_01702_),
    .Y(_01964_));
 sky130_fd_sc_hd__o21ai_1 _21650_ (.A1(_08280_),
    .A2(_01963_),
    .B1(_01964_),
    .Y(_01965_));
 sky130_fd_sc_hd__or4_4 _21651_ (.A(_08810_),
    .B(_08824_),
    .C(_08838_),
    .D(_01720_),
    .X(_01966_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_424 ();
 sky130_fd_sc_hd__nor2_8 _21653_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .Y(_01968_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_423 ();
 sky130_fd_sc_hd__or4_4 _21655_ (.A(_09894_),
    .B(_09884_),
    .C(_09878_),
    .D(_01968_),
    .X(_01970_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_422 ();
 sky130_fd_sc_hd__and2_4 _21657_ (.A(_01966_),
    .B(_01970_),
    .X(_01972_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_420 ();
 sky130_fd_sc_hd__nor2_4 _21660_ (.A(net945),
    .B(_01972_),
    .Y(_01975_));
 sky130_fd_sc_hd__o2111a_4 _21661_ (.A1(_09010_),
    .A2(_09018_),
    .B1(_01968_),
    .C1(_09034_),
    .D1(_09025_),
    .X(_01976_));
 sky130_fd_sc_hd__o2111a_4 _21662_ (.A1(_09729_),
    .A2(_09735_),
    .B1(_01720_),
    .C1(_09750_),
    .D1(_09742_),
    .X(_01977_));
 sky130_fd_sc_hd__or2_4 _21663_ (.A(_01976_),
    .B(_01977_),
    .X(_01978_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_419 ();
 sky130_fd_sc_hd__and4b_4 _21665_ (.A_N(_09763_),
    .B(net1304),
    .C(_09783_),
    .D(net321),
    .X(_01980_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_418 ();
 sky130_fd_sc_hd__a21o_4 _21667_ (.A1(net658),
    .A2(_01712_),
    .B1(_01980_),
    .X(_01982_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_417 ();
 sky130_fd_sc_hd__nor2_8 _21669_ (.A(_01982_),
    .B(net1224),
    .Y(_01984_));
 sky130_fd_sc_hd__maj3_2 _21670_ (.A(_01965_),
    .B(_01975_),
    .C(_01984_),
    .X(_01985_));
 sky130_fd_sc_hd__mux2i_1 _21671_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[51] ),
    .A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[35] ),
    .S(net315),
    .Y(_01986_));
 sky130_fd_sc_hd__nand2_1 _21672_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[51] ),
    .B(net322),
    .Y(_01987_));
 sky130_fd_sc_hd__o21a_1 _21673_ (.A1(_08280_),
    .A2(_01986_),
    .B1(_01987_),
    .X(_01988_));
 sky130_fd_sc_hd__nor2_4 _21674_ (.A(_01972_),
    .B(_01982_),
    .Y(_01989_));
 sky130_fd_sc_hd__nor3_4 _21675_ (.A(_08629_),
    .B(_08617_),
    .C(_01720_),
    .Y(_01990_));
 sky130_fd_sc_hd__and4_4 _21676_ (.A(_09951_),
    .B(_09955_),
    .C(_09968_),
    .D(_01720_),
    .X(_01991_));
 sky130_fd_sc_hd__nor2_8 _21677_ (.A(_01990_),
    .B(_01991_),
    .Y(_01992_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_416 ();
 sky130_fd_sc_hd__nor2_1 _21679_ (.A(_01717_),
    .B(_01992_),
    .Y(_01994_));
 sky130_fd_sc_hd__xnor3_2 _21680_ (.A(_01988_),
    .B(_01989_),
    .C(_01994_),
    .X(_01995_));
 sky130_fd_sc_hd__or4_4 _21681_ (.A(_08873_),
    .B(_08886_),
    .C(_08894_),
    .D(_01720_),
    .X(_01996_));
 sky130_fd_sc_hd__nand4_4 _21682_ (.A(_09799_),
    .B(_09813_),
    .C(_09820_),
    .D(_01720_),
    .Y(_01997_));
 sky130_fd_sc_hd__nand2_8 _21683_ (.A(_01996_),
    .B(_01997_),
    .Y(_01998_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_413 ();
 sky130_fd_sc_hd__o211ai_2 _21687_ (.A1(_08679_),
    .A2(_08685_),
    .B1(_08691_),
    .C1(net320),
    .Y(_02002_));
 sky130_fd_sc_hd__a31oi_4 _21688_ (.A1(_08161_),
    .A2(_08662_),
    .A3(_08678_),
    .B1(_02002_),
    .Y(_02003_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_412 ();
 sky130_fd_sc_hd__a21oi_4 _21690_ (.A1(net303),
    .A2(net322),
    .B1(net1053),
    .Y(_02005_));
 sky130_fd_sc_hd__nand2_1 _21691_ (.A(_01998_),
    .B(_02005_),
    .Y(_02006_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_411 ();
 sky130_fd_sc_hd__a21oi_1 _21693_ (.A1(_08760_),
    .A2(_08763_),
    .B1(net321),
    .Y(_02008_));
 sky130_fd_sc_hd__nor4b_4 _21694_ (.A(_08773_),
    .B(_08784_),
    .C(_08793_),
    .D_N(_02008_),
    .Y(_02009_));
 sky130_fd_sc_hd__a21o_4 _21695_ (.A1(net305),
    .A2(net322),
    .B1(net302),
    .X(_02010_));
 sky130_fd_sc_hd__nor2_2 _21696_ (.A(net1224),
    .B(_02010_),
    .Y(_02011_));
 sky130_fd_sc_hd__xnor2_2 _21697_ (.A(_02006_),
    .B(_02011_),
    .Y(_02012_));
 sky130_fd_sc_hd__xor3_4 _21698_ (.A(_01995_),
    .B(_01985_),
    .C(_02012_),
    .X(_02013_));
 sky130_fd_sc_hd__nor2_8 _21699_ (.A(net1214),
    .B(_01976_),
    .Y(_02014_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_410 ();
 sky130_fd_sc_hd__a21oi_4 _21701_ (.A1(_01712_),
    .A2(net660),
    .B1(net1209),
    .Y(_02016_));
 sky130_fd_sc_hd__mux2i_2 _21702_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[49] ),
    .A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[33] ),
    .S(net315),
    .Y(_02017_));
 sky130_fd_sc_hd__a2bb2oi_4 _21703_ (.A1_N(_08280_),
    .A2_N(_02017_),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[49] ),
    .B2(net322),
    .Y(_02018_));
 sky130_fd_sc_hd__xnor3_1 _21704_ (.A(_02014_),
    .B(_02016_),
    .C(_02018_),
    .X(_02019_));
 sky130_fd_sc_hd__and3_2 _21705_ (.A(_01710_),
    .B(_01726_),
    .C(_02019_),
    .X(_02020_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_407 ();
 sky130_fd_sc_hd__a21oi_4 _21709_ (.A1(net305),
    .A2(net322),
    .B1(net302),
    .Y(_02024_));
 sky130_fd_sc_hd__nand2_1 _21710_ (.A(_01998_),
    .B(_02024_),
    .Y(_02025_));
 sky130_fd_sc_hd__nor2_1 _21711_ (.A(_02020_),
    .B(_02025_),
    .Y(_02026_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_406 ();
 sky130_fd_sc_hd__nand2_1 _21713_ (.A(_01998_),
    .B(_02016_),
    .Y(_02028_));
 sky130_fd_sc_hd__nor3_4 _21714_ (.A(_08909_),
    .B(_08915_),
    .C(net321),
    .Y(_02029_));
 sky130_fd_sc_hd__and3_4 _21715_ (.A(_08926_),
    .B(_08940_),
    .C(_08947_),
    .X(_02030_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_405 ();
 sky130_fd_sc_hd__a22oi_4 _21717_ (.A1(_09856_),
    .A2(net321),
    .B1(_02029_),
    .B2(_02030_),
    .Y(_02032_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_404 ();
 sky130_fd_sc_hd__nand2_1 _21719_ (.A(_02032_),
    .B(_02014_),
    .Y(_02034_));
 sky130_fd_sc_hd__o41ai_2 _21720_ (.A1(net945),
    .A2(net1279),
    .A3(net1224),
    .A4(_01982_),
    .B1(_02018_),
    .Y(_02035_));
 sky130_fd_sc_hd__a21boi_4 _21721_ (.A1(_02028_),
    .A2(_02034_),
    .B1_N(_02035_),
    .Y(_02036_));
 sky130_fd_sc_hd__o21a_1 _21722_ (.A1(_08280_),
    .A2(_01963_),
    .B1(_01964_),
    .X(_02037_));
 sky130_fd_sc_hd__xnor3_2 _21723_ (.A(_02037_),
    .B(_01975_),
    .C(_01984_),
    .X(_02038_));
 sky130_fd_sc_hd__or2_1 _21724_ (.A(_02036_),
    .B(_02038_),
    .X(_02039_));
 sky130_fd_sc_hd__nand2_1 _21725_ (.A(_02036_),
    .B(_02038_),
    .Y(_02040_));
 sky130_fd_sc_hd__and2_0 _21726_ (.A(_02039_),
    .B(_02040_),
    .X(_02041_));
 sky130_fd_sc_hd__nand3_1 _21727_ (.A(_02013_),
    .B(_02026_),
    .C(_02041_),
    .Y(_02042_));
 sky130_fd_sc_hd__a21oi_1 _21728_ (.A1(_02039_),
    .A2(_02020_),
    .B1(_02012_),
    .Y(_02043_));
 sky130_fd_sc_hd__a21oi_1 _21729_ (.A1(_02038_),
    .A2(_02020_),
    .B1(_02036_),
    .Y(_02044_));
 sky130_fd_sc_hd__o21ai_0 _21730_ (.A1(_02038_),
    .A2(_02020_),
    .B1(_02012_),
    .Y(_02045_));
 sky130_fd_sc_hd__xnor2_1 _21731_ (.A(_01985_),
    .B(_01995_),
    .Y(_02046_));
 sky130_fd_sc_hd__o21a_1 _21732_ (.A1(_02044_),
    .A2(_02045_),
    .B1(_02046_),
    .X(_02047_));
 sky130_fd_sc_hd__nor2_1 _21733_ (.A(_02046_),
    .B(_02040_),
    .Y(_02048_));
 sky130_fd_sc_hd__nand2_1 _21734_ (.A(_02024_),
    .B(_02020_),
    .Y(_02049_));
 sky130_fd_sc_hd__mux2_4 _21735_ (.A0(_02040_),
    .A1(_02039_),
    .S(_02013_),
    .X(_02050_));
 sky130_fd_sc_hd__o32a_1 _21736_ (.A1(_02043_),
    .A2(_02047_),
    .A3(_02048_),
    .B1(_02049_),
    .B2(_02050_),
    .X(_02051_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_403 ();
 sky130_fd_sc_hd__o21ai_0 _21738_ (.A1(net946),
    .A2(net781),
    .B1(_02037_),
    .Y(_02053_));
 sky130_fd_sc_hd__o221ai_2 _21739_ (.A1(_02053_),
    .A2(_01984_),
    .B1(_01985_),
    .B2(_02036_),
    .C1(_01995_),
    .Y(_02054_));
 sky130_fd_sc_hd__nand4_1 _21740_ (.A(_01965_),
    .B(_01975_),
    .C(_01984_),
    .D(_02036_),
    .Y(_02055_));
 sky130_fd_sc_hd__nand2_1 _21741_ (.A(_02054_),
    .B(_02055_),
    .Y(_02056_));
 sky130_fd_sc_hd__a221oi_4 _21742_ (.A1(net306),
    .A2(net321),
    .B1(net1200),
    .B2(net741),
    .C1(net302),
    .Y(_02057_));
 sky130_fd_sc_hd__a2111oi_4 _21743_ (.A1(net304),
    .A2(net321),
    .B1(_01976_),
    .C1(net1052),
    .D1(net1214),
    .Y(_02058_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_401 ();
 sky130_fd_sc_hd__and4_4 _21746_ (.A(_10024_),
    .B(_10031_),
    .C(_10039_),
    .D(net321),
    .X(_02061_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_399 ();
 sky130_fd_sc_hd__a221oi_4 _21749_ (.A1(net308),
    .A2(net320),
    .B1(_01996_),
    .B2(_01997_),
    .C1(_02061_),
    .Y(_02064_));
 sky130_fd_sc_hd__xnor2_2 _21750_ (.A(_02058_),
    .B(_02064_),
    .Y(_02065_));
 sky130_fd_sc_hd__xor2_4 _21751_ (.A(net958),
    .B(_02065_),
    .X(_02066_));
 sky130_fd_sc_hd__o21ai_1 _21752_ (.A1(_08280_),
    .A2(_01986_),
    .B1(_01987_),
    .Y(_02067_));
 sky130_fd_sc_hd__maj3_1 _21753_ (.A(_02067_),
    .B(_01989_),
    .C(_01994_),
    .X(_02068_));
 sky130_fd_sc_hd__mux2i_1 _21754_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[52] ),
    .A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[36] ),
    .S(net315),
    .Y(_02069_));
 sky130_fd_sc_hd__nand2_1 _21755_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[52] ),
    .B(net322),
    .Y(_02070_));
 sky130_fd_sc_hd__o21ai_1 _21756_ (.A1(_08280_),
    .A2(_02069_),
    .B1(_02070_),
    .Y(_02071_));
 sky130_fd_sc_hd__nor2_4 _21757_ (.A(_08512_),
    .B(_01968_),
    .Y(_02072_));
 sky130_fd_sc_hd__nand3_1 _21758_ (.A(_10048_),
    .B(_10051_),
    .C(_02072_),
    .Y(_02073_));
 sky130_fd_sc_hd__nor2_4 _21759_ (.A(_08512_),
    .B(_01720_),
    .Y(_02074_));
 sky130_fd_sc_hd__nand3_1 _21760_ (.A(_08558_),
    .B(_08563_),
    .C(_02074_),
    .Y(_02075_));
 sky130_fd_sc_hd__nor2_8 _21761_ (.A(net386),
    .B(_01968_),
    .Y(_02076_));
 sky130_fd_sc_hd__o311ai_4 _21762_ (.A1(net392),
    .A2(_10054_),
    .A3(_10056_),
    .B1(_02076_),
    .C1(_10059_),
    .Y(_02077_));
 sky130_fd_sc_hd__nor2_4 _21763_ (.A(net386),
    .B(_01720_),
    .Y(_02078_));
 sky130_fd_sc_hd__o311ai_4 _21764_ (.A1(net977),
    .A2(_08567_),
    .A3(_08570_),
    .B1(_02078_),
    .C1(_08573_),
    .Y(_02079_));
 sky130_fd_sc_hd__nand4_4 _21765_ (.A(_02073_),
    .B(_02075_),
    .C(_02077_),
    .D(_02079_),
    .Y(_02080_));
 sky130_fd_sc_hd__a221oi_2 _21766_ (.A1(_09856_),
    .A2(net321),
    .B1(_02029_),
    .B2(_02030_),
    .C1(_02080_),
    .Y(_02081_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_398 ();
 sky130_fd_sc_hd__or3_4 _21768_ (.A(_08617_),
    .B(_08629_),
    .C(_01720_),
    .X(_02083_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_397 ();
 sky130_fd_sc_hd__nand4_4 _21770_ (.A(_09951_),
    .B(_09955_),
    .C(_09968_),
    .D(_01720_),
    .Y(_02085_));
 sky130_fd_sc_hd__a221oi_2 _21771_ (.A1(_08995_),
    .A2(net320),
    .B1(_02083_),
    .B2(_02085_),
    .C1(_01980_),
    .Y(_02086_));
 sky130_fd_sc_hd__xor3_2 _21772_ (.A(_02071_),
    .B(_02081_),
    .C(_02086_),
    .X(_02087_));
 sky130_fd_sc_hd__a21o_4 _21773_ (.A1(net303),
    .A2(net322),
    .B1(net1053),
    .X(_02088_));
 sky130_fd_sc_hd__a32oi_4 _21774_ (.A1(_01719_),
    .A2(_09751_),
    .A3(_01720_),
    .B1(_01724_),
    .B2(net562),
    .Y(_02089_));
 sky130_fd_sc_hd__nor3_2 _21775_ (.A(_02010_),
    .B(_02088_),
    .C(_02089_),
    .Y(_02090_));
 sky130_fd_sc_hd__xor2_1 _21776_ (.A(_02087_),
    .B(_02090_),
    .X(_02091_));
 sky130_fd_sc_hd__xnor2_1 _21777_ (.A(_02068_),
    .B(_02091_),
    .Y(_02092_));
 sky130_fd_sc_hd__xor2_1 _21778_ (.A(_02066_),
    .B(_02092_),
    .X(_02093_));
 sky130_fd_sc_hd__xnor2_1 _21779_ (.A(_02056_),
    .B(_02093_),
    .Y(_02094_));
 sky130_fd_sc_hd__a21o_4 _21780_ (.A1(_02051_),
    .A2(_02042_),
    .B1(_02094_),
    .X(_02095_));
 sky130_fd_sc_hd__nand3_1 _21781_ (.A(_02094_),
    .B(_02042_),
    .C(_02051_),
    .Y(_02096_));
 sky130_fd_sc_hd__nand2_2 _21782_ (.A(_02095_),
    .B(_02096_),
    .Y(_02097_));
 sky130_fd_sc_hd__nand2_1 _21783_ (.A(_01700_),
    .B(_02097_),
    .Y(_02098_));
 sky130_fd_sc_hd__o21ai_0 _21784_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[36] ),
    .A2(_01700_),
    .B1(_02098_),
    .Y(_02099_));
 sky130_fd_sc_hd__nand2_2 _21785_ (.A(net312),
    .B(_02099_),
    .Y(_02100_));
 sky130_fd_sc_hd__nand2_2 _21786_ (.A(_01959_),
    .B(_02100_),
    .Y(_02101_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_396 ();
 sky130_fd_sc_hd__nand2_1 _21788_ (.A(\load_store_unit_i.rdata_offset_q[1] ),
    .B(net39),
    .Y(_02103_));
 sky130_fd_sc_hd__nor2_1 _21789_ (.A(\load_store_unit_i.rdata_offset_q[0] ),
    .B(_02103_),
    .Y(_02104_));
 sky130_fd_sc_hd__a21oi_1 _21790_ (.A1(net30),
    .A2(_01672_),
    .B1(_02104_),
    .Y(_02105_));
 sky130_fd_sc_hd__a221oi_1 _21791_ (.A1(\load_store_unit_i.rdata_q[12] ),
    .A2(_01672_),
    .B1(_01683_),
    .B2(\load_store_unit_i.rdata_q[20] ),
    .C1(_01684_),
    .Y(_02106_));
 sky130_fd_sc_hd__a21oi_1 _21792_ (.A1(_01684_),
    .A2(_02105_),
    .B1(_02106_),
    .Y(_02107_));
 sky130_fd_sc_hd__a22oi_1 _21793_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(net47),
    .B1(_01688_),
    .B2(\load_store_unit_i.rdata_q[28] ),
    .Y(_02108_));
 sky130_fd_sc_hd__nand2_1 _21794_ (.A(_01682_),
    .B(net53),
    .Y(_02109_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_395 ();
 sky130_fd_sc_hd__o22ai_1 _21796_ (.A1(_01693_),
    .A2(_02108_),
    .B1(_02109_),
    .B2(\load_store_unit_i.rdata_offset_q[0] ),
    .Y(_02111_));
 sky130_fd_sc_hd__nor3_1 _21797_ (.A(net267),
    .B(_02107_),
    .C(_02111_),
    .Y(_02112_));
 sky130_fd_sc_hd__a31oi_4 _21798_ (.A1(_11885_),
    .A2(net267),
    .A3(_02101_),
    .B1(_02112_),
    .Y(_02113_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_394 ();
 sky130_fd_sc_hd__or2_2 _21800_ (.A(net267),
    .B(_01911_),
    .X(_02115_));
 sky130_fd_sc_hd__nand2_2 _21801_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .B(_02115_),
    .Y(_02116_));
 sky130_fd_sc_hd__or2_4 _21802_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .B(_02116_),
    .X(_02117_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_393 ();
 sky130_fd_sc_hd__nor2_8 _21804_ (.A(_08194_),
    .B(_02117_),
    .Y(_02119_));
 sky130_fd_sc_hd__nand2_1 _21805_ (.A(_02113_),
    .B(_02119_),
    .Y(_02120_));
 sky130_fd_sc_hd__nor3_4 _21806_ (.A(net1020),
    .B(net331),
    .C(net447),
    .Y(_02121_));
 sky130_fd_sc_hd__nor2_8 _21807_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .B(_02116_),
    .Y(_02122_));
 sky130_fd_sc_hd__nand2_8 _21808_ (.A(_02121_),
    .B(_02122_),
    .Y(_02123_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_392 ();
 sky130_fd_sc_hd__nand2_1 _21810_ (.A(\gen_regfile_ff.register_file_i.rf_reg[132] ),
    .B(_02123_),
    .Y(_02125_));
 sky130_fd_sc_hd__nand2_1 _21811_ (.A(_02120_),
    .B(_02125_),
    .Y(_00515_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_390 ();
 sky130_fd_sc_hd__nand2_1 _21814_ (.A(_02066_),
    .B(_02092_),
    .Y(_02128_));
 sky130_fd_sc_hd__o211ai_1 _21815_ (.A1(_02066_),
    .A2(_02092_),
    .B1(_02054_),
    .C1(_02055_),
    .Y(_02129_));
 sky130_fd_sc_hd__nand2_1 _21816_ (.A(_02128_),
    .B(_02129_),
    .Y(_02130_));
 sky130_fd_sc_hd__and4_4 _21817_ (.A(_10089_),
    .B(net902),
    .C(_10109_),
    .D(net321),
    .X(_02131_));
 sky130_fd_sc_hd__a21oi_4 _21818_ (.A1(_10865_),
    .A2(net320),
    .B1(_02131_),
    .Y(_02132_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_389 ();
 sky130_fd_sc_hd__nand2_2 _21820_ (.A(_01998_),
    .B(_02132_),
    .Y(_02134_));
 sky130_fd_sc_hd__a221oi_4 _21821_ (.A1(net305),
    .A2(net321),
    .B1(_02083_),
    .B2(_02085_),
    .C1(net302),
    .Y(_02135_));
 sky130_fd_sc_hd__a221oi_4 _21822_ (.A1(net303),
    .A2(net321),
    .B1(net741),
    .B2(net1200),
    .C1(net1052),
    .Y(_02136_));
 sky130_fd_sc_hd__xor2_2 _21823_ (.A(_02135_),
    .B(_02136_),
    .X(_02137_));
 sky130_fd_sc_hd__a2111oi_4 _21824_ (.A1(net308),
    .A2(net320),
    .B1(_01976_),
    .C1(_02061_),
    .D1(net1214),
    .Y(_02138_));
 sky130_fd_sc_hd__xnor2_2 _21825_ (.A(_02137_),
    .B(net1068),
    .Y(_02139_));
 sky130_fd_sc_hd__xor2_2 _21826_ (.A(_02134_),
    .B(_02139_),
    .X(_02140_));
 sky130_fd_sc_hd__or2_0 _21827_ (.A(_02087_),
    .B(_02090_),
    .X(_02141_));
 sky130_fd_sc_hd__and2_0 _21828_ (.A(_02087_),
    .B(_02090_),
    .X(_02142_));
 sky130_fd_sc_hd__mux2i_1 _21829_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[53] ),
    .A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[37] ),
    .S(net315),
    .Y(_02143_));
 sky130_fd_sc_hd__nand2_1 _21830_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[53] ),
    .B(net322),
    .Y(_02144_));
 sky130_fd_sc_hd__o21ai_1 _21831_ (.A1(_08280_),
    .A2(_02143_),
    .B1(_02144_),
    .Y(_02145_));
 sky130_fd_sc_hd__nand3_1 _21832_ (.A(_10117_),
    .B(_10120_),
    .C(_02072_),
    .Y(_02146_));
 sky130_fd_sc_hd__nand3_2 _21833_ (.A(_09091_),
    .B(_09094_),
    .C(_02074_),
    .Y(_02147_));
 sky130_fd_sc_hd__o311ai_4 _21834_ (.A1(net1075),
    .A2(_10123_),
    .A3(_10125_),
    .B1(_02076_),
    .C1(_10128_),
    .Y(_02148_));
 sky130_fd_sc_hd__o311ai_4 _21835_ (.A1(net976),
    .A2(_09097_),
    .A3(_09099_),
    .B1(_02078_),
    .C1(_09102_),
    .Y(_02149_));
 sky130_fd_sc_hd__nand4_4 _21836_ (.A(_02146_),
    .B(_02147_),
    .C(_02148_),
    .D(_02149_),
    .Y(_02150_));
 sky130_fd_sc_hd__a221oi_2 _21837_ (.A1(_09856_),
    .A2(net321),
    .B1(_02029_),
    .B2(_02030_),
    .C1(_02150_),
    .Y(_02151_));
 sky130_fd_sc_hd__a211oi_1 _21838_ (.A1(_08995_),
    .A2(net320),
    .B1(_01980_),
    .C1(_02080_),
    .Y(_02152_));
 sky130_fd_sc_hd__xor3_1 _21839_ (.A(_02145_),
    .B(_02151_),
    .C(_02152_),
    .X(_02153_));
 sky130_fd_sc_hd__maj3_2 _21840_ (.A(_02058_),
    .B(_02057_),
    .C(_02064_),
    .X(_02154_));
 sky130_fd_sc_hd__maj3_1 _21841_ (.A(_02071_),
    .B(_02081_),
    .C(_02086_),
    .X(_02155_));
 sky130_fd_sc_hd__xor3_1 _21842_ (.A(_02153_),
    .B(_02154_),
    .C(_02155_),
    .X(_02156_));
 sky130_fd_sc_hd__a211oi_2 _21843_ (.A1(_02068_),
    .A2(_02141_),
    .B1(_02142_),
    .C1(_02156_),
    .Y(_02157_));
 sky130_fd_sc_hd__nand2_8 _21844_ (.A(net742),
    .B(net1200),
    .Y(_02158_));
 sky130_fd_sc_hd__nand2_1 _21845_ (.A(_02158_),
    .B(net984),
    .Y(_02159_));
 sky130_fd_sc_hd__nand2_4 _21846_ (.A(_02083_),
    .B(_02085_),
    .Y(_02160_));
 sky130_fd_sc_hd__nand2_1 _21847_ (.A(_02032_),
    .B(_02160_),
    .Y(_02161_));
 sky130_fd_sc_hd__a21oi_1 _21848_ (.A1(_02159_),
    .A2(_02161_),
    .B1(_01988_),
    .Y(_02162_));
 sky130_fd_sc_hd__nor2_1 _21849_ (.A(_02159_),
    .B(_02161_),
    .Y(_02163_));
 sky130_fd_sc_hd__o311a_4 _21850_ (.A1(_02162_),
    .A2(_02163_),
    .A3(_02142_),
    .B1(_02156_),
    .C1(_02141_),
    .X(_02164_));
 sky130_fd_sc_hd__nor2_4 _21851_ (.A(_02157_),
    .B(_02164_),
    .Y(_02165_));
 sky130_fd_sc_hd__xnor2_2 _21852_ (.A(_02140_),
    .B(_02165_),
    .Y(_02166_));
 sky130_fd_sc_hd__xnor2_2 _21853_ (.A(_02130_),
    .B(_02166_),
    .Y(_02167_));
 sky130_fd_sc_hd__xor2_2 _21854_ (.A(_02095_),
    .B(_02167_),
    .X(_02168_));
 sky130_fd_sc_hd__or3_4 _21855_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .C(net316),
    .X(_02169_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_387 ();
 sky130_fd_sc_hd__mux2i_4 _21858_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[37] ),
    .A1(_02168_),
    .S(_02169_),
    .Y(_02172_));
 sky130_fd_sc_hd__nand2_1 _21859_ (.A(net443),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[37] ),
    .Y(_02173_));
 sky130_fd_sc_hd__o21ai_4 _21860_ (.A1(net443),
    .A2(_02172_),
    .B1(_02173_),
    .Y(_02174_));
 sky130_fd_sc_hd__mux2i_4 _21861_ (.A0(_01817_),
    .A1(_01819_),
    .S(net299),
    .Y(_02175_));
 sky130_fd_sc_hd__nor2_1 _21862_ (.A(net299),
    .B(_01821_),
    .Y(_02176_));
 sky130_fd_sc_hd__nor2_1 _21863_ (.A(net1467),
    .B(_01781_),
    .Y(_02177_));
 sky130_fd_sc_hd__nor2_1 _21864_ (.A(_02176_),
    .B(_02177_),
    .Y(_02178_));
 sky130_fd_sc_hd__nand2_1 _21865_ (.A(_01751_),
    .B(_02178_),
    .Y(_02179_));
 sky130_fd_sc_hd__o21ai_2 _21866_ (.A1(_01751_),
    .A2(_02175_),
    .B1(_02179_),
    .Y(_02180_));
 sky130_fd_sc_hd__mux2i_1 _21867_ (.A0(_01784_),
    .A1(_01775_),
    .S(net300),
    .Y(_02181_));
 sky130_fd_sc_hd__nand2_1 _21868_ (.A(_01751_),
    .B(_01935_),
    .Y(_02182_));
 sky130_fd_sc_hd__o21ai_2 _21869_ (.A1(_01751_),
    .A2(_02181_),
    .B1(_02182_),
    .Y(_02183_));
 sky130_fd_sc_hd__mux2i_2 _21870_ (.A0(_02180_),
    .A1(_02183_),
    .S(_01748_),
    .Y(_02184_));
 sky130_fd_sc_hd__nand2_1 _21871_ (.A(_01771_),
    .B(_01936_),
    .Y(_02185_));
 sky130_fd_sc_hd__o21ai_2 _21872_ (.A1(_01771_),
    .A2(_01766_),
    .B1(_02185_),
    .Y(_02186_));
 sky130_fd_sc_hd__a21oi_1 _21873_ (.A1(_01758_),
    .A2(_02186_),
    .B1(_01947_),
    .Y(_02187_));
 sky130_fd_sc_hd__nand2_1 _21874_ (.A(_01826_),
    .B(_02187_),
    .Y(_02188_));
 sky130_fd_sc_hd__o21ai_2 _21875_ (.A1(_01826_),
    .A2(_02184_),
    .B1(_02188_),
    .Y(_02189_));
 sky130_fd_sc_hd__mux2i_4 _21876_ (.A0(_01830_),
    .A1(_01838_),
    .S(net300),
    .Y(_02190_));
 sky130_fd_sc_hd__nand2_1 _21877_ (.A(net1468),
    .B(_01841_),
    .Y(_02191_));
 sky130_fd_sc_hd__o21ai_2 _21878_ (.A1(net1469),
    .A2(_01861_),
    .B1(_02191_),
    .Y(_02192_));
 sky130_fd_sc_hd__mux2i_4 _21879_ (.A0(_02190_),
    .A1(_02192_),
    .S(_01751_),
    .Y(_02193_));
 sky130_fd_sc_hd__nor2_1 _21880_ (.A(_01748_),
    .B(_02193_),
    .Y(_02194_));
 sky130_fd_sc_hd__mux2i_2 _21881_ (.A0(_01862_),
    .A1(_01864_),
    .S(net300),
    .Y(_02195_));
 sky130_fd_sc_hd__mux2i_4 _21882_ (.A0(_01866_),
    .A1(_01869_),
    .S(net299),
    .Y(_02196_));
 sky130_fd_sc_hd__mux2i_2 _21883_ (.A0(_02195_),
    .A1(_02196_),
    .S(_01751_),
    .Y(_02197_));
 sky130_fd_sc_hd__nor2_1 _21884_ (.A(_01758_),
    .B(_02197_),
    .Y(_02198_));
 sky130_fd_sc_hd__xnor2_1 _21885_ (.A(net1466),
    .B(net294),
    .Y(_02199_));
 sky130_fd_sc_hd__mux2i_1 _21886_ (.A0(_09679_),
    .A1(_09825_),
    .S(_02199_),
    .Y(_02200_));
 sky130_fd_sc_hd__nand2_1 _21887_ (.A(net299),
    .B(_01874_),
    .Y(_02201_));
 sky130_fd_sc_hd__o21ai_2 _21888_ (.A1(net299),
    .A2(_01870_),
    .B1(_02201_),
    .Y(_02202_));
 sky130_fd_sc_hd__nand2_1 _21889_ (.A(_01771_),
    .B(_02202_),
    .Y(_02203_));
 sky130_fd_sc_hd__o21ai_1 _21890_ (.A1(_01771_),
    .A2(_02200_),
    .B1(_02203_),
    .Y(_02204_));
 sky130_fd_sc_hd__mux2i_4 _21891_ (.A0(_01811_),
    .A1(_01816_),
    .S(net299),
    .Y(_02205_));
 sky130_fd_sc_hd__nor2_1 _21892_ (.A(net1466),
    .B(_01810_),
    .Y(_02206_));
 sky130_fd_sc_hd__a21oi_1 _21893_ (.A1(net1466),
    .A2(_01807_),
    .B1(_02206_),
    .Y(_02207_));
 sky130_fd_sc_hd__nand2_1 _21894_ (.A(_01771_),
    .B(_02207_),
    .Y(_02208_));
 sky130_fd_sc_hd__o21ai_2 _21895_ (.A1(_01771_),
    .A2(_02205_),
    .B1(_02208_),
    .Y(_02209_));
 sky130_fd_sc_hd__nor2_1 _21896_ (.A(_01758_),
    .B(_02209_),
    .Y(_02210_));
 sky130_fd_sc_hd__a21oi_1 _21897_ (.A1(_01758_),
    .A2(_02204_),
    .B1(_02210_),
    .Y(_02211_));
 sky130_fd_sc_hd__nand2_1 _21898_ (.A(_01826_),
    .B(_02211_),
    .Y(_02212_));
 sky130_fd_sc_hd__o311ai_4 _21899_ (.A1(_01826_),
    .A2(_02194_),
    .A3(_02198_),
    .B1(_02212_),
    .C1(_01743_),
    .Y(_02213_));
 sky130_fd_sc_hd__o21ai_4 _21900_ (.A1(_01743_),
    .A2(_02189_),
    .B1(_02213_),
    .Y(_02214_));
 sky130_fd_sc_hd__nand2_1 _21901_ (.A(_01751_),
    .B(_01794_),
    .Y(_02215_));
 sky130_fd_sc_hd__o21ai_1 _21902_ (.A1(_01751_),
    .A2(_01779_),
    .B1(_02215_),
    .Y(_02216_));
 sky130_fd_sc_hd__nor2_1 _21903_ (.A(_01751_),
    .B(_01798_),
    .Y(_02217_));
 sky130_fd_sc_hd__a21oi_2 _21904_ (.A1(_01756_),
    .A2(_01751_),
    .B1(_02217_),
    .Y(_02218_));
 sky130_fd_sc_hd__nand2_1 _21905_ (.A(_01748_),
    .B(_02218_),
    .Y(_02219_));
 sky130_fd_sc_hd__o21ai_2 _21906_ (.A1(_01748_),
    .A2(_02216_),
    .B1(_02219_),
    .Y(_02220_));
 sky130_fd_sc_hd__nand2_1 _21907_ (.A(_01756_),
    .B(_01746_),
    .Y(_02221_));
 sky130_fd_sc_hd__o21ai_0 _21908_ (.A1(_01746_),
    .A2(_02220_),
    .B1(_02221_),
    .Y(_02222_));
 sky130_fd_sc_hd__nand2_1 _21909_ (.A(net295),
    .B(_02222_),
    .Y(_02223_));
 sky130_fd_sc_hd__o211ai_4 _21910_ (.A1(net295),
    .A2(_02214_),
    .B1(_02223_),
    .C1(_01734_),
    .Y(_02224_));
 sky130_fd_sc_hd__nand2_8 _21911_ (.A(_01890_),
    .B(_01892_),
    .Y(_02225_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_385 ();
 sky130_fd_sc_hd__or2_4 _21914_ (.A(_08429_),
    .B(net647),
    .X(_02228_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_383 ();
 sky130_fd_sc_hd__nand3_1 _21917_ (.A(_09111_),
    .B(_10868_),
    .C(_02228_),
    .Y(_02231_));
 sky130_fd_sc_hd__o21ai_0 _21918_ (.A1(_10868_),
    .A2(_01902_),
    .B1(_02231_),
    .Y(_02232_));
 sky130_fd_sc_hd__nand2_8 _21919_ (.A(_02225_),
    .B(_01896_),
    .Y(_02233_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_381 ();
 sky130_fd_sc_hd__a21oi_1 _21922_ (.A1(_10868_),
    .A2(_02233_),
    .B1(_09111_),
    .Y(_02236_));
 sky130_fd_sc_hd__a21oi_1 _21923_ (.A1(_02225_),
    .A2(_02232_),
    .B1(_02236_),
    .Y(_02237_));
 sky130_fd_sc_hd__a21oi_1 _21924_ (.A1(net176),
    .A2(_01929_),
    .B1(_02237_),
    .Y(_02238_));
 sky130_fd_sc_hd__nand3_1 _21925_ (.A(net739),
    .B(_02224_),
    .C(_02238_),
    .Y(_02239_));
 sky130_fd_sc_hd__o21ai_4 _21926_ (.A1(_08290_),
    .A2(_02174_),
    .B1(_02239_),
    .Y(_02240_));
 sky130_fd_sc_hd__nand2_1 _21927_ (.A(\load_store_unit_i.rdata_offset_q[1] ),
    .B(net40),
    .Y(_02241_));
 sky130_fd_sc_hd__nor2_1 _21928_ (.A(\load_store_unit_i.rdata_offset_q[0] ),
    .B(_02241_),
    .Y(_02242_));
 sky130_fd_sc_hd__a21oi_1 _21929_ (.A1(net31),
    .A2(_01672_),
    .B1(_02242_),
    .Y(_02243_));
 sky130_fd_sc_hd__a221oi_1 _21930_ (.A1(\load_store_unit_i.rdata_q[13] ),
    .A2(_01672_),
    .B1(_01683_),
    .B2(\load_store_unit_i.rdata_q[21] ),
    .C1(_01684_),
    .Y(_02244_));
 sky130_fd_sc_hd__a21oi_1 _21931_ (.A1(_01684_),
    .A2(_02243_),
    .B1(_02244_),
    .Y(_02245_));
 sky130_fd_sc_hd__a22oi_1 _21932_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(net48),
    .B1(_01688_),
    .B2(\load_store_unit_i.rdata_q[29] ),
    .Y(_02246_));
 sky130_fd_sc_hd__nand2_1 _21933_ (.A(_01682_),
    .B(net54),
    .Y(_02247_));
 sky130_fd_sc_hd__o22ai_1 _21934_ (.A1(_01693_),
    .A2(_02246_),
    .B1(_02247_),
    .B2(\load_store_unit_i.rdata_offset_q[0] ),
    .Y(_02248_));
 sky130_fd_sc_hd__nor3_1 _21935_ (.A(net267),
    .B(_02245_),
    .C(_02248_),
    .Y(_02249_));
 sky130_fd_sc_hd__a31oi_4 _21936_ (.A1(_11900_),
    .A2(net267),
    .A3(_02240_),
    .B1(_02249_),
    .Y(_02250_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_380 ();
 sky130_fd_sc_hd__nand2_1 _21938_ (.A(_02119_),
    .B(_02250_),
    .Y(_02252_));
 sky130_fd_sc_hd__nand2_1 _21939_ (.A(\gen_regfile_ff.register_file_i.rf_reg[133] ),
    .B(_02123_),
    .Y(_02253_));
 sky130_fd_sc_hd__nand2_1 _21940_ (.A(_02252_),
    .B(_02253_),
    .Y(_00516_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_379 ();
 sky130_fd_sc_hd__nand2_1 _21942_ (.A(_01751_),
    .B(_01786_),
    .Y(_02255_));
 sky130_fd_sc_hd__o21ai_2 _21943_ (.A1(_01751_),
    .A2(_01822_),
    .B1(_02255_),
    .Y(_02256_));
 sky130_fd_sc_hd__nor2_1 _21944_ (.A(_01748_),
    .B(_02256_),
    .Y(_02257_));
 sky130_fd_sc_hd__nor2_1 _21945_ (.A(_01758_),
    .B(_02216_),
    .Y(_02258_));
 sky130_fd_sc_hd__nor2_1 _21946_ (.A(_02257_),
    .B(_02258_),
    .Y(_02259_));
 sky130_fd_sc_hd__a211oi_1 _21947_ (.A1(_01758_),
    .A2(_02218_),
    .B1(_01947_),
    .C1(_01738_),
    .Y(_02260_));
 sky130_fd_sc_hd__a21o_1 _21948_ (.A1(_01738_),
    .A2(_02259_),
    .B1(_02260_),
    .X(_02261_));
 sky130_fd_sc_hd__mux2i_2 _21949_ (.A0(_01809_),
    .A1(_01876_),
    .S(_01771_),
    .Y(_02262_));
 sky130_fd_sc_hd__mux2i_2 _21950_ (.A0(_01812_),
    .A1(_01818_),
    .S(_01751_),
    .Y(_02263_));
 sky130_fd_sc_hd__mux2i_2 _21951_ (.A0(_02262_),
    .A1(_02263_),
    .S(_01748_),
    .Y(_02264_));
 sky130_fd_sc_hd__mux2i_2 _21952_ (.A0(_01867_),
    .A1(_01871_),
    .S(_01751_),
    .Y(_02265_));
 sky130_fd_sc_hd__nor2_1 _21953_ (.A(_01751_),
    .B(_01843_),
    .Y(_02266_));
 sky130_fd_sc_hd__nor2_1 _21954_ (.A(_01771_),
    .B(_01863_),
    .Y(_02267_));
 sky130_fd_sc_hd__nor2_1 _21955_ (.A(_02266_),
    .B(_02267_),
    .Y(_02268_));
 sky130_fd_sc_hd__nand2_1 _21956_ (.A(_01758_),
    .B(_02268_),
    .Y(_02269_));
 sky130_fd_sc_hd__o211ai_1 _21957_ (.A1(_01758_),
    .A2(_02265_),
    .B1(_02269_),
    .C1(_01738_),
    .Y(_02270_));
 sky130_fd_sc_hd__o211ai_2 _21958_ (.A1(_01738_),
    .A2(_02264_),
    .B1(_02270_),
    .C1(_01743_),
    .Y(_02271_));
 sky130_fd_sc_hd__o21ai_1 _21959_ (.A1(_01743_),
    .A2(_02261_),
    .B1(_02271_),
    .Y(_02272_));
 sky130_fd_sc_hd__nor2_1 _21960_ (.A(_01748_),
    .B(_02183_),
    .Y(_02273_));
 sky130_fd_sc_hd__a21oi_2 _21961_ (.A1(_01748_),
    .A2(_02186_),
    .B1(_02273_),
    .Y(_02274_));
 sky130_fd_sc_hd__a21oi_1 _21962_ (.A1(_01738_),
    .A2(_02274_),
    .B1(_01941_),
    .Y(_02275_));
 sky130_fd_sc_hd__a21oi_1 _21963_ (.A1(_01743_),
    .A2(_02275_),
    .B1(_01943_),
    .Y(_02276_));
 sky130_fd_sc_hd__nor2_1 _21964_ (.A(_01773_),
    .B(_02276_),
    .Y(_02277_));
 sky130_fd_sc_hd__a21oi_2 _21965_ (.A1(_01773_),
    .A2(_02272_),
    .B1(_02277_),
    .Y(_02278_));
 sky130_fd_sc_hd__nor2_1 _21966_ (.A(net928),
    .B(_01898_),
    .Y(_02279_));
 sky130_fd_sc_hd__a22oi_1 _21967_ (.A1(net928),
    .A2(_01896_),
    .B1(_02279_),
    .B2(_08547_),
    .Y(_02280_));
 sky130_fd_sc_hd__nor2_1 _21968_ (.A(net925),
    .B(_01903_),
    .Y(_02281_));
 sky130_fd_sc_hd__o22ai_1 _21969_ (.A1(_01893_),
    .A2(_02280_),
    .B1(_02281_),
    .B2(_08547_),
    .Y(_02282_));
 sky130_fd_sc_hd__o221ai_1 _21970_ (.A1(_09159_),
    .A2(_01889_),
    .B1(_02278_),
    .B2(_01761_),
    .C1(_02282_),
    .Y(_02283_));
 sky130_fd_sc_hd__nand2_1 _21971_ (.A(_10950_),
    .B(_02169_),
    .Y(_02284_));
 sky130_fd_sc_hd__nor2_2 _21972_ (.A(_02095_),
    .B(_02167_),
    .Y(_02285_));
 sky130_fd_sc_hd__a21oi_2 _21973_ (.A1(net309),
    .A2(_01712_),
    .B1(_02061_),
    .Y(_02286_));
 sky130_fd_sc_hd__nand4_4 _21974_ (.A(_09123_),
    .B(_09130_),
    .C(net499),
    .D(net320),
    .Y(_02287_));
 sky130_fd_sc_hd__nand4_4 _21975_ (.A(_10181_),
    .B(_10188_),
    .C(net1217),
    .D(net321),
    .Y(_02288_));
 sky130_fd_sc_hd__nand2_8 _21976_ (.A(_02287_),
    .B(_02288_),
    .Y(_02289_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_378 ();
 sky130_fd_sc_hd__o2111ai_1 _21978_ (.A1(net1224),
    .A2(_02286_),
    .B1(net1006),
    .C1(_02289_),
    .D1(_01998_),
    .Y(_02291_));
 sky130_fd_sc_hd__a21o_4 _21979_ (.A1(net309),
    .A2(_01712_),
    .B1(_02061_),
    .X(_02292_));
 sky130_fd_sc_hd__nand4_1 _21980_ (.A(_02014_),
    .B(_02292_),
    .C(net1006),
    .D(_02289_),
    .Y(_02293_));
 sky130_fd_sc_hd__xnor2_2 _21981_ (.A(_02135_),
    .B(_02136_),
    .Y(_02294_));
 sky130_fd_sc_hd__mux2i_2 _21982_ (.A0(_02291_),
    .A1(_02293_),
    .S(_02294_),
    .Y(_02295_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_377 ();
 sky130_fd_sc_hd__nor2_1 _21984_ (.A(_01725_),
    .B(_02014_),
    .Y(_02297_));
 sky130_fd_sc_hd__nor3_1 _21985_ (.A(net887),
    .B(_02292_),
    .C(_02089_),
    .Y(_02298_));
 sky130_fd_sc_hd__and4_4 _21986_ (.A(_09123_),
    .B(_09130_),
    .C(net499),
    .D(net320),
    .X(_02299_));
 sky130_fd_sc_hd__and4_4 _21987_ (.A(_10181_),
    .B(_10188_),
    .C(net1217),
    .D(net321),
    .X(_02300_));
 sky130_fd_sc_hd__nor2_8 _21988_ (.A(_02299_),
    .B(_02300_),
    .Y(_02301_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_376 ();
 sky130_fd_sc_hd__o211a_1 _21990_ (.A1(_02297_),
    .A2(_02298_),
    .B1(_02294_),
    .C1(net1307),
    .X(_02303_));
 sky130_fd_sc_hd__a32o_2 _21991_ (.A1(_09751_),
    .A2(_01719_),
    .A3(_01720_),
    .B1(_01724_),
    .B2(net563),
    .X(_02304_));
 sky130_fd_sc_hd__nand2_1 _21992_ (.A(_02304_),
    .B(net1307),
    .Y(_02305_));
 sky130_fd_sc_hd__nor3_1 _21993_ (.A(_02294_),
    .B(net1067),
    .C(_02305_),
    .Y(_02306_));
 sky130_fd_sc_hd__nand4_4 _21994_ (.A(_10089_),
    .B(net1174),
    .C(_10109_),
    .D(net321),
    .Y(_02307_));
 sky130_fd_sc_hd__o21ai_4 _21995_ (.A1(net913),
    .A2(net321),
    .B1(_02307_),
    .Y(_02308_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_375 ();
 sky130_fd_sc_hd__nor3_2 _21997_ (.A(_01998_),
    .B(net887),
    .C(net908),
    .Y(_02310_));
 sky130_fd_sc_hd__nor3_1 _21998_ (.A(_01725_),
    .B(net1006),
    .C(_02289_),
    .Y(_02311_));
 sky130_fd_sc_hd__or2_0 _21999_ (.A(_02310_),
    .B(_02311_),
    .X(_02312_));
 sky130_fd_sc_hd__a211oi_2 _22000_ (.A1(net305),
    .A2(net322),
    .B1(net302),
    .C1(_02080_),
    .Y(_02313_));
 sky130_fd_sc_hd__a221oi_4 _22001_ (.A1(net303),
    .A2(net322),
    .B1(_02083_),
    .B2(_02085_),
    .C1(net1053),
    .Y(_02314_));
 sky130_fd_sc_hd__a221oi_4 _22002_ (.A1(net308),
    .A2(net320),
    .B1(net1200),
    .B2(net741),
    .C1(_02061_),
    .Y(_02315_));
 sky130_fd_sc_hd__xnor2_1 _22003_ (.A(_02314_),
    .B(_02315_),
    .Y(_02316_));
 sky130_fd_sc_hd__xnor2_1 _22004_ (.A(_02313_),
    .B(_02316_),
    .Y(_02317_));
 sky130_fd_sc_hd__o41ai_2 _22005_ (.A1(_02312_),
    .A2(_02303_),
    .A3(_02306_),
    .A4(_02295_),
    .B1(_02317_),
    .Y(_02318_));
 sky130_fd_sc_hd__nor3_1 _22006_ (.A(_02089_),
    .B(net1067),
    .C(_02289_),
    .Y(_02319_));
 sky130_fd_sc_hd__a211oi_1 _22007_ (.A1(_02137_),
    .A2(_02319_),
    .B1(_02310_),
    .C1(_02311_),
    .Y(_02320_));
 sky130_fd_sc_hd__or4b_4 _22008_ (.A(_02317_),
    .B(_02295_),
    .C(_02303_),
    .D_N(_02320_),
    .X(_02321_));
 sky130_fd_sc_hd__nand2_2 _22009_ (.A(_02318_),
    .B(_02321_),
    .Y(_02322_));
 sky130_fd_sc_hd__maj3_2 _22010_ (.A(_02135_),
    .B(_02136_),
    .C(_02138_),
    .X(_02323_));
 sky130_fd_sc_hd__mux2i_1 _22011_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[54] ),
    .A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[38] ),
    .S(net315),
    .Y(_02324_));
 sky130_fd_sc_hd__nand2_1 _22012_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[54] ),
    .B(net322),
    .Y(_02325_));
 sky130_fd_sc_hd__o21ai_1 _22013_ (.A1(_08280_),
    .A2(_02324_),
    .B1(_02325_),
    .Y(_02326_));
 sky130_fd_sc_hd__nand3_1 _22014_ (.A(_10155_),
    .B(_10158_),
    .C(_02072_),
    .Y(_02327_));
 sky130_fd_sc_hd__nand3_1 _22015_ (.A(net1073),
    .B(_08525_),
    .C(_02074_),
    .Y(_02328_));
 sky130_fd_sc_hd__o311ai_4 _22016_ (.A1(net976),
    .A2(_10161_),
    .A3(_10163_),
    .B1(_02076_),
    .C1(_10166_),
    .Y(_02329_));
 sky130_fd_sc_hd__o311ai_2 _22017_ (.A1(net975),
    .A2(_08532_),
    .A3(_08536_),
    .B1(_02078_),
    .C1(_08542_),
    .Y(_02330_));
 sky130_fd_sc_hd__nand4_4 _22018_ (.A(_02328_),
    .B(_02327_),
    .C(_02329_),
    .D(_02330_),
    .Y(_02331_));
 sky130_fd_sc_hd__a221oi_2 _22019_ (.A1(_09856_),
    .A2(net321),
    .B1(_02029_),
    .B2(_02030_),
    .C1(_02331_),
    .Y(_02332_));
 sky130_fd_sc_hd__a211oi_1 _22020_ (.A1(_08995_),
    .A2(net320),
    .B1(_01980_),
    .C1(_02150_),
    .Y(_02333_));
 sky130_fd_sc_hd__xor3_1 _22021_ (.A(_02326_),
    .B(_02332_),
    .C(_02333_),
    .X(_02334_));
 sky130_fd_sc_hd__maj3_1 _22022_ (.A(_02145_),
    .B(_02151_),
    .C(_02152_),
    .X(_02335_));
 sky130_fd_sc_hd__xnor3_2 _22023_ (.A(_02335_),
    .B(_02334_),
    .C(_02323_),
    .X(_02336_));
 sky130_fd_sc_hd__maj3_1 _22024_ (.A(_02153_),
    .B(_02154_),
    .C(_02155_),
    .X(_02337_));
 sky130_fd_sc_hd__xnor2_2 _22025_ (.A(_02336_),
    .B(_02337_),
    .Y(_02338_));
 sky130_fd_sc_hd__xnor2_2 _22026_ (.A(_02164_),
    .B(_02338_),
    .Y(_02339_));
 sky130_fd_sc_hd__xnor2_2 _22027_ (.A(_02322_),
    .B(_02339_),
    .Y(_02340_));
 sky130_fd_sc_hd__nor2_1 _22028_ (.A(_02140_),
    .B(_02165_),
    .Y(_02341_));
 sky130_fd_sc_hd__a22oi_2 _22029_ (.A1(_02128_),
    .A2(_02129_),
    .B1(_02140_),
    .B2(_02165_),
    .Y(_02342_));
 sky130_fd_sc_hd__nor2_1 _22030_ (.A(_02341_),
    .B(_02342_),
    .Y(_02343_));
 sky130_fd_sc_hd__xnor2_2 _22031_ (.A(_02340_),
    .B(_02343_),
    .Y(_02344_));
 sky130_fd_sc_hd__xor2_4 _22032_ (.A(_02285_),
    .B(_02344_),
    .X(_02345_));
 sky130_fd_sc_hd__nor2_1 _22033_ (.A(_02284_),
    .B(_02345_),
    .Y(_02346_));
 sky130_fd_sc_hd__nor2_1 _22034_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[38] ),
    .B(_01700_),
    .Y(_02347_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_374 ();
 sky130_fd_sc_hd__o21ai_4 _22036_ (.A1(_02346_),
    .A2(_02347_),
    .B1(net312),
    .Y(_02349_));
 sky130_fd_sc_hd__o21ai_2 _22037_ (.A1(_08272_),
    .A2(_02283_),
    .B1(_02349_),
    .Y(_02350_));
 sky130_fd_sc_hd__nand2_1 _22038_ (.A(\load_store_unit_i.rdata_offset_q[1] ),
    .B(net41),
    .Y(_02351_));
 sky130_fd_sc_hd__nor2_1 _22039_ (.A(\load_store_unit_i.rdata_offset_q[0] ),
    .B(_02351_),
    .Y(_02352_));
 sky130_fd_sc_hd__a21oi_1 _22040_ (.A1(net32),
    .A2(_01672_),
    .B1(_02352_),
    .Y(_02353_));
 sky130_fd_sc_hd__a221oi_1 _22041_ (.A1(\load_store_unit_i.rdata_q[14] ),
    .A2(_01672_),
    .B1(_01683_),
    .B2(\load_store_unit_i.rdata_q[22] ),
    .C1(_01684_),
    .Y(_02354_));
 sky130_fd_sc_hd__a21oi_1 _22042_ (.A1(_01684_),
    .A2(_02353_),
    .B1(_02354_),
    .Y(_02355_));
 sky130_fd_sc_hd__a22oi_1 _22043_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(net50),
    .B1(_01688_),
    .B2(\load_store_unit_i.rdata_q[30] ),
    .Y(_02356_));
 sky130_fd_sc_hd__nand2_1 _22044_ (.A(_01682_),
    .B(net55),
    .Y(_02357_));
 sky130_fd_sc_hd__o22ai_1 _22045_ (.A1(_01693_),
    .A2(_02356_),
    .B1(_02357_),
    .B2(\load_store_unit_i.rdata_offset_q[0] ),
    .Y(_02358_));
 sky130_fd_sc_hd__nor3_1 _22046_ (.A(net267),
    .B(_02355_),
    .C(_02358_),
    .Y(_02359_));
 sky130_fd_sc_hd__a31oi_4 _22047_ (.A1(_11915_),
    .A2(net267),
    .A3(_02350_),
    .B1(_02359_),
    .Y(_02360_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_373 ();
 sky130_fd_sc_hd__nand2_1 _22049_ (.A(_02119_),
    .B(_02360_),
    .Y(_02362_));
 sky130_fd_sc_hd__nand2_1 _22050_ (.A(\gen_regfile_ff.register_file_i.rf_reg[134] ),
    .B(_02123_),
    .Y(_02363_));
 sky130_fd_sc_hd__nand2_1 _22051_ (.A(_02362_),
    .B(_02363_),
    .Y(_00517_));
 sky130_fd_sc_hd__inv_1 _22052_ (.A(_01768_),
    .Y(_02364_));
 sky130_fd_sc_hd__nand2_1 _22053_ (.A(_01771_),
    .B(_02178_),
    .Y(_02365_));
 sky130_fd_sc_hd__o21ai_1 _22054_ (.A1(_01771_),
    .A2(_02181_),
    .B1(_02365_),
    .Y(_02366_));
 sky130_fd_sc_hd__nand2_1 _22055_ (.A(_01748_),
    .B(_01938_),
    .Y(_02367_));
 sky130_fd_sc_hd__o21ai_1 _22056_ (.A1(_01748_),
    .A2(_02366_),
    .B1(_02367_),
    .Y(_02368_));
 sky130_fd_sc_hd__nand2_1 _22057_ (.A(_01771_),
    .B(_02200_),
    .Y(_02369_));
 sky130_fd_sc_hd__nand2_1 _22058_ (.A(_01751_),
    .B(_02207_),
    .Y(_02370_));
 sky130_fd_sc_hd__nand2_2 _22059_ (.A(_02369_),
    .B(_02370_),
    .Y(_02371_));
 sky130_fd_sc_hd__mux2i_4 _22060_ (.A0(_02175_),
    .A1(_02205_),
    .S(_01771_),
    .Y(_02372_));
 sky130_fd_sc_hd__mux2i_1 _22061_ (.A0(_02371_),
    .A1(_02372_),
    .S(_01748_),
    .Y(_02373_));
 sky130_fd_sc_hd__mux2i_2 _22062_ (.A0(_02192_),
    .A1(_02195_),
    .S(_01751_),
    .Y(_02374_));
 sky130_fd_sc_hd__mux2i_4 _22063_ (.A0(_02202_),
    .A1(_02196_),
    .S(_01771_),
    .Y(_02375_));
 sky130_fd_sc_hd__mux2i_1 _22064_ (.A0(_02374_),
    .A1(_02375_),
    .S(_01748_),
    .Y(_02376_));
 sky130_fd_sc_hd__mux4_1 _22065_ (.A0(_02364_),
    .A1(_02368_),
    .A2(_02373_),
    .A3(_02376_),
    .S0(_01738_),
    .S1(_01743_),
    .X(_02377_));
 sky130_fd_sc_hd__o21ai_1 _22066_ (.A1(_01746_),
    .A2(_01802_),
    .B1(_02221_),
    .Y(_02378_));
 sky130_fd_sc_hd__nor2_1 _22067_ (.A(_01773_),
    .B(_02378_),
    .Y(_02379_));
 sky130_fd_sc_hd__a21oi_2 _22068_ (.A1(_01773_),
    .A2(_02377_),
    .B1(_02379_),
    .Y(_02380_));
 sky130_fd_sc_hd__nor2_1 _22069_ (.A(_08497_),
    .B(_01898_),
    .Y(_02381_));
 sky130_fd_sc_hd__a22oi_1 _22070_ (.A1(_08497_),
    .A2(_01896_),
    .B1(_02381_),
    .B2(_08375_),
    .Y(_02382_));
 sky130_fd_sc_hd__nor2_1 _22071_ (.A(_08497_),
    .B(_01903_),
    .Y(_02383_));
 sky130_fd_sc_hd__o22ai_1 _22072_ (.A1(_01893_),
    .A2(_02382_),
    .B1(_02383_),
    .B2(_08375_),
    .Y(_02384_));
 sky130_fd_sc_hd__o221ai_2 _22073_ (.A1(_09157_),
    .A2(_01889_),
    .B1(_02380_),
    .B2(_01761_),
    .C1(_02384_),
    .Y(_02385_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_371 ();
 sky130_fd_sc_hd__o21a_1 _22076_ (.A1(_02341_),
    .A2(_02342_),
    .B1(_02340_),
    .X(_02388_));
 sky130_fd_sc_hd__or3_1 _22077_ (.A(_02341_),
    .B(_02340_),
    .C(_02342_),
    .X(_02389_));
 sky130_fd_sc_hd__o31a_4 _22078_ (.A1(_02388_),
    .A2(_02167_),
    .A3(_02095_),
    .B1(_02389_),
    .X(_02390_));
 sky130_fd_sc_hd__nand3_4 _22079_ (.A(_10219_),
    .B(net1313),
    .C(_02072_),
    .Y(_02391_));
 sky130_fd_sc_hd__nand3_4 _22080_ (.A(_08350_),
    .B(_08357_),
    .C(_02074_),
    .Y(_02392_));
 sky130_fd_sc_hd__o311ai_4 _22081_ (.A1(_10225_),
    .A2(net390),
    .A3(_10227_),
    .B1(_10230_),
    .C1(_02076_),
    .Y(_02393_));
 sky130_fd_sc_hd__nand2_1 _22082_ (.A(_08512_),
    .B(_01968_),
    .Y(_02394_));
 sky130_fd_sc_hd__a311o_4 _22083_ (.A1(_08309_),
    .A2(_08317_),
    .A3(_08323_),
    .B1(_08333_),
    .C1(_02394_),
    .X(_02395_));
 sky130_fd_sc_hd__nand4_4 _22084_ (.A(_02391_),
    .B(_02392_),
    .C(_02395_),
    .D(_02393_),
    .Y(_02396_));
 sky130_fd_sc_hd__a221oi_2 _22085_ (.A1(_09856_),
    .A2(net321),
    .B1(_02029_),
    .B2(_02030_),
    .C1(_02396_),
    .Y(_02397_));
 sky130_fd_sc_hd__mux2i_1 _22086_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[55] ),
    .A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[39] ),
    .S(net315),
    .Y(_02398_));
 sky130_fd_sc_hd__nand2_1 _22087_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[55] ),
    .B(net322),
    .Y(_02399_));
 sky130_fd_sc_hd__o21ai_2 _22088_ (.A1(_08280_),
    .A2(_02398_),
    .B1(_02399_),
    .Y(_02400_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_370 ();
 sky130_fd_sc_hd__a211oi_2 _22090_ (.A1(net699),
    .A2(net320),
    .B1(_01980_),
    .C1(_02331_),
    .Y(_02402_));
 sky130_fd_sc_hd__xor3_1 _22091_ (.A(_02397_),
    .B(_02400_),
    .C(_02402_),
    .X(_02403_));
 sky130_fd_sc_hd__maj3_1 _22092_ (.A(_02326_),
    .B(_02332_),
    .C(_02333_),
    .X(_02404_));
 sky130_fd_sc_hd__maj3_1 _22093_ (.A(_02313_),
    .B(_02314_),
    .C(_02315_),
    .X(_02405_));
 sky130_fd_sc_hd__xnor3_2 _22094_ (.A(_02403_),
    .B(_02404_),
    .C(_02405_),
    .X(_02406_));
 sky130_fd_sc_hd__maj3_2 _22095_ (.A(_02323_),
    .B(_02334_),
    .C(_02335_),
    .X(_02407_));
 sky130_fd_sc_hd__xnor2_2 _22096_ (.A(_02407_),
    .B(_02406_),
    .Y(_02408_));
 sky130_fd_sc_hd__xnor3_2 _22097_ (.A(_02313_),
    .B(_02315_),
    .C(_02314_),
    .X(_02409_));
 sky130_fd_sc_hd__xnor2_1 _22098_ (.A(net1287),
    .B(net1308),
    .Y(_02410_));
 sky130_fd_sc_hd__xnor2_1 _22099_ (.A(_02409_),
    .B(_02410_),
    .Y(_02411_));
 sky130_fd_sc_hd__nor3_2 _22100_ (.A(_02134_),
    .B(_02139_),
    .C(_02411_),
    .Y(_02412_));
 sky130_fd_sc_hd__nor2_1 _22101_ (.A(_02408_),
    .B(_02412_),
    .Y(_02413_));
 sky130_fd_sc_hd__nand2_1 _22102_ (.A(_02408_),
    .B(_02412_),
    .Y(_02414_));
 sky130_fd_sc_hd__nand2b_1 _22103_ (.A_N(_02413_),
    .B(_02414_),
    .Y(_02415_));
 sky130_fd_sc_hd__nand2b_2 _22104_ (.A_N(_02336_),
    .B(_02337_),
    .Y(_02416_));
 sky130_fd_sc_hd__and4_4 _22105_ (.A(_08468_),
    .B(_08480_),
    .C(_08493_),
    .D(net320),
    .X(_02417_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_369 ();
 sky130_fd_sc_hd__and4_4 _22107_ (.A(_10241_),
    .B(net744),
    .C(_10258_),
    .D(net321),
    .X(_02419_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_368 ();
 sky130_fd_sc_hd__nor2_8 _22109_ (.A(_02417_),
    .B(_02419_),
    .Y(_02421_));
 sky130_fd_sc_hd__xnor2_2 _22110_ (.A(_01972_),
    .B(_02421_),
    .Y(_02422_));
 sky130_fd_sc_hd__nor2_4 _22111_ (.A(net788),
    .B(_02289_),
    .Y(_02423_));
 sky130_fd_sc_hd__nand4_4 _22112_ (.A(_08468_),
    .B(_08480_),
    .C(_08493_),
    .D(net320),
    .Y(_02424_));
 sky130_fd_sc_hd__nand4_4 _22113_ (.A(net745),
    .B(_10241_),
    .C(_10258_),
    .D(net321),
    .Y(_02425_));
 sky130_fd_sc_hd__nand2_8 _22114_ (.A(_02424_),
    .B(_02425_),
    .Y(_02426_));
 sky130_fd_sc_hd__a21oi_1 _22115_ (.A1(_02158_),
    .A2(_02132_),
    .B1(_01998_),
    .Y(_02427_));
 sky130_fd_sc_hd__a21oi_1 _22116_ (.A1(net906),
    .A2(_02426_),
    .B1(_02427_),
    .Y(_02428_));
 sky130_fd_sc_hd__nor3_1 _22117_ (.A(net1279),
    .B(net1170),
    .C(net1216),
    .Y(_02429_));
 sky130_fd_sc_hd__nor3_1 _22118_ (.A(_01998_),
    .B(net1172),
    .C(net906),
    .Y(_02430_));
 sky130_fd_sc_hd__o21ai_2 _22119_ (.A1(_02430_),
    .A2(_02429_),
    .B1(_02423_),
    .Y(_02431_));
 sky130_fd_sc_hd__o221ai_4 _22120_ (.A1(_02134_),
    .A2(_02422_),
    .B1(_02423_),
    .B2(_02428_),
    .C1(_02431_),
    .Y(_02432_));
 sky130_fd_sc_hd__o211ai_2 _22121_ (.A1(net887),
    .A2(net907),
    .B1(net1307),
    .C1(_01998_),
    .Y(_02433_));
 sky130_fd_sc_hd__o211ai_2 _22122_ (.A1(net1279),
    .A2(_02289_),
    .B1(net1171),
    .C1(_02014_),
    .Y(_02434_));
 sky130_fd_sc_hd__a21oi_4 _22123_ (.A1(_02433_),
    .A2(_02434_),
    .B1(_02409_),
    .Y(_02435_));
 sky130_fd_sc_hd__and4_4 _22124_ (.A(_02146_),
    .B(_02147_),
    .C(_02148_),
    .D(_02149_),
    .X(_02436_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_367 ();
 sky130_fd_sc_hd__nand2_1 _22126_ (.A(_02024_),
    .B(_02436_),
    .Y(_02438_));
 sky130_fd_sc_hd__nand2_1 _22127_ (.A(_02160_),
    .B(_02286_),
    .Y(_02439_));
 sky130_fd_sc_hd__and4_4 _22128_ (.A(_02073_),
    .B(_02075_),
    .C(_02077_),
    .D(_02079_),
    .X(_02440_));
 sky130_fd_sc_hd__nand2_1 _22129_ (.A(_02005_),
    .B(_02440_),
    .Y(_02441_));
 sky130_fd_sc_hd__xor3_4 _22130_ (.A(_02438_),
    .B(_02439_),
    .C(_02441_),
    .X(_02442_));
 sky130_fd_sc_hd__xnor2_4 _22131_ (.A(_02442_),
    .B(_02435_),
    .Y(_02443_));
 sky130_fd_sc_hd__xor2_4 _22132_ (.A(_02432_),
    .B(_02443_),
    .X(_02444_));
 sky130_fd_sc_hd__xnor2_2 _22133_ (.A(_02416_),
    .B(_02444_),
    .Y(_02445_));
 sky130_fd_sc_hd__xnor2_2 _22134_ (.A(_02445_),
    .B(_02415_),
    .Y(_02446_));
 sky130_fd_sc_hd__inv_1 _22135_ (.A(_02164_),
    .Y(_02447_));
 sky130_fd_sc_hd__inv_1 _22136_ (.A(_02338_),
    .Y(_02448_));
 sky130_fd_sc_hd__maj3_2 _22137_ (.A(_02447_),
    .B(_02322_),
    .C(_02448_),
    .X(_02449_));
 sky130_fd_sc_hd__xnor2_2 _22138_ (.A(_02449_),
    .B(_02446_),
    .Y(_02450_));
 sky130_fd_sc_hd__xnor2_2 _22139_ (.A(_02390_),
    .B(_02450_),
    .Y(_02451_));
 sky130_fd_sc_hd__nand2_1 _22140_ (.A(_02169_),
    .B(_02451_),
    .Y(_02452_));
 sky130_fd_sc_hd__o21ai_4 _22141_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[39] ),
    .A2(_02169_),
    .B1(_02452_),
    .Y(_02453_));
 sky130_fd_sc_hd__nand2_1 _22142_ (.A(net442),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[39] ),
    .Y(_02454_));
 sky130_fd_sc_hd__o211ai_4 _22143_ (.A1(net442),
    .A2(_02453_),
    .B1(_02454_),
    .C1(net312),
    .Y(_02455_));
 sky130_fd_sc_hd__o21ai_2 _22144_ (.A1(_08272_),
    .A2(_02385_),
    .B1(_02455_),
    .Y(_02456_));
 sky130_fd_sc_hd__nand2_1 _22145_ (.A(\load_store_unit_i.rdata_q[15] ),
    .B(_01674_),
    .Y(_02457_));
 sky130_fd_sc_hd__nand2_1 _22146_ (.A(net33),
    .B(_01684_),
    .Y(_02458_));
 sky130_fd_sc_hd__a221oi_1 _22147_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(net51),
    .B1(_01688_),
    .B2(\load_store_unit_i.rdata_q[31] ),
    .C1(_01682_),
    .Y(_02459_));
 sky130_fd_sc_hd__a31oi_1 _22148_ (.A1(_01682_),
    .A2(_02457_),
    .A3(_02458_),
    .B1(_02459_),
    .Y(_02460_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_366 ();
 sky130_fd_sc_hd__nand2_1 _22150_ (.A(\load_store_unit_i.rdata_q[23] ),
    .B(_01674_),
    .Y(_02462_));
 sky130_fd_sc_hd__nand2_1 _22151_ (.A(net42),
    .B(_01684_),
    .Y(_02463_));
 sky130_fd_sc_hd__nor2_1 _22152_ (.A(\load_store_unit_i.rdata_offset_q[1] ),
    .B(net56),
    .Y(_02464_));
 sky130_fd_sc_hd__a311oi_1 _22153_ (.A1(\load_store_unit_i.rdata_offset_q[1] ),
    .A2(_02462_),
    .A3(_02463_),
    .B1(_02464_),
    .C1(\load_store_unit_i.rdata_offset_q[0] ),
    .Y(_02465_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_365 ();
 sky130_fd_sc_hd__a211oi_2 _22155_ (.A1(\load_store_unit_i.rdata_offset_q[0] ),
    .A2(_02460_),
    .B1(_02465_),
    .C1(net267),
    .Y(_02467_));
 sky130_fd_sc_hd__a31oi_4 _22156_ (.A1(_11933_),
    .A2(net267),
    .A3(_02456_),
    .B1(_02467_),
    .Y(_02468_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_364 ();
 sky130_fd_sc_hd__nand2_1 _22158_ (.A(_02119_),
    .B(_02468_),
    .Y(_02470_));
 sky130_fd_sc_hd__nand2_1 _22159_ (.A(\gen_regfile_ff.register_file_i.rf_reg[135] ),
    .B(_02123_),
    .Y(_02471_));
 sky130_fd_sc_hd__nand2_1 _22160_ (.A(_02470_),
    .B(_02471_),
    .Y(_00518_));
 sky130_fd_sc_hd__mux4_2 _22161_ (.A0(_01735_),
    .A1(_01802_),
    .A2(_01824_),
    .A3(_01878_),
    .S0(_01738_),
    .S1(_01743_),
    .X(_02472_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_363 ();
 sky130_fd_sc_hd__nor2_1 _22163_ (.A(_01826_),
    .B(_02368_),
    .Y(_02474_));
 sky130_fd_sc_hd__a21oi_1 _22164_ (.A1(_01768_),
    .A2(_01826_),
    .B1(_02474_),
    .Y(_02475_));
 sky130_fd_sc_hd__a21oi_1 _22165_ (.A1(_01743_),
    .A2(_02475_),
    .B1(_01943_),
    .Y(_02476_));
 sky130_fd_sc_hd__nor2_1 _22166_ (.A(_01773_),
    .B(_02476_),
    .Y(_02477_));
 sky130_fd_sc_hd__a21oi_2 _22167_ (.A1(_01773_),
    .A2(_02472_),
    .B1(_02477_),
    .Y(_02478_));
 sky130_fd_sc_hd__nor2_1 _22168_ (.A(_09222_),
    .B(_01898_),
    .Y(_02479_));
 sky130_fd_sc_hd__a22oi_1 _22169_ (.A1(_09222_),
    .A2(_01896_),
    .B1(_02479_),
    .B2(_09187_),
    .Y(_02480_));
 sky130_fd_sc_hd__nor2_1 _22170_ (.A(_09222_),
    .B(_01903_),
    .Y(_02481_));
 sky130_fd_sc_hd__o22ai_2 _22171_ (.A1(_01893_),
    .A2(_02480_),
    .B1(_02481_),
    .B2(_09187_),
    .Y(_02482_));
 sky130_fd_sc_hd__o221ai_4 _22172_ (.A1(_09303_),
    .A2(_01889_),
    .B1(_02478_),
    .B2(_01761_),
    .C1(_02482_),
    .Y(_02483_));
 sky130_fd_sc_hd__and2_4 _22173_ (.A(_02416_),
    .B(_02444_),
    .X(_02484_));
 sky130_fd_sc_hd__or2_1 _22174_ (.A(_02416_),
    .B(_02444_),
    .X(_02485_));
 sky130_fd_sc_hd__o2111a_2 _22175_ (.A1(_02413_),
    .A2(_02484_),
    .B1(_02449_),
    .C1(_02414_),
    .D1(_02485_),
    .X(_02486_));
 sky130_fd_sc_hd__nand3b_1 _22176_ (.A_N(_02444_),
    .B(_02412_),
    .C(_02408_),
    .Y(_02487_));
 sky130_fd_sc_hd__xor2_1 _22177_ (.A(_02406_),
    .B(_02407_),
    .X(_02488_));
 sky130_fd_sc_hd__a31oi_1 _22178_ (.A1(_02164_),
    .A2(_02318_),
    .A3(_02321_),
    .B1(_02412_),
    .Y(_02489_));
 sky130_fd_sc_hd__or4_4 _22179_ (.A(_02416_),
    .B(_02444_),
    .C(_02488_),
    .D(_02489_),
    .X(_02490_));
 sky130_fd_sc_hd__nand3_1 _22180_ (.A(_02416_),
    .B(_02444_),
    .C(_02413_),
    .Y(_02491_));
 sky130_fd_sc_hd__o211ai_4 _22181_ (.A1(_02449_),
    .A2(_02487_),
    .B1(_02491_),
    .C1(_02490_),
    .Y(_02492_));
 sky130_fd_sc_hd__nor2b_2 _22182_ (.A(_02406_),
    .B_N(_02407_),
    .Y(_02493_));
 sky130_fd_sc_hd__xor2_2 _22183_ (.A(_02432_),
    .B(_02442_),
    .X(_02494_));
 sky130_fd_sc_hd__o32ai_4 _22184_ (.A1(net908),
    .A2(_02305_),
    .A3(_02422_),
    .B1(_02432_),
    .B2(_02442_),
    .Y(_02495_));
 sky130_fd_sc_hd__a21oi_2 _22185_ (.A1(net1297),
    .A2(_02494_),
    .B1(_02495_),
    .Y(_02496_));
 sky130_fd_sc_hd__maj3_2 _22186_ (.A(_02403_),
    .B(_02404_),
    .C(_02405_),
    .X(_02497_));
 sky130_fd_sc_hd__mux2i_2 _22187_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[56] ),
    .A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[40] ),
    .S(net315),
    .Y(_02498_));
 sky130_fd_sc_hd__o22ai_4 _22188_ (.A1(_10343_),
    .A2(_01712_),
    .B1(_02498_),
    .B2(_08280_),
    .Y(_02499_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_362 ();
 sky130_fd_sc_hd__nor2_1 _22190_ (.A(_01982_),
    .B(net1028),
    .Y(_02501_));
 sky130_fd_sc_hd__nand3_4 _22191_ (.A(net1001),
    .B(_09183_),
    .C(_01968_),
    .Y(_02502_));
 sky130_fd_sc_hd__nand4_4 _22192_ (.A(_10349_),
    .B(_10357_),
    .C(_10364_),
    .D(_01720_),
    .Y(_02503_));
 sky130_fd_sc_hd__and2_4 _22193_ (.A(net1035),
    .B(_02503_),
    .X(_02504_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_361 ();
 sky130_fd_sc_hd__nor2_4 _22195_ (.A(net948),
    .B(_02504_),
    .Y(_02506_));
 sky130_fd_sc_hd__xnor3_1 _22196_ (.A(_02499_),
    .B(_02501_),
    .C(_02506_),
    .X(_02507_));
 sky130_fd_sc_hd__a21oi_1 _22197_ (.A1(_02400_),
    .A2(_02402_),
    .B1(_02397_),
    .Y(_02508_));
 sky130_fd_sc_hd__o21bai_2 _22198_ (.A1(_02400_),
    .A2(_02402_),
    .B1_N(_02508_),
    .Y(_02509_));
 sky130_fd_sc_hd__maj3_1 _22199_ (.A(_02438_),
    .B(_02439_),
    .C(_02441_),
    .X(_02510_));
 sky130_fd_sc_hd__xor3_2 _22200_ (.A(_02507_),
    .B(_02509_),
    .C(_02510_),
    .X(_02511_));
 sky130_fd_sc_hd__xnor2_4 _22201_ (.A(_02497_),
    .B(_02511_),
    .Y(_02512_));
 sky130_fd_sc_hd__mux2_8 _22202_ (.A0(_09217_),
    .A1(_10392_),
    .S(net322),
    .X(_02513_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_359 ();
 sky130_fd_sc_hd__nor2_1 _22205_ (.A(net1155),
    .B(_02513_),
    .Y(_02516_));
 sky130_fd_sc_hd__nor2_1 _22206_ (.A(_02010_),
    .B(_02331_),
    .Y(_02517_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_358 ();
 sky130_fd_sc_hd__nor2_2 _22208_ (.A(_02292_),
    .B(_02080_),
    .Y(_02519_));
 sky130_fd_sc_hd__nor2_1 _22209_ (.A(_02088_),
    .B(_02150_),
    .Y(_02520_));
 sky130_fd_sc_hd__xnor3_2 _22210_ (.A(_02517_),
    .B(_02519_),
    .C(_02520_),
    .X(_02521_));
 sky130_fd_sc_hd__o22ai_1 _22211_ (.A1(net1172),
    .A2(net906),
    .B1(_02426_),
    .B2(_01725_),
    .Y(_02522_));
 sky130_fd_sc_hd__nor4_1 _22212_ (.A(_01725_),
    .B(_01972_),
    .C(net906),
    .D(_02426_),
    .Y(_02523_));
 sky130_fd_sc_hd__a21oi_2 _22213_ (.A1(_02423_),
    .A2(_02522_),
    .B1(_02523_),
    .Y(_02524_));
 sky130_fd_sc_hd__nor2_4 _22214_ (.A(net788),
    .B(_02426_),
    .Y(_02525_));
 sky130_fd_sc_hd__nor2_1 _22215_ (.A(_01992_),
    .B(_02308_),
    .Y(_02526_));
 sky130_fd_sc_hd__nor2_1 _22216_ (.A(_01972_),
    .B(_02289_),
    .Y(_02527_));
 sky130_fd_sc_hd__xnor3_2 _22217_ (.A(_02527_),
    .B(_02526_),
    .C(_02525_),
    .X(_02528_));
 sky130_fd_sc_hd__xor2_2 _22218_ (.A(_02524_),
    .B(_02528_),
    .X(_02529_));
 sky130_fd_sc_hd__xnor3_2 _22219_ (.A(_02516_),
    .B(_02521_),
    .C(_02529_),
    .X(_02530_));
 sky130_fd_sc_hd__xnor2_4 _22220_ (.A(_02530_),
    .B(_02512_),
    .Y(_02531_));
 sky130_fd_sc_hd__xnor3_4 _22221_ (.A(_02493_),
    .B(_02496_),
    .C(_02531_),
    .X(_02532_));
 sky130_fd_sc_hd__o21ai_2 _22222_ (.A1(_02486_),
    .A2(_02492_),
    .B1(_02532_),
    .Y(_02533_));
 sky130_fd_sc_hd__or3_1 _22223_ (.A(net1005),
    .B(_02486_),
    .C(_02492_),
    .X(_02534_));
 sky130_fd_sc_hd__nor2_1 _22224_ (.A(_02390_),
    .B(_02450_),
    .Y(_02535_));
 sky130_fd_sc_hd__a21oi_1 _22225_ (.A1(_02533_),
    .A2(_02534_),
    .B1(_02535_),
    .Y(_02536_));
 sky130_fd_sc_hd__nor3_4 _22226_ (.A(_02532_),
    .B(_02486_),
    .C(_02492_),
    .Y(_02537_));
 sky130_fd_sc_hd__nor4b_4 _22227_ (.A(_02450_),
    .B(_02537_),
    .C(_02390_),
    .D_N(_02533_),
    .Y(_02538_));
 sky130_fd_sc_hd__nor2_2 _22228_ (.A(_02536_),
    .B(_02538_),
    .Y(_02539_));
 sky130_fd_sc_hd__mux2i_4 _22229_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[40] ),
    .A1(_02539_),
    .S(_02169_),
    .Y(_02540_));
 sky130_fd_sc_hd__nand2_1 _22230_ (.A(net442),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[40] ),
    .Y(_02541_));
 sky130_fd_sc_hd__o211ai_4 _22231_ (.A1(net442),
    .A2(_02540_),
    .B1(_02541_),
    .C1(net312),
    .Y(_02542_));
 sky130_fd_sc_hd__o21ai_2 _22232_ (.A1(_08272_),
    .A2(_02483_),
    .B1(_02542_),
    .Y(_02543_));
 sky130_fd_sc_hd__mux4_1 _22233_ (.A0(net57),
    .A1(net34),
    .A2(net43),
    .A3(net27),
    .S0(\load_store_unit_i.rdata_offset_q[0] ),
    .S1(\load_store_unit_i.rdata_offset_q[1] ),
    .X(_02544_));
 sky130_fd_sc_hd__mux4_1 _22234_ (.A0(net57),
    .A1(\load_store_unit_i.rdata_q[16] ),
    .A2(\load_store_unit_i.rdata_q[24] ),
    .A3(net27),
    .S0(\load_store_unit_i.rdata_offset_q[0] ),
    .S1(\load_store_unit_i.rdata_offset_q[1] ),
    .X(_02545_));
 sky130_fd_sc_hd__o311a_1 _22235_ (.A1(\load_store_unit_i.rdata_offset_q[0] ),
    .A2(\load_store_unit_i.rdata_offset_q[1] ),
    .A3(net56),
    .B1(\load_store_unit_i.data_sign_ext_q ),
    .C1(\load_store_unit_i.data_type_q[1] ),
    .X(_02546_));
 sky130_fd_sc_hd__mux2i_1 _22236_ (.A0(net33),
    .A1(net51),
    .S(\load_store_unit_i.rdata_offset_q[1] ),
    .Y(_02547_));
 sky130_fd_sc_hd__nand2_1 _22237_ (.A(\load_store_unit_i.rdata_offset_q[0] ),
    .B(_02547_),
    .Y(_02548_));
 sky130_fd_sc_hd__o311a_4 _22238_ (.A1(\load_store_unit_i.rdata_offset_q[0] ),
    .A2(_01682_),
    .A3(net42),
    .B1(_02546_),
    .C1(_02548_),
    .X(_02549_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_357 ();
 sky130_fd_sc_hd__a221o_1 _22240_ (.A1(\load_store_unit_i.data_type_q[2] ),
    .A2(_02544_),
    .B1(_02545_),
    .B2(_01674_),
    .C1(_02549_),
    .X(_02551_));
 sky130_fd_sc_hd__nor2_1 _22241_ (.A(net266),
    .B(_02551_),
    .Y(_02552_));
 sky130_fd_sc_hd__a31oi_4 _22242_ (.A1(_11955_),
    .A2(net265),
    .A3(_02543_),
    .B1(_02552_),
    .Y(_02553_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_356 ();
 sky130_fd_sc_hd__nand2_1 _22244_ (.A(_02119_),
    .B(_02553_),
    .Y(_02555_));
 sky130_fd_sc_hd__nand2_1 _22245_ (.A(\gen_regfile_ff.register_file_i.rf_reg[136] ),
    .B(_02123_),
    .Y(_02556_));
 sky130_fd_sc_hd__nand2_1 _22246_ (.A(_02555_),
    .B(_02556_),
    .Y(_00519_));
 sky130_fd_sc_hd__nand2_1 _22247_ (.A(_11971_),
    .B(_01665_),
    .Y(_02557_));
 sky130_fd_sc_hd__xnor2_4 _22248_ (.A(net974),
    .B(_01742_),
    .Y(_02558_));
 sky130_fd_sc_hd__nand2_1 _22249_ (.A(_01756_),
    .B(_02558_),
    .Y(_02559_));
 sky130_fd_sc_hd__nand2_1 _22250_ (.A(_01743_),
    .B(_02261_),
    .Y(_02560_));
 sky130_fd_sc_hd__nand2_1 _22251_ (.A(_02559_),
    .B(_02560_),
    .Y(_02561_));
 sky130_fd_sc_hd__mux2i_4 _22252_ (.A0(_02180_),
    .A1(_02209_),
    .S(_01758_),
    .Y(_02562_));
 sky130_fd_sc_hd__nor2_1 _22253_ (.A(_01758_),
    .B(_02204_),
    .Y(_02563_));
 sky130_fd_sc_hd__a21oi_2 _22254_ (.A1(_01758_),
    .A2(_02197_),
    .B1(_02563_),
    .Y(_02564_));
 sky130_fd_sc_hd__mux2i_4 _22255_ (.A0(_02562_),
    .A1(_02564_),
    .S(_01738_),
    .Y(_02565_));
 sky130_fd_sc_hd__nor2_1 _22256_ (.A(_01743_),
    .B(_02275_),
    .Y(_02566_));
 sky130_fd_sc_hd__a21oi_1 _22257_ (.A1(_01743_),
    .A2(_02565_),
    .B1(_02566_),
    .Y(_02567_));
 sky130_fd_sc_hd__nand2_1 _22258_ (.A(_01773_),
    .B(_02567_),
    .Y(_02568_));
 sky130_fd_sc_hd__o21ai_0 _22259_ (.A1(_01773_),
    .A2(_02561_),
    .B1(_02568_),
    .Y(_02569_));
 sky130_fd_sc_hd__nand3_1 _22260_ (.A(_09261_),
    .B(_09290_),
    .C(_02228_),
    .Y(_02570_));
 sky130_fd_sc_hd__o21ai_0 _22261_ (.A1(_09261_),
    .A2(_01902_),
    .B1(_02570_),
    .Y(_02571_));
 sky130_fd_sc_hd__a21oi_1 _22262_ (.A1(_09261_),
    .A2(_02233_),
    .B1(_09290_),
    .Y(_02572_));
 sky130_fd_sc_hd__a21oi_1 _22263_ (.A1(_02225_),
    .A2(_02571_),
    .B1(_02572_),
    .Y(_02573_));
 sky130_fd_sc_hd__a221oi_2 _22264_ (.A1(net180),
    .A2(_01929_),
    .B1(_02569_),
    .B2(_01734_),
    .C1(_02573_),
    .Y(_02574_));
 sky130_fd_sc_hd__o211ai_1 _22265_ (.A1(_02413_),
    .A2(_02484_),
    .B1(_02485_),
    .C1(_02414_),
    .Y(_02575_));
 sky130_fd_sc_hd__or3_1 _22266_ (.A(_02416_),
    .B(_02444_),
    .C(_02414_),
    .X(_02576_));
 sky130_fd_sc_hd__nand2_1 _22267_ (.A(_02575_),
    .B(_02576_),
    .Y(_02577_));
 sky130_fd_sc_hd__xnor2_1 _22268_ (.A(net1005),
    .B(_02577_),
    .Y(_02578_));
 sky130_fd_sc_hd__maj3_1 _22269_ (.A(_02390_),
    .B(_02446_),
    .C(_02449_),
    .X(_02579_));
 sky130_fd_sc_hd__nor2_2 _22270_ (.A(_02578_),
    .B(_02579_),
    .Y(_02580_));
 sky130_fd_sc_hd__inv_1 _22271_ (.A(_02575_),
    .Y(_02581_));
 sky130_fd_sc_hd__o21ai_2 _22272_ (.A1(net1005),
    .A2(_02581_),
    .B1(_02576_),
    .Y(_02582_));
 sky130_fd_sc_hd__inv_1 _22273_ (.A(_02511_),
    .Y(_02583_));
 sky130_fd_sc_hd__nand2_1 _22274_ (.A(_02497_),
    .B(_02583_),
    .Y(_02584_));
 sky130_fd_sc_hd__maj3_2 _22275_ (.A(_02499_),
    .B(_02501_),
    .C(_02506_),
    .X(_02585_));
 sky130_fd_sc_hd__or4_4 _22276_ (.A(_09267_),
    .B(_09272_),
    .C(_09282_),
    .D(_01720_),
    .X(_02586_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_355 ();
 sky130_fd_sc_hd__nand4_4 _22278_ (.A(_10283_),
    .B(_10291_),
    .C(_10298_),
    .D(_01720_),
    .Y(_02588_));
 sky130_fd_sc_hd__nand2_2 _22279_ (.A(_02586_),
    .B(_02588_),
    .Y(_02589_));
 sky130_fd_sc_hd__nand2_1 _22280_ (.A(_02032_),
    .B(_02589_),
    .Y(_02590_));
 sky130_fd_sc_hd__mux2i_2 _22281_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[57] ),
    .A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[41] ),
    .S(net315),
    .Y(_02591_));
 sky130_fd_sc_hd__nand2_1 _22282_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[57] ),
    .B(net322),
    .Y(_02592_));
 sky130_fd_sc_hd__o21ai_4 _22283_ (.A1(_08280_),
    .A2(_02591_),
    .B1(_02592_),
    .Y(_02593_));
 sky130_fd_sc_hd__a221oi_4 _22284_ (.A1(net658),
    .A2(_01712_),
    .B1(_02503_),
    .B2(net1035),
    .C1(net780),
    .Y(_02594_));
 sky130_fd_sc_hd__xor2_1 _22285_ (.A(_02593_),
    .B(_02594_),
    .X(_02595_));
 sky130_fd_sc_hd__xnor2_1 _22286_ (.A(_02590_),
    .B(_02595_),
    .Y(_02596_));
 sky130_fd_sc_hd__maj3_1 _22287_ (.A(_02517_),
    .B(_02519_),
    .C(_02520_),
    .X(_02597_));
 sky130_fd_sc_hd__xor2_1 _22288_ (.A(_02597_),
    .B(_02596_),
    .X(_02598_));
 sky130_fd_sc_hd__xnor2_2 _22289_ (.A(_02598_),
    .B(_02585_),
    .Y(_02599_));
 sky130_fd_sc_hd__maj3_2 _22290_ (.A(_02507_),
    .B(_02509_),
    .C(_02510_),
    .X(_02600_));
 sky130_fd_sc_hd__xor2_2 _22291_ (.A(_02600_),
    .B(_02599_),
    .X(_02601_));
 sky130_fd_sc_hd__xor2_2 _22292_ (.A(_02584_),
    .B(_02601_),
    .X(_02602_));
 sky130_fd_sc_hd__xnor2_1 _22293_ (.A(_02521_),
    .B(_02529_),
    .Y(_02603_));
 sky130_fd_sc_hd__maj3_2 _22294_ (.A(_02495_),
    .B(_02516_),
    .C(_02603_),
    .X(_02604_));
 sky130_fd_sc_hd__o22ai_1 _22295_ (.A1(_01992_),
    .A2(_02308_),
    .B1(_02289_),
    .B2(net1172),
    .Y(_02605_));
 sky130_fd_sc_hd__nor4_1 _22296_ (.A(_01972_),
    .B(net1050),
    .C(_02308_),
    .D(_02289_),
    .Y(_02606_));
 sky130_fd_sc_hd__a21oi_1 _22297_ (.A1(net1219),
    .A2(_02605_),
    .B1(_02606_),
    .Y(_02607_));
 sky130_fd_sc_hd__a211oi_2 _22298_ (.A1(net306),
    .A2(net321),
    .B1(net735),
    .C1(net1027),
    .Y(_02608_));
 sky130_fd_sc_hd__a211oi_2 _22299_ (.A1(net479),
    .A2(net320),
    .B1(_02061_),
    .C1(_02150_),
    .Y(_02609_));
 sky130_fd_sc_hd__a211oi_1 _22300_ (.A1(net304),
    .A2(net321),
    .B1(_02003_),
    .C1(_02331_),
    .Y(_02610_));
 sky130_fd_sc_hd__xnor2_1 _22301_ (.A(_02609_),
    .B(_02610_),
    .Y(_02611_));
 sky130_fd_sc_hd__xor2_1 _22302_ (.A(_02608_),
    .B(_02611_),
    .X(_02612_));
 sky130_fd_sc_hd__a211o_1 _22303_ (.A1(_01966_),
    .A2(_01970_),
    .B1(_02417_),
    .C1(_02419_),
    .X(_02613_));
 sky130_fd_sc_hd__o211ai_2 _22304_ (.A1(net914),
    .A2(net321),
    .B1(_02440_),
    .C1(_02307_),
    .Y(_02614_));
 sky130_fd_sc_hd__o211ai_4 _22305_ (.A1(net1057),
    .A2(_01991_),
    .B1(_02287_),
    .C1(_02288_),
    .Y(_02615_));
 sky130_fd_sc_hd__xor3_1 _22306_ (.A(_02615_),
    .B(_02614_),
    .C(_02613_),
    .X(_02616_));
 sky130_fd_sc_hd__xor3_4 _22307_ (.A(_02616_),
    .B(_02612_),
    .C(_02607_),
    .X(_02617_));
 sky130_fd_sc_hd__maj3_2 _22308_ (.A(_02524_),
    .B(_02528_),
    .C(_02521_),
    .X(_02618_));
 sky130_fd_sc_hd__and4_4 _22309_ (.A(_09240_),
    .B(_09245_),
    .C(_09252_),
    .D(_09259_),
    .X(_02619_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_354 ();
 sky130_fd_sc_hd__and4b_4 _22311_ (.A_N(_10311_),
    .B(_10318_),
    .C(_10331_),
    .D(net321),
    .X(_02621_));
 sky130_fd_sc_hd__a21o_4 _22312_ (.A1(_02619_),
    .A2(_01712_),
    .B1(_02621_),
    .X(_02622_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_353 ();
 sky130_fd_sc_hd__nor2_1 _22314_ (.A(net1155),
    .B(net1194),
    .Y(_02624_));
 sky130_fd_sc_hd__nor2_1 _22315_ (.A(net789),
    .B(_02513_),
    .Y(_02625_));
 sky130_fd_sc_hd__xor2_1 _22316_ (.A(_02624_),
    .B(_02625_),
    .X(_02626_));
 sky130_fd_sc_hd__xnor2_2 _22317_ (.A(_02626_),
    .B(_02618_),
    .Y(_02627_));
 sky130_fd_sc_hd__xnor2_2 _22318_ (.A(_02617_),
    .B(_02627_),
    .Y(_02628_));
 sky130_fd_sc_hd__xnor2_2 _22319_ (.A(_02604_),
    .B(_02628_),
    .Y(_02629_));
 sky130_fd_sc_hd__xnor2_2 _22320_ (.A(_02629_),
    .B(_02602_),
    .Y(_02630_));
 sky130_fd_sc_hd__nand2_1 _22321_ (.A(_02435_),
    .B(_02494_),
    .Y(_02631_));
 sky130_fd_sc_hd__xnor2_2 _22322_ (.A(_02495_),
    .B(_02530_),
    .Y(_02632_));
 sky130_fd_sc_hd__nand2_1 _22323_ (.A(_02631_),
    .B(_02632_),
    .Y(_02633_));
 sky130_fd_sc_hd__a31oi_1 _22324_ (.A1(_02435_),
    .A2(_02494_),
    .A3(_02530_),
    .B1(_02512_),
    .Y(_02634_));
 sky130_fd_sc_hd__a21oi_2 _22325_ (.A1(_02631_),
    .A2(_02632_),
    .B1(_02634_),
    .Y(_02635_));
 sky130_fd_sc_hd__and2_0 _22326_ (.A(_02493_),
    .B(_02512_),
    .X(_02636_));
 sky130_fd_sc_hd__nand4_2 _22327_ (.A(_02435_),
    .B(_02494_),
    .C(_02530_),
    .D(_02636_),
    .Y(_02637_));
 sky130_fd_sc_hd__o221ai_4 _22328_ (.A1(net959),
    .A2(_02633_),
    .B1(_02635_),
    .B2(_02493_),
    .C1(_02637_),
    .Y(_02638_));
 sky130_fd_sc_hd__xor2_4 _22329_ (.A(_02638_),
    .B(_02630_),
    .X(_02639_));
 sky130_fd_sc_hd__xor2_2 _22330_ (.A(_02582_),
    .B(_02639_),
    .X(_02640_));
 sky130_fd_sc_hd__xnor2_4 _22331_ (.A(_02580_),
    .B(_02640_),
    .Y(_02641_));
 sky130_fd_sc_hd__nor2_1 _22332_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[41] ),
    .B(_02169_),
    .Y(_02642_));
 sky130_fd_sc_hd__a211oi_4 _22333_ (.A1(_02169_),
    .A2(_02641_),
    .B1(_02642_),
    .C1(_13335_),
    .Y(_02643_));
 sky130_fd_sc_hd__a211oi_4 _22334_ (.A1(net442),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[41] ),
    .B1(net739),
    .C1(_02643_),
    .Y(_02644_));
 sky130_fd_sc_hd__a21oi_2 _22335_ (.A1(_08290_),
    .A2(_02574_),
    .B1(_02644_),
    .Y(_02645_));
 sky130_fd_sc_hd__or3_4 _22336_ (.A(_11197_),
    .B(_12128_),
    .C(_01664_),
    .X(_02646_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_350 ();
 sky130_fd_sc_hd__mux4_1 _22340_ (.A0(net58),
    .A1(net35),
    .A2(net44),
    .A3(net38),
    .S0(\load_store_unit_i.rdata_offset_q[0] ),
    .S1(\load_store_unit_i.rdata_offset_q[1] ),
    .X(_02650_));
 sky130_fd_sc_hd__mux4_1 _22341_ (.A0(net58),
    .A1(\load_store_unit_i.rdata_q[17] ),
    .A2(\load_store_unit_i.rdata_q[25] ),
    .A3(net38),
    .S0(\load_store_unit_i.rdata_offset_q[0] ),
    .S1(\load_store_unit_i.rdata_offset_q[1] ),
    .X(_02651_));
 sky130_fd_sc_hd__a221oi_4 _22342_ (.A1(\load_store_unit_i.data_type_q[2] ),
    .A2(_02650_),
    .B1(_02651_),
    .B2(_01674_),
    .C1(_02549_),
    .Y(_02652_));
 sky130_fd_sc_hd__a2bb2oi_4 _22343_ (.A1_N(_02557_),
    .A2_N(_02645_),
    .B1(_02646_),
    .B2(_02652_),
    .Y(_02653_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_349 ();
 sky130_fd_sc_hd__nand2_1 _22345_ (.A(_02119_),
    .B(_02653_),
    .Y(_02655_));
 sky130_fd_sc_hd__nand2_1 _22346_ (.A(\gen_regfile_ff.register_file_i.rf_reg[137] ),
    .B(_02123_),
    .Y(_02656_));
 sky130_fd_sc_hd__nand2_1 _22347_ (.A(_02655_),
    .B(_02656_),
    .Y(_00520_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_348 ();
 sky130_fd_sc_hd__nand2_1 _22349_ (.A(_01735_),
    .B(_02558_),
    .Y(_02658_));
 sky130_fd_sc_hd__o21a_1 _22350_ (.A1(_02558_),
    .A2(_02189_),
    .B1(_02658_),
    .X(_02659_));
 sky130_fd_sc_hd__mux2i_2 _22351_ (.A0(_02256_),
    .A1(_02263_),
    .S(_01758_),
    .Y(_02660_));
 sky130_fd_sc_hd__mux2i_2 _22352_ (.A0(_02262_),
    .A1(_02265_),
    .S(_01758_),
    .Y(_02661_));
 sky130_fd_sc_hd__mux4_1 _22353_ (.A0(_01735_),
    .A1(_02220_),
    .A2(_02660_),
    .A3(_02661_),
    .S0(_01738_),
    .S1(_01743_),
    .X(_02662_));
 sky130_fd_sc_hd__nand2_1 _22354_ (.A(_01773_),
    .B(_02662_),
    .Y(_02663_));
 sky130_fd_sc_hd__o21ai_2 _22355_ (.A1(_01773_),
    .A2(_02659_),
    .B1(_02663_),
    .Y(_02664_));
 sky130_fd_sc_hd__nand3_1 _22356_ (.A(_09385_),
    .B(_10852_),
    .C(_02228_),
    .Y(_02665_));
 sky130_fd_sc_hd__o21ai_0 _22357_ (.A1(_10852_),
    .A2(_01902_),
    .B1(_02665_),
    .Y(_02666_));
 sky130_fd_sc_hd__a21oi_1 _22358_ (.A1(_10852_),
    .A2(_02233_),
    .B1(_09385_),
    .Y(_02667_));
 sky130_fd_sc_hd__a21oi_1 _22359_ (.A1(_02225_),
    .A2(_02666_),
    .B1(_02667_),
    .Y(_02668_));
 sky130_fd_sc_hd__a221o_1 _22360_ (.A1(net151),
    .A2(_01929_),
    .B1(_02664_),
    .B2(_01734_),
    .C1(_02668_),
    .X(_02669_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_347 ();
 sky130_fd_sc_hd__nand2_1 _22362_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[42] ),
    .B(_01698_),
    .Y(_02671_));
 sky130_fd_sc_hd__nor2_1 _22363_ (.A(_02582_),
    .B(_02639_),
    .Y(_02672_));
 sky130_fd_sc_hd__o21ai_1 _22364_ (.A1(_02532_),
    .A2(_02484_),
    .B1(_02413_),
    .Y(_02673_));
 sky130_fd_sc_hd__nand2_1 _22365_ (.A(_02532_),
    .B(_02485_),
    .Y(_02674_));
 sky130_fd_sc_hd__a22o_1 _22366_ (.A1(_02408_),
    .A2(_02412_),
    .B1(_02674_),
    .B2(_02673_),
    .X(_02675_));
 sky130_fd_sc_hd__o211ai_2 _22367_ (.A1(_02532_),
    .A2(_02581_),
    .B1(_02576_),
    .C1(_02449_),
    .Y(_02676_));
 sky130_fd_sc_hd__nand2_1 _22368_ (.A(net1005),
    .B(_02484_),
    .Y(_02677_));
 sky130_fd_sc_hd__a41oi_4 _22369_ (.A1(_02675_),
    .A2(_02639_),
    .A3(_02676_),
    .A4(_02677_),
    .B1(_02538_),
    .Y(_02678_));
 sky130_fd_sc_hd__nor2_1 _22370_ (.A(_02672_),
    .B(_02678_),
    .Y(_02679_));
 sky130_fd_sc_hd__a211oi_1 _22371_ (.A1(_02493_),
    .A2(_02633_),
    .B1(_02635_),
    .C1(_02636_),
    .Y(_02680_));
 sky130_fd_sc_hd__o21ai_2 _22372_ (.A1(net1275),
    .A2(_02680_),
    .B1(_02637_),
    .Y(_02681_));
 sky130_fd_sc_hd__inv_1 _22373_ (.A(_02584_),
    .Y(_02682_));
 sky130_fd_sc_hd__maj3_2 _22374_ (.A(_02604_),
    .B(_02601_),
    .C(_02628_),
    .X(_02683_));
 sky130_fd_sc_hd__nand3_1 _22375_ (.A(_02497_),
    .B(_02583_),
    .C(_02604_),
    .Y(_02684_));
 sky130_fd_sc_hd__nand2_1 _22376_ (.A(_02601_),
    .B(_02628_),
    .Y(_02685_));
 sky130_fd_sc_hd__or3_1 _22377_ (.A(_02604_),
    .B(_02601_),
    .C(_02628_),
    .X(_02686_));
 sky130_fd_sc_hd__o221ai_2 _22378_ (.A1(_02683_),
    .A2(_02682_),
    .B1(_02684_),
    .B2(_02685_),
    .C1(_02686_),
    .Y(_02687_));
 sky130_fd_sc_hd__nand3_1 _22379_ (.A(_10444_),
    .B(_10447_),
    .C(_02072_),
    .Y(_02688_));
 sky130_fd_sc_hd__nand3_2 _22380_ (.A(_09364_),
    .B(_09368_),
    .C(_02074_),
    .Y(_02689_));
 sky130_fd_sc_hd__o311ai_4 _22381_ (.A1(net1152),
    .A2(_10450_),
    .A3(_10452_),
    .B1(_10455_),
    .C1(_02076_),
    .Y(_02690_));
 sky130_fd_sc_hd__o311ai_4 _22382_ (.A1(net1152),
    .A2(_09372_),
    .A3(_09374_),
    .B1(_09378_),
    .C1(_02078_),
    .Y(_02691_));
 sky130_fd_sc_hd__nand4_4 _22383_ (.A(_02688_),
    .B(_02689_),
    .C(_02690_),
    .D(_02691_),
    .Y(_02692_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_346 ();
 sky130_fd_sc_hd__a221oi_2 _22385_ (.A1(_09856_),
    .A2(net321),
    .B1(_02029_),
    .B2(_02030_),
    .C1(_02692_),
    .Y(_02694_));
 sky130_fd_sc_hd__mux2i_2 _22386_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[58] ),
    .A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[42] ),
    .S(net315),
    .Y(_02695_));
 sky130_fd_sc_hd__nand2_1 _22387_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[58] ),
    .B(net322),
    .Y(_02696_));
 sky130_fd_sc_hd__o21ai_4 _22388_ (.A1(_08280_),
    .A2(_02695_),
    .B1(_02696_),
    .Y(_02697_));
 sky130_fd_sc_hd__a221oi_2 _22389_ (.A1(_08995_),
    .A2(net320),
    .B1(_02586_),
    .B2(_02588_),
    .C1(net1268),
    .Y(_02698_));
 sky130_fd_sc_hd__xor2_1 _22390_ (.A(_02697_),
    .B(_02698_),
    .X(_02699_));
 sky130_fd_sc_hd__xnor2_1 _22391_ (.A(_02694_),
    .B(_02699_),
    .Y(_02700_));
 sky130_fd_sc_hd__a21oi_1 _22392_ (.A1(_02608_),
    .A2(_02609_),
    .B1(_02610_),
    .Y(_02701_));
 sky130_fd_sc_hd__o21bai_1 _22393_ (.A1(_02608_),
    .A2(_02609_),
    .B1_N(_02701_),
    .Y(_02702_));
 sky130_fd_sc_hd__nand2_1 _22394_ (.A(_02593_),
    .B(_02594_),
    .Y(_02703_));
 sky130_fd_sc_hd__nor2_1 _22395_ (.A(_02593_),
    .B(_02594_),
    .Y(_02704_));
 sky130_fd_sc_hd__a21o_1 _22396_ (.A1(_02590_),
    .A2(_02703_),
    .B1(_02704_),
    .X(_02705_));
 sky130_fd_sc_hd__xnor3_1 _22397_ (.A(_02700_),
    .B(_02702_),
    .C(_02705_),
    .X(_02706_));
 sky130_fd_sc_hd__maj3_2 _22398_ (.A(_02597_),
    .B(_02596_),
    .C(_02585_),
    .X(_02707_));
 sky130_fd_sc_hd__xnor2_2 _22399_ (.A(_02706_),
    .B(_02707_),
    .Y(_02708_));
 sky130_fd_sc_hd__nor3_2 _22400_ (.A(net1159),
    .B(_02600_),
    .C(_02708_),
    .Y(_02709_));
 sky130_fd_sc_hd__o21ai_1 _22401_ (.A1(net1159),
    .A2(_02600_),
    .B1(_02708_),
    .Y(_02710_));
 sky130_fd_sc_hd__nor2b_4 _22402_ (.A(_02709_),
    .B_N(_02710_),
    .Y(_02711_));
 sky130_fd_sc_hd__a211oi_1 _22403_ (.A1(_02083_),
    .A2(_02085_),
    .B1(_02417_),
    .C1(_02419_),
    .Y(_02712_));
 sky130_fd_sc_hd__a211oi_1 _22404_ (.A1(_10865_),
    .A2(net320),
    .B1(_02131_),
    .C1(_02150_),
    .Y(_02713_));
 sky130_fd_sc_hd__nor3_2 _22405_ (.A(_02080_),
    .B(_02299_),
    .C(_02300_),
    .Y(_02714_));
 sky130_fd_sc_hd__xnor3_1 _22406_ (.A(_02714_),
    .B(_02713_),
    .C(_02712_),
    .X(_02715_));
 sky130_fd_sc_hd__a211oi_1 _22407_ (.A1(net476),
    .A2(net320),
    .B1(_02061_),
    .C1(_02331_),
    .Y(_02716_));
 sky130_fd_sc_hd__a211oi_1 _22408_ (.A1(net304),
    .A2(net321),
    .B1(_02003_),
    .C1(net1027),
    .Y(_02717_));
 sky130_fd_sc_hd__a221oi_4 _22409_ (.A1(net306),
    .A2(net321),
    .B1(net1035),
    .B2(_02503_),
    .C1(net734),
    .Y(_02718_));
 sky130_fd_sc_hd__xnor3_1 _22410_ (.A(_02716_),
    .B(_02717_),
    .C(_02718_),
    .X(_02719_));
 sky130_fd_sc_hd__maj3_1 _22411_ (.A(_02613_),
    .B(_02614_),
    .C(_02615_),
    .X(_02720_));
 sky130_fd_sc_hd__xnor2_1 _22412_ (.A(_02719_),
    .B(_02720_),
    .Y(_02721_));
 sky130_fd_sc_hd__xnor2_2 _22413_ (.A(net936),
    .B(_02721_),
    .Y(_02722_));
 sky130_fd_sc_hd__and4_4 _22414_ (.A(_09392_),
    .B(net1079),
    .C(_09412_),
    .D(net320),
    .X(_02723_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_345 ();
 sky130_fd_sc_hd__and4_4 _22416_ (.A(_10416_),
    .B(net884),
    .C(_10423_),
    .D(net321),
    .X(_02725_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_344 ();
 sky130_fd_sc_hd__nor2_8 _22418_ (.A(_02723_),
    .B(_02725_),
    .Y(_02727_));
 sky130_fd_sc_hd__xnor2_1 _22419_ (.A(_02158_),
    .B(_02727_),
    .Y(_02728_));
 sky130_fd_sc_hd__nor2_1 _22420_ (.A(net790),
    .B(net1194),
    .Y(_02729_));
 sky130_fd_sc_hd__or2_4 _22421_ (.A(_02725_),
    .B(_02723_),
    .X(_02730_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_343 ();
 sky130_fd_sc_hd__nor2_1 _22423_ (.A(net1155),
    .B(net1213),
    .Y(_02732_));
 sky130_fd_sc_hd__nor2_1 _22424_ (.A(net1172),
    .B(_02513_),
    .Y(_02733_));
 sky130_fd_sc_hd__a22o_1 _22425_ (.A1(net1161),
    .A2(_02732_),
    .B1(_02733_),
    .B2(net1176),
    .X(_02734_));
 sky130_fd_sc_hd__nand2_1 _22426_ (.A(net1161),
    .B(net1158),
    .Y(_02735_));
 sky130_fd_sc_hd__o21ai_0 _22427_ (.A1(net781),
    .A2(net1161),
    .B1(net1155),
    .Y(_02736_));
 sky130_fd_sc_hd__a21oi_1 _22428_ (.A1(_02735_),
    .A2(_02736_),
    .B1(_02729_),
    .Y(_02737_));
 sky130_fd_sc_hd__a221o_1 _22429_ (.A1(_02516_),
    .A2(_02728_),
    .B1(_02729_),
    .B2(_02734_),
    .C1(_02737_),
    .X(_02738_));
 sky130_fd_sc_hd__maj3_1 _22430_ (.A(_02607_),
    .B(_02612_),
    .C(_02616_),
    .X(_02739_));
 sky130_fd_sc_hd__xnor2_1 _22431_ (.A(_02738_),
    .B(_02739_),
    .Y(_02740_));
 sky130_fd_sc_hd__xnor2_2 _22432_ (.A(_02722_),
    .B(_02740_),
    .Y(_02741_));
 sky130_fd_sc_hd__inv_1 _22433_ (.A(_02626_),
    .Y(_02742_));
 sky130_fd_sc_hd__maj3_2 _22434_ (.A(_02618_),
    .B(_02617_),
    .C(_02742_),
    .X(_02743_));
 sky130_fd_sc_hd__inv_1 _22435_ (.A(_02743_),
    .Y(_02744_));
 sky130_fd_sc_hd__xnor2_2 _22436_ (.A(_02741_),
    .B(_02744_),
    .Y(_02745_));
 sky130_fd_sc_hd__xnor2_4 _22437_ (.A(_02711_),
    .B(_02745_),
    .Y(_02746_));
 sky130_fd_sc_hd__xor2_2 _22438_ (.A(_02746_),
    .B(_02687_),
    .X(_02747_));
 sky130_fd_sc_hd__xor2_2 _22439_ (.A(_02747_),
    .B(_02681_),
    .X(_02748_));
 sky130_fd_sc_hd__nor2_1 _22440_ (.A(_02679_),
    .B(_02748_),
    .Y(_02749_));
 sky130_fd_sc_hd__nor3b_4 _22441_ (.A(_02678_),
    .B(_02672_),
    .C_N(_02748_),
    .Y(_02750_));
 sky130_fd_sc_hd__nor2_2 _22442_ (.A(_02749_),
    .B(_02750_),
    .Y(_02751_));
 sky130_fd_sc_hd__nand2_1 _22443_ (.A(_02169_),
    .B(_02751_),
    .Y(_02752_));
 sky130_fd_sc_hd__nand2_2 _22444_ (.A(_02671_),
    .B(_02752_),
    .Y(_02753_));
 sky130_fd_sc_hd__mux2i_1 _22445_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[42] ),
    .A1(_02753_),
    .S(_08100_),
    .Y(_02754_));
 sky130_fd_sc_hd__nand2_2 _22446_ (.A(net313),
    .B(_02754_),
    .Y(_02755_));
 sky130_fd_sc_hd__o21ai_2 _22447_ (.A1(_08272_),
    .A2(_02669_),
    .B1(_02755_),
    .Y(_02756_));
 sky130_fd_sc_hd__mux4_1 _22448_ (.A0(net28),
    .A1(net36),
    .A2(net45),
    .A3(net49),
    .S0(\load_store_unit_i.rdata_offset_q[0] ),
    .S1(\load_store_unit_i.rdata_offset_q[1] ),
    .X(_02757_));
 sky130_fd_sc_hd__mux4_1 _22449_ (.A0(net28),
    .A1(\load_store_unit_i.rdata_q[18] ),
    .A2(\load_store_unit_i.rdata_q[26] ),
    .A3(net49),
    .S0(\load_store_unit_i.rdata_offset_q[0] ),
    .S1(\load_store_unit_i.rdata_offset_q[1] ),
    .X(_02758_));
 sky130_fd_sc_hd__a221o_1 _22450_ (.A1(\load_store_unit_i.data_type_q[2] ),
    .A2(_02757_),
    .B1(_02758_),
    .B2(_01674_),
    .C1(_02549_),
    .X(_02759_));
 sky130_fd_sc_hd__nor2_1 _22451_ (.A(net267),
    .B(_02759_),
    .Y(_02760_));
 sky130_fd_sc_hd__a31oi_4 _22452_ (.A1(_11354_),
    .A2(_01665_),
    .A3(_02756_),
    .B1(_02760_),
    .Y(_02761_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_342 ();
 sky130_fd_sc_hd__nand2_1 _22454_ (.A(_02119_),
    .B(_02761_),
    .Y(_02763_));
 sky130_fd_sc_hd__nand2_1 _22455_ (.A(\gen_regfile_ff.register_file_i.rf_reg[138] ),
    .B(_02123_),
    .Y(_02764_));
 sky130_fd_sc_hd__nand2_1 _22456_ (.A(_02763_),
    .B(_02764_),
    .Y(_00521_));
 sky130_fd_sc_hd__mux4_1 _22457_ (.A0(net29),
    .A1(net37),
    .A2(net46),
    .A3(net52),
    .S0(\load_store_unit_i.rdata_offset_q[0] ),
    .S1(\load_store_unit_i.rdata_offset_q[1] ),
    .X(_02765_));
 sky130_fd_sc_hd__mux4_1 _22458_ (.A0(net29),
    .A1(\load_store_unit_i.rdata_q[19] ),
    .A2(\load_store_unit_i.rdata_q[27] ),
    .A3(net52),
    .S0(\load_store_unit_i.rdata_offset_q[0] ),
    .S1(\load_store_unit_i.rdata_offset_q[1] ),
    .X(_02766_));
 sky130_fd_sc_hd__a221oi_2 _22459_ (.A1(\load_store_unit_i.data_type_q[2] ),
    .A2(_02765_),
    .B1(_02766_),
    .B2(_01674_),
    .C1(_02549_),
    .Y(_02767_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_341 ();
 sky130_fd_sc_hd__o21ai_0 _22461_ (.A1(_02709_),
    .A2(_02744_),
    .B1(_02710_),
    .Y(_02769_));
 sky130_fd_sc_hd__or4_1 _22462_ (.A(net1159),
    .B(_02600_),
    .C(_02708_),
    .D(_02743_),
    .X(_02770_));
 sky130_fd_sc_hd__o22ai_1 _22463_ (.A1(_02710_),
    .A2(_02744_),
    .B1(_02770_),
    .B2(_02741_),
    .Y(_02771_));
 sky130_fd_sc_hd__a21oi_1 _22464_ (.A1(_02741_),
    .A2(_02769_),
    .B1(_02771_),
    .Y(_02772_));
 sky130_fd_sc_hd__nor4_4 _22465_ (.A(_10521_),
    .B(_10514_),
    .C(_10509_),
    .D(net320),
    .Y(_02773_));
 sky130_fd_sc_hd__a21oi_4 _22466_ (.A1(net307),
    .A2(_01712_),
    .B1(net1221),
    .Y(_02774_));
 sky130_fd_sc_hd__nand2_1 _22467_ (.A(_01998_),
    .B(_02774_),
    .Y(_02775_));
 sky130_fd_sc_hd__nor2_4 _22468_ (.A(net1213),
    .B(net790),
    .Y(_02776_));
 sky130_fd_sc_hd__nor2_1 _22469_ (.A(_01992_),
    .B(_02513_),
    .Y(_02777_));
 sky130_fd_sc_hd__nor2_1 _22470_ (.A(net781),
    .B(net1194),
    .Y(_02778_));
 sky130_fd_sc_hd__xor3_2 _22471_ (.A(_02778_),
    .B(_02777_),
    .C(_02776_),
    .X(_02779_));
 sky130_fd_sc_hd__maj3_1 _22472_ (.A(_02729_),
    .B(_02732_),
    .C(_02733_),
    .X(_02780_));
 sky130_fd_sc_hd__xor3_1 _22473_ (.A(_02775_),
    .B(_02779_),
    .C(_02780_),
    .X(_02781_));
 sky130_fd_sc_hd__maj3_1 _22474_ (.A(_02715_),
    .B(_02719_),
    .C(_02720_),
    .X(_02782_));
 sky130_fd_sc_hd__nor3_1 _22475_ (.A(_02080_),
    .B(_02417_),
    .C(_02419_),
    .Y(_02783_));
 sky130_fd_sc_hd__nor3_2 _22476_ (.A(_02150_),
    .B(_02299_),
    .C(_02300_),
    .Y(_02784_));
 sky130_fd_sc_hd__a211oi_2 _22477_ (.A1(_10865_),
    .A2(net320),
    .B1(_02131_),
    .C1(_02331_),
    .Y(_02785_));
 sky130_fd_sc_hd__xnor3_1 _22478_ (.A(_02785_),
    .B(_02784_),
    .C(_02783_),
    .X(_02786_));
 sky130_fd_sc_hd__a221oi_1 _22479_ (.A1(net306),
    .A2(net322),
    .B1(_02586_),
    .B2(_02588_),
    .C1(net735),
    .Y(_02787_));
 sky130_fd_sc_hd__a211oi_1 _22480_ (.A1(net309),
    .A2(net320),
    .B1(_02061_),
    .C1(net1027),
    .Y(_02788_));
 sky130_fd_sc_hd__a221oi_4 _22481_ (.A1(net749),
    .A2(net322),
    .B1(net1035),
    .B2(_02503_),
    .C1(net1051),
    .Y(_02789_));
 sky130_fd_sc_hd__xnor3_1 _22482_ (.A(_02787_),
    .B(_02788_),
    .C(_02789_),
    .X(_02790_));
 sky130_fd_sc_hd__maj3_1 _22483_ (.A(_02712_),
    .B(_02713_),
    .C(_02714_),
    .X(_02791_));
 sky130_fd_sc_hd__xnor3_1 _22484_ (.A(_02786_),
    .B(_02790_),
    .C(_02791_),
    .X(_02792_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_339 ();
 sky130_fd_sc_hd__nor4b_1 _22487_ (.A(_02089_),
    .B(net1161),
    .C(net1173),
    .D_N(_02728_),
    .Y(_02795_));
 sky130_fd_sc_hd__xnor3_2 _22488_ (.A(_02782_),
    .B(_02792_),
    .C(_02795_),
    .X(_02796_));
 sky130_fd_sc_hd__xnor2_4 _22489_ (.A(_02796_),
    .B(_02781_),
    .Y(_02797_));
 sky130_fd_sc_hd__maj3_1 _22490_ (.A(_02722_),
    .B(_02738_),
    .C(_02739_),
    .X(_02798_));
 sky130_fd_sc_hd__nand2_2 _22491_ (.A(_02706_),
    .B(_02707_),
    .Y(_02799_));
 sky130_fd_sc_hd__mux4_4 _22492_ (.A0(_09340_),
    .A1(_09348_),
    .A2(_10484_),
    .A3(_10492_),
    .S0(_08512_),
    .S1(_01720_),
    .X(_02800_));
 sky130_fd_sc_hd__a221oi_2 _22493_ (.A1(_09856_),
    .A2(net321),
    .B1(_02029_),
    .B2(_02030_),
    .C1(_02800_),
    .Y(_02801_));
 sky130_fd_sc_hd__mux2i_2 _22494_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[59] ),
    .A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[43] ),
    .S(net315),
    .Y(_02802_));
 sky130_fd_sc_hd__nand2_1 _22495_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[59] ),
    .B(net322),
    .Y(_02803_));
 sky130_fd_sc_hd__o21ai_4 _22496_ (.A1(_08280_),
    .A2(_02802_),
    .B1(_02803_),
    .Y(_02804_));
 sky130_fd_sc_hd__a211oi_1 _22497_ (.A1(net699),
    .A2(net320),
    .B1(net1268),
    .C1(_02692_),
    .Y(_02805_));
 sky130_fd_sc_hd__xnor2_1 _22498_ (.A(_02804_),
    .B(_02805_),
    .Y(_02806_));
 sky130_fd_sc_hd__xnor2_1 _22499_ (.A(_02801_),
    .B(_02806_),
    .Y(_02807_));
 sky130_fd_sc_hd__maj3_1 _22500_ (.A(_02716_),
    .B(_02717_),
    .C(_02718_),
    .X(_02808_));
 sky130_fd_sc_hd__maj3_1 _22501_ (.A(_02697_),
    .B(_02694_),
    .C(_02698_),
    .X(_02809_));
 sky130_fd_sc_hd__xor2_1 _22502_ (.A(_02808_),
    .B(_02809_),
    .X(_02810_));
 sky130_fd_sc_hd__xnor2_1 _22503_ (.A(_02807_),
    .B(_02810_),
    .Y(_02811_));
 sky130_fd_sc_hd__maj3_1 _22504_ (.A(_02700_),
    .B(_02702_),
    .C(_02705_),
    .X(_02812_));
 sky130_fd_sc_hd__xor2_2 _22505_ (.A(_02811_),
    .B(_02812_),
    .X(_02813_));
 sky130_fd_sc_hd__xor2_1 _22506_ (.A(_02799_),
    .B(_02813_),
    .X(_02814_));
 sky130_fd_sc_hd__xnor2_1 _22507_ (.A(_02798_),
    .B(_02814_),
    .Y(_02815_));
 sky130_fd_sc_hd__xnor2_2 _22508_ (.A(net888),
    .B(_02815_),
    .Y(_02816_));
 sky130_fd_sc_hd__xor2_2 _22509_ (.A(_02772_),
    .B(_02816_),
    .X(_02817_));
 sky130_fd_sc_hd__o21ai_0 _22510_ (.A1(_02601_),
    .A2(_02628_),
    .B1(_02604_),
    .Y(_02818_));
 sky130_fd_sc_hd__nand2_1 _22511_ (.A(_02682_),
    .B(_02686_),
    .Y(_02819_));
 sky130_fd_sc_hd__a21o_1 _22512_ (.A1(_02818_),
    .A2(_02819_),
    .B1(net1267),
    .X(_02820_));
 sky130_fd_sc_hd__a21o_1 _22513_ (.A1(_02684_),
    .A2(_02746_),
    .B1(_02685_),
    .X(_02821_));
 sky130_fd_sc_hd__nand3_4 _22514_ (.A(_02817_),
    .B(_02820_),
    .C(_02821_),
    .Y(_02822_));
 sky130_fd_sc_hd__a21o_1 _22515_ (.A1(_02820_),
    .A2(_02821_),
    .B1(_02817_),
    .X(_02823_));
 sky130_fd_sc_hd__nand2_2 _22516_ (.A(_02822_),
    .B(_02823_),
    .Y(_02824_));
 sky130_fd_sc_hd__nand2_1 _22517_ (.A(_02681_),
    .B(_02747_),
    .Y(_02825_));
 sky130_fd_sc_hd__nand2b_1 _22518_ (.A_N(_02750_),
    .B(_02825_),
    .Y(_02826_));
 sky130_fd_sc_hd__xor2_4 _22519_ (.A(_02824_),
    .B(_02826_),
    .X(_02827_));
 sky130_fd_sc_hd__nor2_1 _22520_ (.A(_01698_),
    .B(_02827_),
    .Y(_02828_));
 sky130_fd_sc_hd__a21oi_2 _22521_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[43] ),
    .A2(_01698_),
    .B1(_02828_),
    .Y(_02829_));
 sky130_fd_sc_hd__nor2_1 _22522_ (.A(net442),
    .B(_02829_),
    .Y(_02830_));
 sky130_fd_sc_hd__a21oi_4 _22523_ (.A1(net442),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[43] ),
    .B1(_02830_),
    .Y(_02831_));
 sky130_fd_sc_hd__o21ai_1 _22524_ (.A1(_02558_),
    .A2(_01950_),
    .B1(_02658_),
    .Y(_02832_));
 sky130_fd_sc_hd__mux2i_1 _22525_ (.A0(_02366_),
    .A1(_02372_),
    .S(_01758_),
    .Y(_02833_));
 sky130_fd_sc_hd__nor2_1 _22526_ (.A(_01738_),
    .B(_02833_),
    .Y(_02834_));
 sky130_fd_sc_hd__mux2i_1 _22527_ (.A0(_02371_),
    .A1(_02375_),
    .S(_01758_),
    .Y(_02835_));
 sky130_fd_sc_hd__nor2_1 _22528_ (.A(_01826_),
    .B(_02835_),
    .Y(_02836_));
 sky130_fd_sc_hd__o21ai_0 _22529_ (.A1(_02834_),
    .A2(_02836_),
    .B1(_01743_),
    .Y(_02837_));
 sky130_fd_sc_hd__o21ai_0 _22530_ (.A1(_01743_),
    .A2(_01942_),
    .B1(_02837_),
    .Y(_02838_));
 sky130_fd_sc_hd__nor2_1 _22531_ (.A(_01762_),
    .B(_02838_),
    .Y(_02839_));
 sky130_fd_sc_hd__a21oi_1 _22532_ (.A1(_01762_),
    .A2(_02832_),
    .B1(_02839_),
    .Y(_02840_));
 sky130_fd_sc_hd__nor3_1 _22533_ (.A(net1139),
    .B(_09357_),
    .C(_01898_),
    .Y(_02841_));
 sky130_fd_sc_hd__a21oi_1 _22534_ (.A1(_09357_),
    .A2(_01896_),
    .B1(_02841_),
    .Y(_02842_));
 sky130_fd_sc_hd__o21ai_0 _22535_ (.A1(_09357_),
    .A2(_01903_),
    .B1(net1139),
    .Y(_02843_));
 sky130_fd_sc_hd__o21ai_0 _22536_ (.A1(_01893_),
    .A2(_02842_),
    .B1(_02843_),
    .Y(_02844_));
 sky130_fd_sc_hd__o221ai_1 _22537_ (.A1(net1590),
    .A2(_01889_),
    .B1(_02840_),
    .B2(_01761_),
    .C1(_02844_),
    .Y(_02845_));
 sky130_fd_sc_hd__nor2_1 _22538_ (.A(net1103),
    .B(_02845_),
    .Y(_02846_));
 sky130_fd_sc_hd__a21oi_2 _22539_ (.A1(net1104),
    .A2(_02831_),
    .B1(_02846_),
    .Y(_02847_));
 sky130_fd_sc_hd__nor3_2 _22540_ (.A(_11389_),
    .B(_02646_),
    .C(_02847_),
    .Y(_02848_));
 sky130_fd_sc_hd__a21oi_4 _22541_ (.A1(_02646_),
    .A2(_02767_),
    .B1(_02848_),
    .Y(_02849_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_338 ();
 sky130_fd_sc_hd__nand2_1 _22543_ (.A(_02119_),
    .B(_02849_),
    .Y(_02851_));
 sky130_fd_sc_hd__nand2_1 _22544_ (.A(\gen_regfile_ff.register_file_i.rf_reg[139] ),
    .B(_02123_),
    .Y(_02852_));
 sky130_fd_sc_hd__nand2_1 _22545_ (.A(_02851_),
    .B(_02852_),
    .Y(_00522_));
 sky130_fd_sc_hd__nand3_1 _22546_ (.A(\load_store_unit_i.rdata_offset_q[0] ),
    .B(_01682_),
    .C(net39),
    .Y(_02853_));
 sky130_fd_sc_hd__nand2_1 _22547_ (.A(net47),
    .B(_01683_),
    .Y(_02854_));
 sky130_fd_sc_hd__a221oi_1 _22548_ (.A1(_01682_),
    .A2(\load_store_unit_i.rdata_q[20] ),
    .B1(_01683_),
    .B2(\load_store_unit_i.rdata_q[28] ),
    .C1(\load_store_unit_i.data_type_q[2] ),
    .Y(_02855_));
 sky130_fd_sc_hd__a31oi_1 _22549_ (.A1(\load_store_unit_i.data_type_q[2] ),
    .A2(_02853_),
    .A3(_02854_),
    .B1(_02855_),
    .Y(_02856_));
 sky130_fd_sc_hd__a21oi_1 _22550_ (.A1(\load_store_unit_i.rdata_offset_q[1] ),
    .A2(net53),
    .B1(_02856_),
    .Y(_02857_));
 sky130_fd_sc_hd__nor2_1 _22551_ (.A(\load_store_unit_i.rdata_offset_q[0] ),
    .B(\load_store_unit_i.rdata_offset_q[1] ),
    .Y(_02858_));
 sky130_fd_sc_hd__a22oi_1 _22552_ (.A1(net30),
    .A2(_02858_),
    .B1(_02856_),
    .B2(\load_store_unit_i.rdata_offset_q[1] ),
    .Y(_02859_));
 sky130_fd_sc_hd__o21ai_0 _22553_ (.A1(_01670_),
    .A2(_02857_),
    .B1(_02859_),
    .Y(_02860_));
 sky130_fd_sc_hd__a21oi_1 _22554_ (.A1(_01688_),
    .A2(_02860_),
    .B1(_02549_),
    .Y(_02861_));
 sky130_fd_sc_hd__nor2_1 _22555_ (.A(_01826_),
    .B(_02833_),
    .Y(_02862_));
 sky130_fd_sc_hd__a21oi_1 _22556_ (.A1(_01826_),
    .A2(_01940_),
    .B1(_02862_),
    .Y(_02863_));
 sky130_fd_sc_hd__a21oi_1 _22557_ (.A1(_01743_),
    .A2(_02863_),
    .B1(_01943_),
    .Y(_02864_));
 sky130_fd_sc_hd__a21oi_1 _22558_ (.A1(_01758_),
    .A2(_01738_),
    .B1(_01756_),
    .Y(_02865_));
 sky130_fd_sc_hd__a31oi_1 _22559_ (.A1(_01758_),
    .A2(_01738_),
    .A3(_01800_),
    .B1(_02865_),
    .Y(_02866_));
 sky130_fd_sc_hd__nor2_1 _22560_ (.A(_01738_),
    .B(_01946_),
    .Y(_02867_));
 sky130_fd_sc_hd__nor2_1 _22561_ (.A(_01826_),
    .B(_01951_),
    .Y(_02868_));
 sky130_fd_sc_hd__or3_1 _22562_ (.A(_02558_),
    .B(_02867_),
    .C(_02868_),
    .X(_02869_));
 sky130_fd_sc_hd__o21ai_1 _22563_ (.A1(_01743_),
    .A2(_02866_),
    .B1(_02869_),
    .Y(_02870_));
 sky130_fd_sc_hd__nand2_1 _22564_ (.A(_01773_),
    .B(_02870_),
    .Y(_02871_));
 sky130_fd_sc_hd__o21ai_0 _22565_ (.A1(_01773_),
    .A2(_02864_),
    .B1(_02871_),
    .Y(_02872_));
 sky130_fd_sc_hd__nand3_1 _22566_ (.A(_09526_),
    .B(_09562_),
    .C(_02228_),
    .Y(_02873_));
 sky130_fd_sc_hd__o21ai_0 _22567_ (.A1(_09562_),
    .A2(_01902_),
    .B1(_02873_),
    .Y(_02874_));
 sky130_fd_sc_hd__a21oi_1 _22568_ (.A1(_09562_),
    .A2(_02233_),
    .B1(_09526_),
    .Y(_02875_));
 sky130_fd_sc_hd__a21oi_1 _22569_ (.A1(_02225_),
    .A2(_02874_),
    .B1(_02875_),
    .Y(_02876_));
 sky130_fd_sc_hd__a221oi_1 _22570_ (.A1(net153),
    .A2(_01929_),
    .B1(_02872_),
    .B2(_01734_),
    .C1(_02876_),
    .Y(_02877_));
 sky130_fd_sc_hd__nand2_1 _22571_ (.A(_02798_),
    .B(_02797_),
    .Y(_02878_));
 sky130_fd_sc_hd__nor2_1 _22572_ (.A(_02798_),
    .B(_02797_),
    .Y(_02879_));
 sky130_fd_sc_hd__a21o_1 _22573_ (.A1(_02813_),
    .A2(_02878_),
    .B1(_02879_),
    .X(_02880_));
 sky130_fd_sc_hd__inv_1 _22574_ (.A(_02799_),
    .Y(_02881_));
 sky130_fd_sc_hd__nand3_1 _22575_ (.A(_02881_),
    .B(_02813_),
    .C(_02879_),
    .Y(_02882_));
 sky130_fd_sc_hd__o221ai_1 _22576_ (.A1(_02813_),
    .A2(_02878_),
    .B1(_02880_),
    .B2(_02881_),
    .C1(_02882_),
    .Y(_02883_));
 sky130_fd_sc_hd__nor2_1 _22577_ (.A(_02781_),
    .B(_02796_),
    .Y(_02884_));
 sky130_fd_sc_hd__inv_1 _22578_ (.A(_02884_),
    .Y(_02885_));
 sky130_fd_sc_hd__or2_4 _22579_ (.A(_02811_),
    .B(_02812_),
    .X(_02886_));
 sky130_fd_sc_hd__maj3_1 _22580_ (.A(_02807_),
    .B(_02808_),
    .C(_02809_),
    .X(_02887_));
 sky130_fd_sc_hd__a22o_1 _22581_ (.A1(_09340_),
    .A2(_02074_),
    .B1(_02078_),
    .B2(_09348_),
    .X(_02888_));
 sky130_fd_sc_hd__a221oi_4 _22582_ (.A1(_10484_),
    .A2(_02072_),
    .B1(_02076_),
    .B2(_10492_),
    .C1(_02888_),
    .Y(_02889_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_337 ();
 sky130_fd_sc_hd__nand2_1 _22584_ (.A(_02016_),
    .B(_02889_),
    .Y(_02891_));
 sky130_fd_sc_hd__mux2i_2 _22585_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[60] ),
    .A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[44] ),
    .S(net315),
    .Y(_02892_));
 sky130_fd_sc_hd__nand2_1 _22586_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[60] ),
    .B(net322),
    .Y(_02893_));
 sky130_fd_sc_hd__o21ai_4 _22587_ (.A1(_08280_),
    .A2(_02892_),
    .B1(_02893_),
    .Y(_02894_));
 sky130_fd_sc_hd__nand4_4 _22588_ (.A(_09534_),
    .B(_09542_),
    .C(_09552_),
    .D(_01968_),
    .Y(_02895_));
 sky130_fd_sc_hd__nand4_4 _22589_ (.A(_10628_),
    .B(_10636_),
    .C(_10643_),
    .D(_01720_),
    .Y(_02896_));
 sky130_fd_sc_hd__nand2_2 _22590_ (.A(_02895_),
    .B(_02896_),
    .Y(_02897_));
 sky130_fd_sc_hd__nand2_1 _22591_ (.A(_02032_),
    .B(_02897_),
    .Y(_02898_));
 sky130_fd_sc_hd__xnor3_2 _22592_ (.A(_02891_),
    .B(_02894_),
    .C(_02898_),
    .X(_02899_));
 sky130_fd_sc_hd__maj3_2 _22593_ (.A(_02801_),
    .B(_02804_),
    .C(_02805_),
    .X(_02900_));
 sky130_fd_sc_hd__maj3_1 _22594_ (.A(_02787_),
    .B(_02788_),
    .C(_02789_),
    .X(_02901_));
 sky130_fd_sc_hd__xnor2_1 _22595_ (.A(_02900_),
    .B(_02901_),
    .Y(_02902_));
 sky130_fd_sc_hd__xnor2_1 _22596_ (.A(_02899_),
    .B(_02902_),
    .Y(_02903_));
 sky130_fd_sc_hd__xor2_1 _22597_ (.A(_02903_),
    .B(_02887_),
    .X(_02904_));
 sky130_fd_sc_hd__xor2_1 _22598_ (.A(_02886_),
    .B(_02904_),
    .X(_02905_));
 sky130_fd_sc_hd__nand2_1 _22599_ (.A(_02782_),
    .B(_02792_),
    .Y(_02906_));
 sky130_fd_sc_hd__nand2_1 _22600_ (.A(_02795_),
    .B(_02906_),
    .Y(_02907_));
 sky130_fd_sc_hd__o21ai_1 _22601_ (.A1(_02782_),
    .A2(_02792_),
    .B1(_02907_),
    .Y(_02908_));
 sky130_fd_sc_hd__xnor2_2 _22602_ (.A(_02908_),
    .B(_02905_),
    .Y(_02909_));
 sky130_fd_sc_hd__nand2_1 _22603_ (.A(_02786_),
    .B(_02790_),
    .Y(_02910_));
 sky130_fd_sc_hd__nor2_1 _22604_ (.A(_02786_),
    .B(_02790_),
    .Y(_02911_));
 sky130_fd_sc_hd__a21oi_1 _22605_ (.A1(_02791_),
    .A2(_02910_),
    .B1(_02911_),
    .Y(_02912_));
 sky130_fd_sc_hd__nand2_2 _22606_ (.A(_02780_),
    .B(_02779_),
    .Y(_02913_));
 sky130_fd_sc_hd__a211oi_1 _22607_ (.A1(net306),
    .A2(net322),
    .B1(net735),
    .C1(_02692_),
    .Y(_02914_));
 sky130_fd_sc_hd__a221oi_4 _22608_ (.A1(net1186),
    .A2(_01712_),
    .B1(_02503_),
    .B2(net1035),
    .C1(_02061_),
    .Y(_02915_));
 sky130_fd_sc_hd__a221oi_2 _22609_ (.A1(net748),
    .A2(net322),
    .B1(_02586_),
    .B2(_02588_),
    .C1(net1051),
    .Y(_02916_));
 sky130_fd_sc_hd__xnor3_2 _22610_ (.A(_02914_),
    .B(_02916_),
    .C(_02915_),
    .X(_02917_));
 sky130_fd_sc_hd__and4_4 _22611_ (.A(_02391_),
    .B(_02392_),
    .C(_02393_),
    .D(_02395_),
    .X(_02918_));
 sky130_fd_sc_hd__o211ai_2 _22612_ (.A1(net913),
    .A2(net321),
    .B1(_02307_),
    .C1(_02918_),
    .Y(_02919_));
 sky130_fd_sc_hd__nand3_2 _22613_ (.A(_02436_),
    .B(_02424_),
    .C(_02425_),
    .Y(_02920_));
 sky130_fd_sc_hd__or3_4 _22614_ (.A(_02300_),
    .B(_02299_),
    .C(net1069),
    .X(_02921_));
 sky130_fd_sc_hd__xnor3_1 _22615_ (.A(_02919_),
    .B(_02920_),
    .C(_02921_),
    .X(_02922_));
 sky130_fd_sc_hd__maj3_2 _22616_ (.A(_02783_),
    .B(_02784_),
    .C(_02785_),
    .X(_02923_));
 sky130_fd_sc_hd__xnor2_1 _22617_ (.A(_02922_),
    .B(_02923_),
    .Y(_02924_));
 sky130_fd_sc_hd__xnor2_2 _22618_ (.A(net1510),
    .B(_02924_),
    .Y(_02925_));
 sky130_fd_sc_hd__xor2_2 _22619_ (.A(_02925_),
    .B(_02913_),
    .X(_02926_));
 sky130_fd_sc_hd__xnor2_2 _22620_ (.A(_02926_),
    .B(_02912_),
    .Y(_02927_));
 sky130_fd_sc_hd__nor2_1 _22621_ (.A(_02779_),
    .B(_02780_),
    .Y(_02928_));
 sky130_fd_sc_hd__nor3b_2 _22622_ (.A(_02775_),
    .B(_02928_),
    .C_N(_02913_),
    .Y(_02929_));
 sky130_fd_sc_hd__o31ai_4 _22623_ (.A1(_09505_),
    .A2(_09518_),
    .A3(_09523_),
    .B1(net320),
    .Y(_02930_));
 sky130_fd_sc_hd__nand4_4 _22624_ (.A(_10603_),
    .B(_10614_),
    .C(_10619_),
    .D(net321),
    .Y(_02931_));
 sky130_fd_sc_hd__and2_4 _22625_ (.A(_02931_),
    .B(net1223),
    .X(_02932_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_335 ();
 sky130_fd_sc_hd__nor2_1 _22628_ (.A(net1177),
    .B(_02932_),
    .Y(_02935_));
 sky130_fd_sc_hd__a21o_4 _22629_ (.A1(net307),
    .A2(_01712_),
    .B1(net1221),
    .X(_02936_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_333 ();
 sky130_fd_sc_hd__nor2_1 _22632_ (.A(net790),
    .B(_02936_),
    .Y(_02939_));
 sky130_fd_sc_hd__xnor2_1 _22633_ (.A(_02935_),
    .B(_02939_),
    .Y(_02940_));
 sky130_fd_sc_hd__o22ai_1 _22634_ (.A1(net939),
    .A2(_02513_),
    .B1(net1194),
    .B2(net781),
    .Y(_02941_));
 sky130_fd_sc_hd__nor4_1 _22635_ (.A(net1172),
    .B(net939),
    .C(_02513_),
    .D(net1194),
    .Y(_02942_));
 sky130_fd_sc_hd__a21oi_1 _22636_ (.A1(_02776_),
    .A2(_02941_),
    .B1(_02942_),
    .Y(_02943_));
 sky130_fd_sc_hd__nor2_1 _22637_ (.A(_02080_),
    .B(_02513_),
    .Y(_02944_));
 sky130_fd_sc_hd__a211o_2 _22638_ (.A1(_01966_),
    .A2(_01970_),
    .B1(_02723_),
    .C1(net1157),
    .X(_02945_));
 sky130_fd_sc_hd__a221o_2 _22639_ (.A1(_02619_),
    .A2(_01712_),
    .B1(_02083_),
    .B2(_02085_),
    .C1(_02621_),
    .X(_02946_));
 sky130_fd_sc_hd__xnor2_1 _22640_ (.A(_02945_),
    .B(_02946_),
    .Y(_02947_));
 sky130_fd_sc_hd__xnor2_1 _22641_ (.A(_02944_),
    .B(_02947_),
    .Y(_02948_));
 sky130_fd_sc_hd__xor2_1 _22642_ (.A(_02943_),
    .B(_02948_),
    .X(_02949_));
 sky130_fd_sc_hd__xnor2_1 _22643_ (.A(_02940_),
    .B(_02949_),
    .Y(_02950_));
 sky130_fd_sc_hd__xnor2_1 _22644_ (.A(_02929_),
    .B(_02950_),
    .Y(_02951_));
 sky130_fd_sc_hd__xnor2_1 _22645_ (.A(_02927_),
    .B(_02951_),
    .Y(_02952_));
 sky130_fd_sc_hd__xnor3_2 _22646_ (.A(_02885_),
    .B(_02909_),
    .C(_02952_),
    .X(_02953_));
 sky130_fd_sc_hd__xor2_1 _22647_ (.A(_02883_),
    .B(_02953_),
    .X(_02954_));
 sky130_fd_sc_hd__nor2_1 _22648_ (.A(_02618_),
    .B(_02617_),
    .Y(_02955_));
 sky130_fd_sc_hd__o21ai_0 _22649_ (.A1(_02709_),
    .A2(_02955_),
    .B1(_02710_),
    .Y(_02956_));
 sky130_fd_sc_hd__nor2_1 _22650_ (.A(_02741_),
    .B(_02743_),
    .Y(_02957_));
 sky130_fd_sc_hd__nand2_1 _22651_ (.A(_02618_),
    .B(_02617_),
    .Y(_02958_));
 sky130_fd_sc_hd__nand2_1 _22652_ (.A(_02626_),
    .B(_02958_),
    .Y(_02959_));
 sky130_fd_sc_hd__a21oi_1 _22653_ (.A1(_02741_),
    .A2(_02959_),
    .B1(_02955_),
    .Y(_02960_));
 sky130_fd_sc_hd__mux2i_1 _22654_ (.A0(_02957_),
    .A1(_02960_),
    .S(_02711_),
    .Y(_02961_));
 sky130_fd_sc_hd__maj3_1 _22655_ (.A(_02956_),
    .B(_02961_),
    .C(_02816_),
    .X(_02962_));
 sky130_fd_sc_hd__nor2_2 _22656_ (.A(_02954_),
    .B(_02962_),
    .Y(_02963_));
 sky130_fd_sc_hd__and2_2 _22657_ (.A(_02954_),
    .B(_02962_),
    .X(_02964_));
 sky130_fd_sc_hd__nor2_4 _22658_ (.A(_02963_),
    .B(_02964_),
    .Y(_02965_));
 sky130_fd_sc_hd__nand2_2 _22659_ (.A(_02823_),
    .B(_02825_),
    .Y(_02966_));
 sky130_fd_sc_hd__o21ai_4 _22660_ (.A1(_02750_),
    .A2(_02966_),
    .B1(_02822_),
    .Y(_02967_));
 sky130_fd_sc_hd__xnor2_4 _22661_ (.A(_02965_),
    .B(_02967_),
    .Y(_02968_));
 sky130_fd_sc_hd__mux2i_4 _22662_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[44] ),
    .A1(_02968_),
    .S(_02169_),
    .Y(_02969_));
 sky130_fd_sc_hd__nor2_1 _22663_ (.A(net442),
    .B(_02969_),
    .Y(_02970_));
 sky130_fd_sc_hd__a211oi_4 _22664_ (.A1(net442),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[44] ),
    .B1(net739),
    .C1(_02970_),
    .Y(_02971_));
 sky130_fd_sc_hd__a21oi_2 _22665_ (.A1(net739),
    .A2(_02877_),
    .B1(_02971_),
    .Y(_02972_));
 sky130_fd_sc_hd__nor3_2 _22666_ (.A(_11426_),
    .B(_02646_),
    .C(_02972_),
    .Y(_02973_));
 sky130_fd_sc_hd__a21oi_4 _22667_ (.A1(_02646_),
    .A2(_02861_),
    .B1(_02973_),
    .Y(_02974_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_332 ();
 sky130_fd_sc_hd__nand2_1 _22669_ (.A(_02119_),
    .B(_02974_),
    .Y(_02976_));
 sky130_fd_sc_hd__nand2_1 _22670_ (.A(\gen_regfile_ff.register_file_i.rf_reg[140] ),
    .B(_02123_),
    .Y(_02977_));
 sky130_fd_sc_hd__nand2_1 _22671_ (.A(_02976_),
    .B(_02977_),
    .Y(_00523_));
 sky130_fd_sc_hd__mux4_1 _22672_ (.A0(net31),
    .A1(net40),
    .A2(net48),
    .A3(net54),
    .S0(\load_store_unit_i.rdata_offset_q[0] ),
    .S1(\load_store_unit_i.rdata_offset_q[1] ),
    .X(_02978_));
 sky130_fd_sc_hd__mux4_1 _22673_ (.A0(net31),
    .A1(\load_store_unit_i.rdata_q[21] ),
    .A2(\load_store_unit_i.rdata_q[29] ),
    .A3(net54),
    .S0(\load_store_unit_i.rdata_offset_q[0] ),
    .S1(\load_store_unit_i.rdata_offset_q[1] ),
    .X(_02979_));
 sky130_fd_sc_hd__a221oi_4 _22674_ (.A1(\load_store_unit_i.data_type_q[2] ),
    .A2(_02978_),
    .B1(_02979_),
    .B2(_01674_),
    .C1(_02549_),
    .Y(_02980_));
 sky130_fd_sc_hd__nor2_1 _22675_ (.A(_01738_),
    .B(_02184_),
    .Y(_02981_));
 sky130_fd_sc_hd__a21oi_1 _22676_ (.A1(_01738_),
    .A2(_02211_),
    .B1(_02981_),
    .Y(_02982_));
 sky130_fd_sc_hd__a31oi_1 _22677_ (.A1(_01758_),
    .A2(_01738_),
    .A3(_02186_),
    .B1(_02865_),
    .Y(_02983_));
 sky130_fd_sc_hd__nand2_1 _22678_ (.A(_02558_),
    .B(_02983_),
    .Y(_02984_));
 sky130_fd_sc_hd__o21ai_1 _22679_ (.A1(_02558_),
    .A2(_02982_),
    .B1(_02984_),
    .Y(_02985_));
 sky130_fd_sc_hd__mux2i_1 _22680_ (.A0(_02220_),
    .A1(_02660_),
    .S(_01738_),
    .Y(_02986_));
 sky130_fd_sc_hd__o21ai_1 _22681_ (.A1(_02558_),
    .A2(_02986_),
    .B1(_02658_),
    .Y(_02987_));
 sky130_fd_sc_hd__nand2_1 _22682_ (.A(net295),
    .B(_02987_),
    .Y(_02988_));
 sky130_fd_sc_hd__o21ai_1 _22683_ (.A1(net295),
    .A2(_02985_),
    .B1(_02988_),
    .Y(_02989_));
 sky130_fd_sc_hd__nand3_1 _22684_ (.A(net1465),
    .B(_09484_),
    .C(_02228_),
    .Y(_02990_));
 sky130_fd_sc_hd__o21ai_0 _22685_ (.A1(_09484_),
    .A2(_01902_),
    .B1(_02990_),
    .Y(_02991_));
 sky130_fd_sc_hd__a21oi_1 _22686_ (.A1(_09484_),
    .A2(_02233_),
    .B1(net1465),
    .Y(_02992_));
 sky130_fd_sc_hd__a21oi_1 _22687_ (.A1(_02225_),
    .A2(_02991_),
    .B1(_02992_),
    .Y(_02993_));
 sky130_fd_sc_hd__a221oi_2 _22688_ (.A1(net1569),
    .A2(_01929_),
    .B1(_02989_),
    .B2(_01734_),
    .C1(_02993_),
    .Y(_02994_));
 sky130_fd_sc_hd__nand2_1 _22689_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[45] ),
    .B(_01698_),
    .Y(_02995_));
 sky130_fd_sc_hd__inv_1 _22690_ (.A(_02963_),
    .Y(_02996_));
 sky130_fd_sc_hd__a21oi_2 _22691_ (.A1(_02996_),
    .A2(_02967_),
    .B1(_02964_),
    .Y(_02997_));
 sky130_fd_sc_hd__nor2_1 _22692_ (.A(_02940_),
    .B(_02949_),
    .Y(_02998_));
 sky130_fd_sc_hd__nor2b_2 _22693_ (.A(_02943_),
    .B_N(_02948_),
    .Y(_02999_));
 sky130_fd_sc_hd__inv_1 _22694_ (.A(_02917_),
    .Y(_03000_));
 sky130_fd_sc_hd__maj3_1 _22695_ (.A(_02922_),
    .B(_03000_),
    .C(_02923_),
    .X(_03001_));
 sky130_fd_sc_hd__or3_4 _22696_ (.A(net1069),
    .B(_02417_),
    .C(_02419_),
    .X(_03002_));
 sky130_fd_sc_hd__nand2_1 _22697_ (.A(_02301_),
    .B(_02918_),
    .Y(_03003_));
 sky130_fd_sc_hd__nand2_2 _22698_ (.A(net1035),
    .B(_02503_),
    .Y(_03004_));
 sky130_fd_sc_hd__nand2_1 _22699_ (.A(net1180),
    .B(_03004_),
    .Y(_03005_));
 sky130_fd_sc_hd__xnor3_1 _22700_ (.A(_03002_),
    .B(_03003_),
    .C(_03005_),
    .X(_03006_));
 sky130_fd_sc_hd__a211oi_2 _22701_ (.A1(net306),
    .A2(net322),
    .B1(net736),
    .C1(_02800_),
    .Y(_03007_));
 sky130_fd_sc_hd__a221oi_4 _22702_ (.A1(net309),
    .A2(_01712_),
    .B1(_02586_),
    .B2(_02588_),
    .C1(_02061_),
    .Y(_03008_));
 sky130_fd_sc_hd__a211oi_2 _22703_ (.A1(net750),
    .A2(net322),
    .B1(net1051),
    .C1(_02692_),
    .Y(_03009_));
 sky130_fd_sc_hd__xnor3_2 _22704_ (.A(_03007_),
    .B(_03008_),
    .C(_03009_),
    .X(_03010_));
 sky130_fd_sc_hd__maj3_2 _22705_ (.A(_02919_),
    .B(_02921_),
    .C(_02920_),
    .X(_03011_));
 sky130_fd_sc_hd__xnor2_2 _22706_ (.A(_03010_),
    .B(_03011_),
    .Y(_03012_));
 sky130_fd_sc_hd__xnor2_1 _22707_ (.A(_03012_),
    .B(_03006_),
    .Y(_03013_));
 sky130_fd_sc_hd__xor3_1 _22708_ (.A(_02999_),
    .B(_03001_),
    .C(_03013_),
    .X(_03014_));
 sky130_fd_sc_hd__nand2_1 _22709_ (.A(net1223),
    .B(_02931_),
    .Y(_03015_));
 sky130_fd_sc_hd__nand2_1 _22710_ (.A(_02014_),
    .B(_03015_),
    .Y(_03016_));
 sky130_fd_sc_hd__mux2_4 _22711_ (.A0(_09482_),
    .A1(_10590_),
    .S(net322),
    .X(_03017_));
 sky130_fd_sc_hd__nand2_1 _22712_ (.A(_01998_),
    .B(_03017_),
    .Y(_03018_));
 sky130_fd_sc_hd__nand2_1 _22713_ (.A(_02158_),
    .B(_02774_),
    .Y(_03019_));
 sky130_fd_sc_hd__xor2_1 _22714_ (.A(_03018_),
    .B(_03019_),
    .X(_03020_));
 sky130_fd_sc_hd__xnor2_2 _22715_ (.A(_03016_),
    .B(_03020_),
    .Y(_03021_));
 sky130_fd_sc_hd__nand2_1 _22716_ (.A(_02160_),
    .B(_02727_),
    .Y(_03022_));
 sky130_fd_sc_hd__nand2b_1 _22717_ (.A_N(_02513_),
    .B(_02436_),
    .Y(_03023_));
 sky130_fd_sc_hd__or2_0 _22718_ (.A(_02080_),
    .B(_02622_),
    .X(_03024_));
 sky130_fd_sc_hd__xor3_1 _22719_ (.A(_03022_),
    .B(_03023_),
    .C(_03024_),
    .X(_03025_));
 sky130_fd_sc_hd__nor3_1 _22720_ (.A(_02089_),
    .B(_02936_),
    .C(_02932_),
    .Y(_03026_));
 sky130_fd_sc_hd__o31a_1 _22721_ (.A1(_02080_),
    .A2(_02513_),
    .A3(_02945_),
    .B1(_02946_),
    .X(_03027_));
 sky130_fd_sc_hd__o21a_1 _22722_ (.A1(_02080_),
    .A2(_02513_),
    .B1(_02945_),
    .X(_03028_));
 sky130_fd_sc_hd__o2111ai_1 _22723_ (.A1(_02945_),
    .A2(_02946_),
    .B1(_02774_),
    .C1(_02304_),
    .D1(_03015_),
    .Y(_03029_));
 sky130_fd_sc_hd__a211oi_1 _22724_ (.A1(_02945_),
    .A2(_02946_),
    .B1(_02080_),
    .C1(_02513_),
    .Y(_03030_));
 sky130_fd_sc_hd__o32ai_2 _22725_ (.A1(_03026_),
    .A2(_03027_),
    .A3(_03028_),
    .B1(_03029_),
    .B2(_03030_),
    .Y(_03031_));
 sky130_fd_sc_hd__xnor2_1 _22726_ (.A(_03025_),
    .B(_03031_),
    .Y(_03032_));
 sky130_fd_sc_hd__xor2_1 _22727_ (.A(_03021_),
    .B(_03032_),
    .X(_03033_));
 sky130_fd_sc_hd__xor3_1 _22728_ (.A(_02998_),
    .B(_03014_),
    .C(_03033_),
    .X(_03034_));
 sky130_fd_sc_hd__inv_1 _22729_ (.A(_02929_),
    .Y(_03035_));
 sky130_fd_sc_hd__inv_1 _22730_ (.A(_02927_),
    .Y(_03036_));
 sky130_fd_sc_hd__maj3_2 _22731_ (.A(_03036_),
    .B(_03035_),
    .C(_02950_),
    .X(_03037_));
 sky130_fd_sc_hd__maj3_1 _22732_ (.A(_02913_),
    .B(_02912_),
    .C(_02925_),
    .X(_03038_));
 sky130_fd_sc_hd__or4_4 _22733_ (.A(_09432_),
    .B(_09437_),
    .C(_09444_),
    .D(_01720_),
    .X(_03039_));
 sky130_fd_sc_hd__nand4_4 _22734_ (.A(_10541_),
    .B(_10549_),
    .C(_10556_),
    .D(_01720_),
    .Y(_03040_));
 sky130_fd_sc_hd__nand2_4 _22735_ (.A(_03039_),
    .B(_03040_),
    .Y(_03041_));
 sky130_fd_sc_hd__nand2_1 _22736_ (.A(_02032_),
    .B(_03041_),
    .Y(_03042_));
 sky130_fd_sc_hd__mux2_1 _22737_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[61] ),
    .A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[45] ),
    .S(_13441_),
    .X(_03043_));
 sky130_fd_sc_hd__a22oi_4 _22738_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[61] ),
    .A2(_01702_),
    .B1(_03043_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .Y(_03044_));
 sky130_fd_sc_hd__a221oi_4 _22739_ (.A1(net659),
    .A2(_01712_),
    .B1(_02895_),
    .B2(_02896_),
    .C1(net780),
    .Y(_03045_));
 sky130_fd_sc_hd__xnor2_1 _22740_ (.A(_03044_),
    .B(_03045_),
    .Y(_03046_));
 sky130_fd_sc_hd__xnor2_2 _22741_ (.A(_03042_),
    .B(_03046_),
    .Y(_03047_));
 sky130_fd_sc_hd__maj3_1 _22742_ (.A(_02914_),
    .B(_02915_),
    .C(_02916_),
    .X(_03048_));
 sky130_fd_sc_hd__nand3_1 _22743_ (.A(_02016_),
    .B(_02889_),
    .C(_02894_),
    .Y(_03049_));
 sky130_fd_sc_hd__a21oi_1 _22744_ (.A1(_02016_),
    .A2(_02889_),
    .B1(_02894_),
    .Y(_03050_));
 sky130_fd_sc_hd__a21oi_1 _22745_ (.A1(_02898_),
    .A2(_03049_),
    .B1(_03050_),
    .Y(_03051_));
 sky130_fd_sc_hd__xnor2_1 _22746_ (.A(_03048_),
    .B(_03051_),
    .Y(_03052_));
 sky130_fd_sc_hd__xnor2_2 _22747_ (.A(_03047_),
    .B(_03052_),
    .Y(_03053_));
 sky130_fd_sc_hd__nor2_1 _22748_ (.A(_02900_),
    .B(_02901_),
    .Y(_03054_));
 sky130_fd_sc_hd__nand2_1 _22749_ (.A(_02900_),
    .B(_02901_),
    .Y(_03055_));
 sky130_fd_sc_hd__o21ai_2 _22750_ (.A1(_02899_),
    .A2(_03054_),
    .B1(_03055_),
    .Y(_03056_));
 sky130_fd_sc_hd__xnor2_1 _22751_ (.A(_03053_),
    .B(_03056_),
    .Y(_03057_));
 sky130_fd_sc_hd__nand2b_1 _22752_ (.A_N(_02903_),
    .B(_02887_),
    .Y(_03058_));
 sky130_fd_sc_hd__xnor2_1 _22753_ (.A(_03057_),
    .B(_03058_),
    .Y(_03059_));
 sky130_fd_sc_hd__xnor2_1 _22754_ (.A(_03038_),
    .B(_03059_),
    .Y(_03060_));
 sky130_fd_sc_hd__xnor3_4 _22755_ (.A(_03060_),
    .B(_03037_),
    .C(_03034_),
    .X(_03061_));
 sky130_fd_sc_hd__maj3_2 _22756_ (.A(_02885_),
    .B(_02909_),
    .C(_02952_),
    .X(_03062_));
 sky130_fd_sc_hd__nand2_1 _22757_ (.A(_02886_),
    .B(_02904_),
    .Y(_03063_));
 sky130_fd_sc_hd__nor2_1 _22758_ (.A(_02886_),
    .B(_02904_),
    .Y(_03064_));
 sky130_fd_sc_hd__a21oi_2 _22759_ (.A1(_03063_),
    .A2(_02908_),
    .B1(_03064_),
    .Y(_03065_));
 sky130_fd_sc_hd__xor2_2 _22760_ (.A(_03062_),
    .B(_03065_),
    .X(_03066_));
 sky130_fd_sc_hd__xnor2_4 _22761_ (.A(_03061_),
    .B(_03066_),
    .Y(_03067_));
 sky130_fd_sc_hd__o21ai_2 _22762_ (.A1(_02879_),
    .A2(_02953_),
    .B1(_02813_),
    .Y(_03068_));
 sky130_fd_sc_hd__a21oi_1 _22763_ (.A1(_02798_),
    .A2(_02797_),
    .B1(_02799_),
    .Y(_03069_));
 sky130_fd_sc_hd__o21ai_1 _22764_ (.A1(_02880_),
    .A2(_03069_),
    .B1(_02953_),
    .Y(_03070_));
 sky130_fd_sc_hd__o21ai_4 _22765_ (.A1(_02799_),
    .A2(_03068_),
    .B1(_03070_),
    .Y(_03071_));
 sky130_fd_sc_hd__xor2_4 _22766_ (.A(_03071_),
    .B(_03067_),
    .X(_03072_));
 sky130_fd_sc_hd__xor2_4 _22767_ (.A(_02997_),
    .B(_03072_),
    .X(_03073_));
 sky130_fd_sc_hd__nand2_1 _22768_ (.A(_02169_),
    .B(_03073_),
    .Y(_03074_));
 sky130_fd_sc_hd__nand2_2 _22769_ (.A(_02995_),
    .B(_03074_),
    .Y(_03075_));
 sky130_fd_sc_hd__nand2b_1 _22770_ (.A_N(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[45] ),
    .B(net442),
    .Y(_03076_));
 sky130_fd_sc_hd__o211ai_4 _22771_ (.A1(net442),
    .A2(_03075_),
    .B1(_03076_),
    .C1(net313),
    .Y(_03077_));
 sky130_fd_sc_hd__o21ai_4 _22772_ (.A1(net313),
    .A2(_02994_),
    .B1(_03077_),
    .Y(_03078_));
 sky130_fd_sc_hd__o21ai_2 _22773_ (.A1(_11446_),
    .A2(_03078_),
    .B1(net1483),
    .Y(_03079_));
 sky130_fd_sc_hd__o21ai_4 _22774_ (.A1(net266),
    .A2(_02980_),
    .B1(_03079_),
    .Y(_03080_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_331 ();
 sky130_fd_sc_hd__nand2_1 _22776_ (.A(_02119_),
    .B(_03080_),
    .Y(_03082_));
 sky130_fd_sc_hd__nand2_1 _22777_ (.A(\gen_regfile_ff.register_file_i.rf_reg[141] ),
    .B(_02123_),
    .Y(_03083_));
 sky130_fd_sc_hd__nand2_1 _22778_ (.A(_03082_),
    .B(_03083_),
    .Y(_00524_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_330 ();
 sky130_fd_sc_hd__nand2_1 _22780_ (.A(_01916_),
    .B(_02761_),
    .Y(_03085_));
 sky130_fd_sc_hd__nand2_1 _22781_ (.A(\gen_regfile_ff.register_file_i.rf_reg[42] ),
    .B(_01921_),
    .Y(_03086_));
 sky130_fd_sc_hd__nand2_1 _22782_ (.A(_03085_),
    .B(_03086_),
    .Y(_00525_));
 sky130_fd_sc_hd__mux4_1 _22783_ (.A0(net32),
    .A1(net41),
    .A2(net50),
    .A3(net55),
    .S0(\load_store_unit_i.rdata_offset_q[0] ),
    .S1(\load_store_unit_i.rdata_offset_q[1] ),
    .X(_03087_));
 sky130_fd_sc_hd__mux4_1 _22784_ (.A0(net32),
    .A1(\load_store_unit_i.rdata_q[22] ),
    .A2(\load_store_unit_i.rdata_q[30] ),
    .A3(net55),
    .S0(\load_store_unit_i.rdata_offset_q[0] ),
    .S1(\load_store_unit_i.rdata_offset_q[1] ),
    .X(_03088_));
 sky130_fd_sc_hd__a221oi_2 _22785_ (.A1(\load_store_unit_i.data_type_q[2] ),
    .A2(_03087_),
    .B1(_03088_),
    .B2(_01674_),
    .C1(_02549_),
    .Y(_03089_));
 sky130_fd_sc_hd__nand2_1 _22786_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[46] ),
    .B(_01698_),
    .Y(_03090_));
 sky130_fd_sc_hd__maj3_2 _22787_ (.A(_03062_),
    .B(_03061_),
    .C(_03065_),
    .X(_03091_));
 sky130_fd_sc_hd__inv_1 _22788_ (.A(_03034_),
    .Y(_03092_));
 sky130_fd_sc_hd__maj3_1 _22789_ (.A(_03092_),
    .B(_03037_),
    .C(_03060_),
    .X(_03093_));
 sky130_fd_sc_hd__and2_1 _22790_ (.A(_03053_),
    .B(_03056_),
    .X(_03094_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_329 ();
 sky130_fd_sc_hd__maj3_2 _22792_ (.A(_02999_),
    .B(_03001_),
    .C(net1183),
    .X(_03096_));
 sky130_fd_sc_hd__and2_4 _22793_ (.A(_02895_),
    .B(_02896_),
    .X(_03097_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_328 ();
 sky130_fd_sc_hd__maj3_1 _22795_ (.A(net949),
    .B(_03097_),
    .C(_03044_),
    .X(_03099_));
 sky130_fd_sc_hd__and2_4 _22796_ (.A(_03039_),
    .B(_03040_),
    .X(_03100_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_327 ();
 sky130_fd_sc_hd__nor2_2 _22798_ (.A(_01982_),
    .B(_03100_),
    .Y(_03102_));
 sky130_fd_sc_hd__nor4_1 _22799_ (.A(net857),
    .B(_03097_),
    .C(_03041_),
    .D(_03044_),
    .Y(_03103_));
 sky130_fd_sc_hd__nor4_1 _22800_ (.A(net949),
    .B(_02016_),
    .C(_03100_),
    .D(_03044_),
    .Y(_03104_));
 sky130_fd_sc_hd__a211o_1 _22801_ (.A1(_03099_),
    .A2(_03102_),
    .B1(_03103_),
    .C1(_03104_),
    .X(_03105_));
 sky130_fd_sc_hd__mux2_1 _22802_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[62] ),
    .A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[46] ),
    .S(_13441_),
    .X(_03106_));
 sky130_fd_sc_hd__a22oi_4 _22803_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[62] ),
    .A2(_01702_),
    .B1(_03106_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .Y(_03107_));
 sky130_fd_sc_hd__nor4b_1 _22804_ (.A(net389),
    .B(_10768_),
    .C(_01968_),
    .D_N(_10771_),
    .Y(_03108_));
 sky130_fd_sc_hd__nor2_1 _22805_ (.A(net1282),
    .B(_01720_),
    .Y(_03109_));
 sky130_fd_sc_hd__a31oi_1 _22806_ (.A1(_09617_),
    .A2(_09620_),
    .A3(_03109_),
    .B1(_08512_),
    .Y(_03110_));
 sky130_fd_sc_hd__nand3_1 _22807_ (.A(net1140),
    .B(_09613_),
    .C(_01968_),
    .Y(_03111_));
 sky130_fd_sc_hd__nand3_1 _22808_ (.A(net1140),
    .B(_10775_),
    .C(_01720_),
    .Y(_03112_));
 sky130_fd_sc_hd__and4b_4 _22809_ (.A_N(_03108_),
    .B(_03110_),
    .C(_03111_),
    .D(_03112_),
    .X(_03113_));
 sky130_fd_sc_hd__o211ai_2 _22810_ (.A1(_10780_),
    .A2(_10782_),
    .B1(_01720_),
    .C1(_08309_),
    .Y(_03114_));
 sky130_fd_sc_hd__nand3_1 _22811_ (.A(net1140),
    .B(_10786_),
    .C(_01720_),
    .Y(_03115_));
 sky130_fd_sc_hd__or3_1 _22812_ (.A(_08309_),
    .B(_09624_),
    .C(_01720_),
    .X(_03116_));
 sky130_fd_sc_hd__o21ai_1 _22813_ (.A1(_09627_),
    .A2(_09629_),
    .B1(_03109_),
    .Y(_03117_));
 sky130_fd_sc_hd__a41oi_4 _22814_ (.A1(_03115_),
    .A2(_03114_),
    .A3(_03116_),
    .A4(_03117_),
    .B1(net383),
    .Y(_03118_));
 sky130_fd_sc_hd__or2_4 _22815_ (.A(_03113_),
    .B(net1063),
    .X(_03119_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_326 ();
 sky130_fd_sc_hd__or3_1 _22817_ (.A(net950),
    .B(_03107_),
    .C(_03119_),
    .X(_03121_));
 sky130_fd_sc_hd__o21ai_2 _22818_ (.A1(net949),
    .A2(_03119_),
    .B1(_03107_),
    .Y(_03122_));
 sky130_fd_sc_hd__maj3_1 _22819_ (.A(_03007_),
    .B(_03008_),
    .C(_03009_),
    .X(_03123_));
 sky130_fd_sc_hd__nand3_1 _22820_ (.A(_03121_),
    .B(_03122_),
    .C(_03123_),
    .Y(_03124_));
 sky130_fd_sc_hd__or2_0 _22821_ (.A(_03008_),
    .B(_03009_),
    .X(_03125_));
 sky130_fd_sc_hd__and2_0 _22822_ (.A(_03008_),
    .B(_03009_),
    .X(_03126_));
 sky130_fd_sc_hd__a221o_1 _22823_ (.A1(_03121_),
    .A2(_03122_),
    .B1(_03125_),
    .B2(_03007_),
    .C1(_03126_),
    .X(_03127_));
 sky130_fd_sc_hd__nand3_1 _22824_ (.A(_03105_),
    .B(_03124_),
    .C(_03127_),
    .Y(_03128_));
 sky130_fd_sc_hd__a21o_1 _22825_ (.A1(_03124_),
    .A2(_03127_),
    .B1(_03105_),
    .X(_03129_));
 sky130_fd_sc_hd__maj3_1 _22826_ (.A(_03047_),
    .B(_03048_),
    .C(_03051_),
    .X(_03130_));
 sky130_fd_sc_hd__a21oi_2 _22827_ (.A1(_03128_),
    .A2(_03129_),
    .B1(_03130_),
    .Y(_03131_));
 sky130_fd_sc_hd__and3_4 _22828_ (.A(_03128_),
    .B(_03129_),
    .C(_03130_),
    .X(_03132_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_325 ();
 sky130_fd_sc_hd__nor2_1 _22830_ (.A(_03131_),
    .B(_03132_),
    .Y(_03134_));
 sky130_fd_sc_hd__xnor3_1 _22831_ (.A(_03094_),
    .B(_03096_),
    .C(_03134_),
    .X(_03135_));
 sky130_fd_sc_hd__maj3_2 _22832_ (.A(_03003_),
    .B(_03002_),
    .C(_03005_),
    .X(_03136_));
 sky130_fd_sc_hd__a211oi_1 _22833_ (.A1(net748),
    .A2(net322),
    .B1(net1051),
    .C1(net1335),
    .Y(_03137_));
 sky130_fd_sc_hd__a211oi_2 _22834_ (.A1(net309),
    .A2(_01712_),
    .B1(_02061_),
    .C1(_02692_),
    .Y(_03138_));
 sky130_fd_sc_hd__a221oi_2 _22835_ (.A1(net306),
    .A2(net322),
    .B1(_02895_),
    .B2(_02896_),
    .C1(net735),
    .Y(_03139_));
 sky130_fd_sc_hd__xnor2_1 _22836_ (.A(_03138_),
    .B(_03139_),
    .Y(_03140_));
 sky130_fd_sc_hd__xor2_1 _22837_ (.A(_03137_),
    .B(_03140_),
    .X(_03141_));
 sky130_fd_sc_hd__and2_4 _22838_ (.A(_02586_),
    .B(_02588_),
    .X(_03142_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_324 ();
 sky130_fd_sc_hd__nor2_1 _22840_ (.A(net1286),
    .B(_03142_),
    .Y(_03144_));
 sky130_fd_sc_hd__nor2_1 _22841_ (.A(net1031),
    .B(_02426_),
    .Y(_03145_));
 sky130_fd_sc_hd__nor2_4 _22842_ (.A(_02289_),
    .B(net1277),
    .Y(_03146_));
 sky130_fd_sc_hd__xnor3_1 _22843_ (.A(_03144_),
    .B(_03145_),
    .C(_03146_),
    .X(_03147_));
 sky130_fd_sc_hd__xor3_1 _22844_ (.A(_03136_),
    .B(_03141_),
    .C(_03147_),
    .X(_03148_));
 sky130_fd_sc_hd__inv_1 _22845_ (.A(_03026_),
    .Y(_03149_));
 sky130_fd_sc_hd__o21ai_0 _22846_ (.A1(_02080_),
    .A2(_02513_),
    .B1(_02946_),
    .Y(_03150_));
 sky130_fd_sc_hd__o31ai_1 _22847_ (.A1(_02080_),
    .A2(_02513_),
    .A3(_02946_),
    .B1(_02945_),
    .Y(_03151_));
 sky130_fd_sc_hd__nand2_1 _22848_ (.A(_03150_),
    .B(_03151_),
    .Y(_03152_));
 sky130_fd_sc_hd__maj3_1 _22849_ (.A(_03025_),
    .B(_03149_),
    .C(_03152_),
    .X(_03153_));
 sky130_fd_sc_hd__nor2_1 _22850_ (.A(_03010_),
    .B(_03011_),
    .Y(_03154_));
 sky130_fd_sc_hd__nand2_1 _22851_ (.A(_03010_),
    .B(_03011_),
    .Y(_03155_));
 sky130_fd_sc_hd__o21ai_2 _22852_ (.A1(_03006_),
    .A2(_03154_),
    .B1(_03155_),
    .Y(_03156_));
 sky130_fd_sc_hd__xnor3_2 _22853_ (.A(_03156_),
    .B(_03153_),
    .C(net1160),
    .X(_03157_));
 sky130_fd_sc_hd__and2_0 _22854_ (.A(_03021_),
    .B(_03032_),
    .X(_03158_));
 sky130_fd_sc_hd__nor4_2 _22855_ (.A(_09592_),
    .B(_09594_),
    .C(_09597_),
    .D(net321),
    .Y(_03159_));
 sky130_fd_sc_hd__and4_4 _22856_ (.A(_09584_),
    .B(_09589_),
    .C(_09605_),
    .D(_03159_),
    .X(_03160_));
 sky130_fd_sc_hd__a21oi_4 _22857_ (.A1(net1163),
    .A2(net322),
    .B1(_03160_),
    .Y(_03161_));
 sky130_fd_sc_hd__nand2_2 _22858_ (.A(_01998_),
    .B(_03161_),
    .Y(_03162_));
 sky130_fd_sc_hd__nor2_1 _22859_ (.A(_01972_),
    .B(_02932_),
    .Y(_03163_));
 sky130_fd_sc_hd__nor2_1 _22860_ (.A(net1060),
    .B(_02936_),
    .Y(_03164_));
 sky130_fd_sc_hd__mux2i_4 _22861_ (.A0(_09482_),
    .A1(_10590_),
    .S(net322),
    .Y(_03165_));
 sky130_fd_sc_hd__nor2_4 _22862_ (.A(_03165_),
    .B(net790),
    .Y(_03166_));
 sky130_fd_sc_hd__xnor3_2 _22863_ (.A(_03163_),
    .B(_03164_),
    .C(_03166_),
    .X(_03167_));
 sky130_fd_sc_hd__xnor2_4 _22864_ (.A(_03162_),
    .B(_03167_),
    .Y(_03168_));
 sky130_fd_sc_hd__maj3_2 _22865_ (.A(_03016_),
    .B(_03018_),
    .C(_03019_),
    .X(_03169_));
 sky130_fd_sc_hd__nor2_1 _22866_ (.A(_02080_),
    .B(_02730_),
    .Y(_03170_));
 sky130_fd_sc_hd__nor2_1 _22867_ (.A(net1069),
    .B(_02513_),
    .Y(_03171_));
 sky130_fd_sc_hd__nor2_1 _22868_ (.A(_02150_),
    .B(net1193),
    .Y(_03172_));
 sky130_fd_sc_hd__xnor3_1 _22869_ (.A(_03172_),
    .B(_03171_),
    .C(_03170_),
    .X(_03173_));
 sky130_fd_sc_hd__maj3_1 _22870_ (.A(_03022_),
    .B(_03023_),
    .C(_03024_),
    .X(_03174_));
 sky130_fd_sc_hd__xor3_2 _22871_ (.A(_03174_),
    .B(_03173_),
    .C(_03169_),
    .X(_03175_));
 sky130_fd_sc_hd__xor2_4 _22872_ (.A(_03168_),
    .B(_03175_),
    .X(_03176_));
 sky130_fd_sc_hd__xnor3_4 _22873_ (.A(_03176_),
    .B(_03158_),
    .C(_03157_),
    .X(_03177_));
 sky130_fd_sc_hd__maj3_2 _22874_ (.A(_03014_),
    .B(_02998_),
    .C(_03033_),
    .X(_03178_));
 sky130_fd_sc_hd__xor2_1 _22875_ (.A(_03178_),
    .B(_03177_),
    .X(_03179_));
 sky130_fd_sc_hd__xnor2_1 _22876_ (.A(_03135_),
    .B(_03179_),
    .Y(_03180_));
 sky130_fd_sc_hd__maj3_1 _22877_ (.A(_03038_),
    .B(_03057_),
    .C(_03058_),
    .X(_03181_));
 sky130_fd_sc_hd__xnor2_1 _22878_ (.A(_03181_),
    .B(_03180_),
    .Y(_03182_));
 sky130_fd_sc_hd__xnor2_1 _22879_ (.A(_03093_),
    .B(_03182_),
    .Y(_03183_));
 sky130_fd_sc_hd__or2_0 _22880_ (.A(_03091_),
    .B(_03183_),
    .X(_03184_));
 sky130_fd_sc_hd__nand2_2 _22881_ (.A(_03091_),
    .B(_03183_),
    .Y(_03185_));
 sky130_fd_sc_hd__nand2_2 _22882_ (.A(_03184_),
    .B(_03185_),
    .Y(_03186_));
 sky130_fd_sc_hd__o2111ai_4 _22883_ (.A1(_02966_),
    .A2(_02750_),
    .B1(_03072_),
    .C1(_02822_),
    .D1(_02965_),
    .Y(_03187_));
 sky130_fd_sc_hd__nor2_4 _22884_ (.A(_03067_),
    .B(_03071_),
    .Y(_03188_));
 sky130_fd_sc_hd__nand2_1 _22885_ (.A(_03067_),
    .B(_03071_),
    .Y(_03189_));
 sky130_fd_sc_hd__o21a_2 _22886_ (.A1(_02996_),
    .A2(_03188_),
    .B1(_03189_),
    .X(_03190_));
 sky130_fd_sc_hd__nand2_1 _22887_ (.A(_03187_),
    .B(_03190_),
    .Y(_03191_));
 sky130_fd_sc_hd__xnor2_4 _22888_ (.A(_03186_),
    .B(_03191_),
    .Y(_03192_));
 sky130_fd_sc_hd__nand2_1 _22889_ (.A(_02169_),
    .B(_03192_),
    .Y(_03193_));
 sky130_fd_sc_hd__a21oi_2 _22890_ (.A1(_03090_),
    .A2(_03193_),
    .B1(_13335_),
    .Y(_03194_));
 sky130_fd_sc_hd__a21oi_2 _22891_ (.A1(net442),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[46] ),
    .B1(_03194_),
    .Y(_03195_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_323 ();
 sky130_fd_sc_hd__or2_0 _22893_ (.A(_09640_),
    .B(_01902_),
    .X(_03197_));
 sky130_fd_sc_hd__nand3_1 _22894_ (.A(_09608_),
    .B(_09640_),
    .C(_02228_),
    .Y(_03198_));
 sky130_fd_sc_hd__a21oi_1 _22895_ (.A1(_03197_),
    .A2(_03198_),
    .B1(_01893_),
    .Y(_03199_));
 sky130_fd_sc_hd__a21oi_1 _22896_ (.A1(_09640_),
    .A2(_02233_),
    .B1(_09608_),
    .Y(_03200_));
 sky130_fd_sc_hd__a31oi_1 _22897_ (.A1(_01758_),
    .A2(_01738_),
    .A3(_02218_),
    .B1(_02865_),
    .Y(_03201_));
 sky130_fd_sc_hd__nand2_1 _22898_ (.A(_01826_),
    .B(_02259_),
    .Y(_03202_));
 sky130_fd_sc_hd__o211ai_1 _22899_ (.A1(_01826_),
    .A2(_02264_),
    .B1(_03202_),
    .C1(_01743_),
    .Y(_03203_));
 sky130_fd_sc_hd__o21ai_0 _22900_ (.A1(_01743_),
    .A2(_03201_),
    .B1(_03203_),
    .Y(_03204_));
 sky130_fd_sc_hd__nor2_1 _22901_ (.A(_01826_),
    .B(_02562_),
    .Y(_03205_));
 sky130_fd_sc_hd__a21oi_1 _22902_ (.A1(_01826_),
    .A2(_02274_),
    .B1(_03205_),
    .Y(_03206_));
 sky130_fd_sc_hd__a21oi_1 _22903_ (.A1(_01743_),
    .A2(_03206_),
    .B1(_01943_),
    .Y(_03207_));
 sky130_fd_sc_hd__nor2_1 _22904_ (.A(_01773_),
    .B(_03207_),
    .Y(_03208_));
 sky130_fd_sc_hd__a21oi_1 _22905_ (.A1(_01773_),
    .A2(_03204_),
    .B1(_03208_),
    .Y(_03209_));
 sky130_fd_sc_hd__o22ai_1 _22906_ (.A1(_03199_),
    .A2(_03200_),
    .B1(_03209_),
    .B2(_01761_),
    .Y(_03210_));
 sky130_fd_sc_hd__a211oi_1 _22907_ (.A1(net155),
    .A2(_01929_),
    .B1(_03210_),
    .C1(net313),
    .Y(_03211_));
 sky130_fd_sc_hd__a21oi_2 _22908_ (.A1(_08272_),
    .A2(_03195_),
    .B1(_03211_),
    .Y(_03212_));
 sky130_fd_sc_hd__o21ai_4 _22909_ (.A1(_11463_),
    .A2(_03212_),
    .B1(net1485),
    .Y(_03213_));
 sky130_fd_sc_hd__o21ai_4 _22910_ (.A1(net266),
    .A2(_03089_),
    .B1(_03213_),
    .Y(_03214_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_322 ();
 sky130_fd_sc_hd__nand2_1 _22912_ (.A(_02119_),
    .B(_03214_),
    .Y(_03216_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_321 ();
 sky130_fd_sc_hd__nand2_1 _22914_ (.A(\gen_regfile_ff.register_file_i.rf_reg[142] ),
    .B(_02123_),
    .Y(_03218_));
 sky130_fd_sc_hd__nand2_1 _22915_ (.A(_03216_),
    .B(_03218_),
    .Y(_00526_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_320 ();
 sky130_fd_sc_hd__nand2_1 _22917_ (.A(_01682_),
    .B(net42),
    .Y(_03220_));
 sky130_fd_sc_hd__nand2_1 _22918_ (.A(\load_store_unit_i.rdata_offset_q[0] ),
    .B(_03220_),
    .Y(_03221_));
 sky130_fd_sc_hd__o21ai_0 _22919_ (.A1(\load_store_unit_i.rdata_offset_q[0] ),
    .A2(net51),
    .B1(_03221_),
    .Y(_03222_));
 sky130_fd_sc_hd__a221oi_1 _22920_ (.A1(\load_store_unit_i.rdata_q[23] ),
    .A2(_01672_),
    .B1(_01683_),
    .B2(\load_store_unit_i.rdata_q[31] ),
    .C1(\load_store_unit_i.data_type_q[2] ),
    .Y(_03223_));
 sky130_fd_sc_hd__a21oi_1 _22921_ (.A1(\load_store_unit_i.data_type_q[2] ),
    .A2(_03222_),
    .B1(_03223_),
    .Y(_03224_));
 sky130_fd_sc_hd__a21oi_1 _22922_ (.A1(\load_store_unit_i.rdata_offset_q[1] ),
    .A2(net56),
    .B1(_03224_),
    .Y(_03225_));
 sky130_fd_sc_hd__a22oi_1 _22923_ (.A1(net33),
    .A2(_02858_),
    .B1(_03224_),
    .B2(\load_store_unit_i.rdata_offset_q[1] ),
    .Y(_03226_));
 sky130_fd_sc_hd__o21ai_0 _22924_ (.A1(_01670_),
    .A2(_03225_),
    .B1(_03226_),
    .Y(_03227_));
 sky130_fd_sc_hd__a21oi_2 _22925_ (.A1(_01688_),
    .A2(_03227_),
    .B1(_02549_),
    .Y(_03228_));
 sky130_fd_sc_hd__nor2_1 _22926_ (.A(_02558_),
    .B(_02373_),
    .Y(_03229_));
 sky130_fd_sc_hd__a21oi_1 _22927_ (.A1(_01768_),
    .A2(_02558_),
    .B1(_03229_),
    .Y(_03230_));
 sky130_fd_sc_hd__o21ai_0 _22928_ (.A1(_02558_),
    .A2(_02368_),
    .B1(_02559_),
    .Y(_03231_));
 sky130_fd_sc_hd__nand2_1 _22929_ (.A(_01826_),
    .B(_03231_),
    .Y(_03232_));
 sky130_fd_sc_hd__o21ai_2 _22930_ (.A1(_01826_),
    .A2(_03230_),
    .B1(_03232_),
    .Y(_03233_));
 sky130_fd_sc_hd__o21ai_0 _22931_ (.A1(_02558_),
    .A2(_01825_),
    .B1(_02658_),
    .Y(_03234_));
 sky130_fd_sc_hd__nand2_1 _22932_ (.A(net295),
    .B(_03234_),
    .Y(_03235_));
 sky130_fd_sc_hd__o21ai_1 _22933_ (.A1(net295),
    .A2(_03233_),
    .B1(_03235_),
    .Y(_03236_));
 sky130_fd_sc_hd__nand3_1 _22934_ (.A(_09679_),
    .B(_09713_),
    .C(_02228_),
    .Y(_03237_));
 sky130_fd_sc_hd__o21ai_0 _22935_ (.A1(_09679_),
    .A2(_01902_),
    .B1(_03237_),
    .Y(_03238_));
 sky130_fd_sc_hd__a21oi_1 _22936_ (.A1(_09679_),
    .A2(_02233_),
    .B1(_09713_),
    .Y(_03239_));
 sky130_fd_sc_hd__a21oi_1 _22937_ (.A1(_02225_),
    .A2(_03238_),
    .B1(_03239_),
    .Y(_03240_));
 sky130_fd_sc_hd__a221oi_1 _22938_ (.A1(net721),
    .A2(_01929_),
    .B1(_03236_),
    .B2(_01734_),
    .C1(_03240_),
    .Y(_03241_));
 sky130_fd_sc_hd__nand2_1 _22939_ (.A(_03184_),
    .B(_03189_),
    .Y(_03242_));
 sky130_fd_sc_hd__nand4bb_4 _22940_ (.A_N(_02672_),
    .B_N(_02678_),
    .C(_02748_),
    .D(_02822_),
    .Y(_03243_));
 sky130_fd_sc_hd__a21bo_1 _22941_ (.A1(_02823_),
    .A2(_02825_),
    .B1_N(_02822_),
    .X(_03244_));
 sky130_fd_sc_hd__a311oi_4 _22942_ (.A1(_02996_),
    .A2(_03243_),
    .A3(_03244_),
    .B1(_03188_),
    .C1(_02964_),
    .Y(_03245_));
 sky130_fd_sc_hd__o21a_1 _22943_ (.A1(_03242_),
    .A2(_03245_),
    .B1(_03185_),
    .X(_03246_));
 sky130_fd_sc_hd__maj3_2 _22944_ (.A(_03093_),
    .B(_03180_),
    .C(_03181_),
    .X(_03247_));
 sky130_fd_sc_hd__a21o_1 _22945_ (.A1(_03157_),
    .A2(_03176_),
    .B1(_03158_),
    .X(_03248_));
 sky130_fd_sc_hd__o21ai_4 _22946_ (.A1(_03157_),
    .A2(_03176_),
    .B1(_03248_),
    .Y(_03249_));
 sky130_fd_sc_hd__nand2_2 _22947_ (.A(_03121_),
    .B(_03122_),
    .Y(_03250_));
 sky130_fd_sc_hd__xnor2_1 _22948_ (.A(net857),
    .B(_03250_),
    .Y(_03251_));
 sky130_fd_sc_hd__nor3_2 _22949_ (.A(_03042_),
    .B(_03044_),
    .C(_03251_),
    .Y(_03252_));
 sky130_fd_sc_hd__a22o_2 _22950_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[61] ),
    .A2(net322),
    .B1(_03043_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .X(_03253_));
 sky130_fd_sc_hd__nand2_1 _22951_ (.A(_03100_),
    .B(_03253_),
    .Y(_03254_));
 sky130_fd_sc_hd__o21ai_0 _22952_ (.A1(_02032_),
    .A2(_03253_),
    .B1(_03041_),
    .Y(_03255_));
 sky130_fd_sc_hd__mux2i_1 _22953_ (.A0(_03254_),
    .A1(_03255_),
    .S(_03250_),
    .Y(_03256_));
 sky130_fd_sc_hd__a21o_1 _22954_ (.A1(_03045_),
    .A2(_03256_),
    .B1(_03123_),
    .X(_03257_));
 sky130_fd_sc_hd__nor2_1 _22955_ (.A(_03253_),
    .B(_03045_),
    .Y(_03258_));
 sky130_fd_sc_hd__nor2_1 _22956_ (.A(net949),
    .B(_03258_),
    .Y(_03259_));
 sky130_fd_sc_hd__a21oi_1 _22957_ (.A1(net984),
    .A2(_03250_),
    .B1(_03259_),
    .Y(_03260_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_319 ();
 sky130_fd_sc_hd__nand2_1 _22959_ (.A(_03253_),
    .B(_03045_),
    .Y(_03262_));
 sky130_fd_sc_hd__o221ai_4 _22960_ (.A1(_03102_),
    .A2(_03250_),
    .B1(_03260_),
    .B2(_03100_),
    .C1(_03262_),
    .Y(_03263_));
 sky130_fd_sc_hd__o21ai_4 _22961_ (.A1(_03252_),
    .A2(_03257_),
    .B1(_03263_),
    .Y(_03264_));
 sky130_fd_sc_hd__nor2_8 _22962_ (.A(_03113_),
    .B(net1064),
    .Y(_03265_));
 sky130_fd_sc_hd__nand2_1 _22963_ (.A(_02016_),
    .B(_03265_),
    .Y(_03266_));
 sky130_fd_sc_hd__nand2_1 _22964_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[47] ),
    .B(net316),
    .Y(_03267_));
 sky130_fd_sc_hd__o21ai_1 _22965_ (.A1(_10727_),
    .A2(net316),
    .B1(_03267_),
    .Y(_03268_));
 sky130_fd_sc_hd__a22oi_4 _22966_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[63] ),
    .A2(_01702_),
    .B1(_03268_),
    .B2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .Y(_03269_));
 sky130_fd_sc_hd__a31o_1 _22967_ (.A1(_08179_),
    .A2(_09653_),
    .A3(_09656_),
    .B1(_01720_),
    .X(_03270_));
 sky130_fd_sc_hd__or3_4 _22968_ (.A(_09669_),
    .B(_09674_),
    .C(_03270_),
    .X(_03271_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_318 ();
 sky130_fd_sc_hd__nand4_4 _22970_ (.A(_10676_),
    .B(_10683_),
    .C(_10690_),
    .D(_01720_),
    .Y(_03273_));
 sky130_fd_sc_hd__nand2_4 _22971_ (.A(_03271_),
    .B(_03273_),
    .Y(_03274_));
 sky130_fd_sc_hd__nand2_1 _22972_ (.A(_02032_),
    .B(_03274_),
    .Y(_03275_));
 sky130_fd_sc_hd__xor3_4 _22973_ (.A(_03266_),
    .B(_03269_),
    .C(_03275_),
    .X(_03276_));
 sky130_fd_sc_hd__nor3_1 _22974_ (.A(net951),
    .B(_03107_),
    .C(_03119_),
    .Y(_03277_));
 sky130_fd_sc_hd__maj3_1 _22975_ (.A(_03137_),
    .B(_03138_),
    .C(_03139_),
    .X(_03278_));
 sky130_fd_sc_hd__o211a_1 _22976_ (.A1(_03102_),
    .A2(_03277_),
    .B1(_03122_),
    .C1(_03278_),
    .X(_03279_));
 sky130_fd_sc_hd__a311oi_2 _22977_ (.A1(net984),
    .A2(_03041_),
    .A3(_03122_),
    .B1(_03278_),
    .C1(_03277_),
    .Y(_03280_));
 sky130_fd_sc_hd__nor2_1 _22978_ (.A(_03279_),
    .B(_03280_),
    .Y(_03281_));
 sky130_fd_sc_hd__xnor2_4 _22979_ (.A(_03276_),
    .B(_03281_),
    .Y(_03282_));
 sky130_fd_sc_hd__maj3_2 _22980_ (.A(_03148_),
    .B(_03153_),
    .C(_03156_),
    .X(_03283_));
 sky130_fd_sc_hd__xnor2_2 _22981_ (.A(_03283_),
    .B(_03132_),
    .Y(_03284_));
 sky130_fd_sc_hd__xnor3_2 _22982_ (.A(_03264_),
    .B(_03282_),
    .C(_03284_),
    .X(_03285_));
 sky130_fd_sc_hd__nor2_1 _22983_ (.A(net1286),
    .B(_02692_),
    .Y(_03286_));
 sky130_fd_sc_hd__nor2_1 _22984_ (.A(net1216),
    .B(net1277),
    .Y(_03287_));
 sky130_fd_sc_hd__nor2_1 _22985_ (.A(_02289_),
    .B(_03142_),
    .Y(_03288_));
 sky130_fd_sc_hd__xor3_1 _22986_ (.A(_03286_),
    .B(_03287_),
    .C(_03288_),
    .X(_03289_));
 sky130_fd_sc_hd__maj3_1 _22987_ (.A(_03144_),
    .B(_03145_),
    .C(_03146_),
    .X(_03290_));
 sky130_fd_sc_hd__nor2_1 _22988_ (.A(_02088_),
    .B(_03097_),
    .Y(_03291_));
 sky130_fd_sc_hd__nor2_1 _22989_ (.A(_02010_),
    .B(_03100_),
    .Y(_03292_));
 sky130_fd_sc_hd__nor2_1 _22990_ (.A(_02292_),
    .B(net1336),
    .Y(_03293_));
 sky130_fd_sc_hd__xor3_4 _22991_ (.A(_03291_),
    .B(_03292_),
    .C(_03293_),
    .X(_03294_));
 sky130_fd_sc_hd__xor3_1 _22992_ (.A(_03289_),
    .B(_03290_),
    .C(_03294_),
    .X(_03295_));
 sky130_fd_sc_hd__inv_1 _22993_ (.A(_03295_),
    .Y(_03296_));
 sky130_fd_sc_hd__maj3_1 _22994_ (.A(_03169_),
    .B(_03173_),
    .C(_03174_),
    .X(_03297_));
 sky130_fd_sc_hd__maj3_1 _22995_ (.A(_03136_),
    .B(_03141_),
    .C(_03147_),
    .X(_03298_));
 sky130_fd_sc_hd__xnor2_2 _22996_ (.A(_03297_),
    .B(_03298_),
    .Y(_03299_));
 sky130_fd_sc_hd__xnor2_2 _22997_ (.A(_03296_),
    .B(_03299_),
    .Y(_03300_));
 sky130_fd_sc_hd__nor2_1 _22998_ (.A(_03168_),
    .B(_03175_),
    .Y(_03301_));
 sky130_fd_sc_hd__maj3_2 _22999_ (.A(_03166_),
    .B(_03164_),
    .C(_03163_),
    .X(_03302_));
 sky130_fd_sc_hd__nand2_1 _23000_ (.A(_02436_),
    .B(_02727_),
    .Y(_03303_));
 sky130_fd_sc_hd__nand2b_1 _23001_ (.A_N(_02513_),
    .B(_02918_),
    .Y(_03304_));
 sky130_fd_sc_hd__or2_0 _23002_ (.A(net1069),
    .B(_02622_),
    .X(_03305_));
 sky130_fd_sc_hd__xor3_1 _23003_ (.A(_03303_),
    .B(_03304_),
    .C(_03305_),
    .X(_03306_));
 sky130_fd_sc_hd__maj3_1 _23004_ (.A(_03170_),
    .B(_03171_),
    .C(_03172_),
    .X(_03307_));
 sky130_fd_sc_hd__xnor3_1 _23005_ (.A(_03302_),
    .B(_03306_),
    .C(_03307_),
    .X(_03308_));
 sky130_fd_sc_hd__nand4_4 _23006_ (.A(_10700_),
    .B(_10707_),
    .C(_10720_),
    .D(net321),
    .Y(_03309_));
 sky130_fd_sc_hd__o21a_4 _23007_ (.A1(_09707_),
    .A2(net322),
    .B1(_03309_),
    .X(_03310_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_317 ();
 sky130_fd_sc_hd__nand2_1 _23009_ (.A(_01998_),
    .B(_03310_),
    .Y(_03312_));
 sky130_fd_sc_hd__a21o_4 _23010_ (.A1(net1163),
    .A2(net322),
    .B1(_03160_),
    .X(_03313_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_316 ();
 sky130_fd_sc_hd__nor2_1 _23012_ (.A(net790),
    .B(_03313_),
    .Y(_03315_));
 sky130_fd_sc_hd__xnor2_1 _23013_ (.A(_03312_),
    .B(_03315_),
    .Y(_03316_));
 sky130_fd_sc_hd__nor2_1 _23014_ (.A(net1060),
    .B(_02932_),
    .Y(_03317_));
 sky130_fd_sc_hd__nand2_1 _23015_ (.A(_02440_),
    .B(_02774_),
    .Y(_03318_));
 sky130_fd_sc_hd__nor2_1 _23016_ (.A(net781),
    .B(_03165_),
    .Y(_03319_));
 sky130_fd_sc_hd__xnor3_1 _23017_ (.A(_03317_),
    .B(_03318_),
    .C(_03319_),
    .X(_03320_));
 sky130_fd_sc_hd__xor2_2 _23018_ (.A(_03316_),
    .B(_03320_),
    .X(_03321_));
 sky130_fd_sc_hd__nor2_2 _23019_ (.A(_03162_),
    .B(_03167_),
    .Y(_03322_));
 sky130_fd_sc_hd__xnor3_2 _23020_ (.A(_03308_),
    .B(_03321_),
    .C(_03322_),
    .X(_03323_));
 sky130_fd_sc_hd__xor2_2 _23021_ (.A(_03301_),
    .B(_03323_),
    .X(_03324_));
 sky130_fd_sc_hd__xnor2_2 _23022_ (.A(_03300_),
    .B(_03324_),
    .Y(_03325_));
 sky130_fd_sc_hd__xor2_4 _23023_ (.A(_03285_),
    .B(_03325_),
    .X(_03326_));
 sky130_fd_sc_hd__xnor2_4 _23024_ (.A(_03249_),
    .B(_03326_),
    .Y(_03327_));
 sky130_fd_sc_hd__o21bai_1 _23025_ (.A1(_03131_),
    .A2(_03132_),
    .B1_N(_03096_),
    .Y(_03328_));
 sky130_fd_sc_hd__and2_0 _23026_ (.A(_03094_),
    .B(_03328_),
    .X(_03329_));
 sky130_fd_sc_hd__nor3b_2 _23027_ (.A(_03131_),
    .B(_03132_),
    .C_N(_03096_),
    .Y(_03330_));
 sky130_fd_sc_hd__o32ai_2 _23028_ (.A1(_03178_),
    .A2(_03329_),
    .A3(_03330_),
    .B1(_03328_),
    .B2(_03094_),
    .Y(_03331_));
 sky130_fd_sc_hd__nand2_1 _23029_ (.A(_03094_),
    .B(_03330_),
    .Y(_03332_));
 sky130_fd_sc_hd__o211ai_1 _23030_ (.A1(_03094_),
    .A2(_03330_),
    .B1(_03328_),
    .C1(_03178_),
    .Y(_03333_));
 sky130_fd_sc_hd__a21oi_2 _23031_ (.A1(_03332_),
    .A2(_03333_),
    .B1(net903),
    .Y(_03334_));
 sky130_fd_sc_hd__nor2_1 _23032_ (.A(_03096_),
    .B(_03134_),
    .Y(_03335_));
 sky130_fd_sc_hd__nor2_1 _23033_ (.A(_03094_),
    .B(_03178_),
    .Y(_03336_));
 sky130_fd_sc_hd__nand2_1 _23034_ (.A(_03094_),
    .B(_03178_),
    .Y(_03337_));
 sky130_fd_sc_hd__nand2_1 _23035_ (.A(_03096_),
    .B(_03134_),
    .Y(_03338_));
 sky130_fd_sc_hd__o2bb2ai_1 _23036_ (.A1_N(_03335_),
    .A2_N(_03336_),
    .B1(_03337_),
    .B2(_03338_),
    .Y(_03339_));
 sky130_fd_sc_hd__a211oi_4 _23037_ (.A1(_03331_),
    .A2(net903),
    .B1(_03334_),
    .C1(_03339_),
    .Y(_03340_));
 sky130_fd_sc_hd__xor2_4 _23038_ (.A(_03327_),
    .B(_03340_),
    .X(_03341_));
 sky130_fd_sc_hd__xor2_4 _23039_ (.A(_03247_),
    .B(_03341_),
    .X(_03342_));
 sky130_fd_sc_hd__xnor2_4 _23040_ (.A(_03246_),
    .B(_03342_),
    .Y(_03343_));
 sky130_fd_sc_hd__o21ai_0 _23041_ (.A1(net441),
    .A2(_01698_),
    .B1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[47] ),
    .Y(_03344_));
 sky130_fd_sc_hd__o311a_1 _23042_ (.A1(net441),
    .A2(_01698_),
    .A3(_03343_),
    .B1(_03344_),
    .C1(net312),
    .X(_03345_));
 sky130_fd_sc_hd__a21oi_2 _23043_ (.A1(_08290_),
    .A2(_03241_),
    .B1(_03345_),
    .Y(_03346_));
 sky130_fd_sc_hd__nor3_1 _23044_ (.A(_11486_),
    .B(_02646_),
    .C(_03346_),
    .Y(_03347_));
 sky130_fd_sc_hd__a21oi_4 _23045_ (.A1(_02646_),
    .A2(_03228_),
    .B1(_03347_),
    .Y(_03348_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_315 ();
 sky130_fd_sc_hd__nand2_1 _23047_ (.A(_02119_),
    .B(_03348_),
    .Y(_03350_));
 sky130_fd_sc_hd__nand2_1 _23048_ (.A(\gen_regfile_ff.register_file_i.rf_reg[143] ),
    .B(_02123_),
    .Y(_03351_));
 sky130_fd_sc_hd__nand2_1 _23049_ (.A(_03350_),
    .B(_03351_),
    .Y(_00527_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_314 ();
 sky130_fd_sc_hd__nor2_1 _23051_ (.A(_03091_),
    .B(_03183_),
    .Y(_03353_));
 sky130_fd_sc_hd__nor2_2 _23052_ (.A(_03247_),
    .B(_03341_),
    .Y(_03354_));
 sky130_fd_sc_hd__nor2_2 _23053_ (.A(_03354_),
    .B(_03353_),
    .Y(_03355_));
 sky130_fd_sc_hd__nand2_1 _23054_ (.A(_03247_),
    .B(_03341_),
    .Y(_03356_));
 sky130_fd_sc_hd__a21oi_4 _23055_ (.A1(_03185_),
    .A2(_03356_),
    .B1(_03354_),
    .Y(_03357_));
 sky130_fd_sc_hd__a31oi_4 _23056_ (.A1(_03187_),
    .A2(_03190_),
    .A3(_03355_),
    .B1(_03357_),
    .Y(_03358_));
 sky130_fd_sc_hd__maj3_1 _23057_ (.A(_03308_),
    .B(_03321_),
    .C(_03322_),
    .X(_03359_));
 sky130_fd_sc_hd__nand2_1 _23058_ (.A(_02440_),
    .B(_03015_),
    .Y(_03360_));
 sky130_fd_sc_hd__nand2_1 _23059_ (.A(_02436_),
    .B(_02774_),
    .Y(_03361_));
 sky130_fd_sc_hd__nand2_1 _23060_ (.A(_02160_),
    .B(_03017_),
    .Y(_03362_));
 sky130_fd_sc_hd__xnor3_1 _23061_ (.A(_03360_),
    .B(_03361_),
    .C(_03362_),
    .X(_03363_));
 sky130_fd_sc_hd__nor2_1 _23062_ (.A(net1172),
    .B(_03313_),
    .Y(_03364_));
 sky130_fd_sc_hd__nor3_2 _23063_ (.A(_08163_),
    .B(_10697_),
    .C(_10699_),
    .Y(_03365_));
 sky130_fd_sc_hd__and3_2 _23064_ (.A(net698),
    .B(_10703_),
    .C(_10706_),
    .X(_03366_));
 sky130_fd_sc_hd__or4_4 _23065_ (.A(_10710_),
    .B(_10713_),
    .C(_10716_),
    .D(_10719_),
    .X(_03367_));
 sky130_fd_sc_hd__nor3_4 _23066_ (.A(_08294_),
    .B(_08265_),
    .C(_08399_),
    .Y(_03368_));
 sky130_fd_sc_hd__o31a_4 _23067_ (.A1(_03365_),
    .A2(_03366_),
    .A3(_03367_),
    .B1(_03368_),
    .X(_03369_));
 sky130_fd_sc_hd__nand2_8 _23068_ (.A(net322),
    .B(_03369_),
    .Y(_03370_));
 sky130_fd_sc_hd__nand4_1 _23069_ (.A(net781),
    .B(net1287),
    .C(_03310_),
    .D(_03370_),
    .Y(_03371_));
 sky130_fd_sc_hd__o31ai_1 _23070_ (.A1(net1287),
    .A2(_03364_),
    .A3(_03370_),
    .B1(_03371_),
    .Y(_03372_));
 sky130_fd_sc_hd__o21ai_4 _23071_ (.A1(_09707_),
    .A2(net322),
    .B1(_03309_),
    .Y(_03373_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_313 ();
 sky130_fd_sc_hd__o31ai_4 _23073_ (.A1(_03365_),
    .A2(_03366_),
    .A3(_03367_),
    .B1(_03368_),
    .Y(_03375_));
 sky130_fd_sc_hd__nor2_8 _23074_ (.A(_01712_),
    .B(net1205),
    .Y(_03376_));
 sky130_fd_sc_hd__nor3_2 _23075_ (.A(net791),
    .B(_03373_),
    .C(_03376_),
    .Y(_03377_));
 sky130_fd_sc_hd__or3_4 _23076_ (.A(_08294_),
    .B(_08265_),
    .C(_08399_),
    .X(_03378_));
 sky130_fd_sc_hd__nand3b_2 _23077_ (.A_N(_03378_),
    .B(net322),
    .C(_10721_),
    .Y(_03379_));
 sky130_fd_sc_hd__nor2_1 _23078_ (.A(_02014_),
    .B(_03379_),
    .Y(_03380_));
 sky130_fd_sc_hd__nor4_2 _23079_ (.A(net781),
    .B(_03313_),
    .C(_03380_),
    .D(_03377_),
    .Y(_03381_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_312 ();
 sky130_fd_sc_hd__nand2_1 _23081_ (.A(net1287),
    .B(_03310_),
    .Y(_03383_));
 sky130_fd_sc_hd__a311oi_4 _23082_ (.A1(_10700_),
    .A2(_10707_),
    .A3(_10720_),
    .B1(net320),
    .C1(_03378_),
    .Y(_03384_));
 sky130_fd_sc_hd__nor3_1 _23083_ (.A(_03161_),
    .B(_03383_),
    .C(_03384_),
    .Y(_03385_));
 sky130_fd_sc_hd__nor3_1 _23084_ (.A(_03373_),
    .B(_03161_),
    .C(net792),
    .Y(_03386_));
 sky130_fd_sc_hd__o21a_1 _23085_ (.A1(_03364_),
    .A2(_03386_),
    .B1(_01998_),
    .X(_03387_));
 sky130_fd_sc_hd__a2111oi_2 _23086_ (.A1(net1178),
    .A2(_03372_),
    .B1(_03387_),
    .C1(_03385_),
    .D1(_03381_),
    .Y(_03388_));
 sky130_fd_sc_hd__xnor2_1 _23087_ (.A(_03388_),
    .B(_03363_),
    .Y(_03389_));
 sky130_fd_sc_hd__nand2_1 _23088_ (.A(_03316_),
    .B(_03320_),
    .Y(_03390_));
 sky130_fd_sc_hd__nor4_1 _23089_ (.A(net1172),
    .B(_02080_),
    .C(_02936_),
    .D(_03165_),
    .Y(_03391_));
 sky130_fd_sc_hd__o22ai_1 _23090_ (.A1(_02080_),
    .A2(_02936_),
    .B1(_03165_),
    .B2(net781),
    .Y(_03392_));
 sky130_fd_sc_hd__o21ai_1 _23091_ (.A1(_03317_),
    .A2(_03391_),
    .B1(_03392_),
    .Y(_03393_));
 sky130_fd_sc_hd__or3_1 _23092_ (.A(net1069),
    .B(_02723_),
    .C(_02725_),
    .X(_03394_));
 sky130_fd_sc_hd__or2_0 _23093_ (.A(net1277),
    .B(_02513_),
    .X(_03395_));
 sky130_fd_sc_hd__or2_0 _23094_ (.A(net1031),
    .B(_02622_),
    .X(_03396_));
 sky130_fd_sc_hd__xor3_1 _23095_ (.A(_03394_),
    .B(_03396_),
    .C(_03395_),
    .X(_03397_));
 sky130_fd_sc_hd__maj3_1 _23096_ (.A(_03303_),
    .B(_03304_),
    .C(_03305_),
    .X(_03398_));
 sky130_fd_sc_hd__xnor3_1 _23097_ (.A(_03393_),
    .B(_03397_),
    .C(_03398_),
    .X(_03399_));
 sky130_fd_sc_hd__xor2_1 _23098_ (.A(_03390_),
    .B(_03399_),
    .X(_03400_));
 sky130_fd_sc_hd__xnor2_1 _23099_ (.A(_03389_),
    .B(_03400_),
    .Y(_03401_));
 sky130_fd_sc_hd__nand2_1 _23100_ (.A(_03302_),
    .B(_03307_),
    .Y(_03402_));
 sky130_fd_sc_hd__nor2_1 _23101_ (.A(_03302_),
    .B(_03307_),
    .Y(_03403_));
 sky130_fd_sc_hd__a21oi_1 _23102_ (.A1(_03306_),
    .A2(_03402_),
    .B1(_03403_),
    .Y(_03404_));
 sky130_fd_sc_hd__nand2_1 _23103_ (.A(net1180),
    .B(_02889_),
    .Y(_03405_));
 sky130_fd_sc_hd__nand2_1 _23104_ (.A(_02421_),
    .B(_02589_),
    .Y(_03406_));
 sky130_fd_sc_hd__and4_4 _23105_ (.A(_02688_),
    .B(_02689_),
    .C(_02690_),
    .D(_02691_),
    .X(_03407_));
 sky130_fd_sc_hd__nand2_1 _23106_ (.A(_02301_),
    .B(_03407_),
    .Y(_03408_));
 sky130_fd_sc_hd__xnor3_1 _23107_ (.A(_03405_),
    .B(_03406_),
    .C(_03408_),
    .X(_03409_));
 sky130_fd_sc_hd__nor2_1 _23108_ (.A(_02292_),
    .B(_03097_),
    .Y(_03410_));
 sky130_fd_sc_hd__nor2_1 _23109_ (.A(_02010_),
    .B(_03119_),
    .Y(_03411_));
 sky130_fd_sc_hd__nor2_1 _23110_ (.A(_02088_),
    .B(_03100_),
    .Y(_03412_));
 sky130_fd_sc_hd__xor3_2 _23111_ (.A(_03410_),
    .B(_03411_),
    .C(_03412_),
    .X(_03413_));
 sky130_fd_sc_hd__maj3_1 _23112_ (.A(_03286_),
    .B(_03287_),
    .C(_03288_),
    .X(_03414_));
 sky130_fd_sc_hd__xor3_2 _23113_ (.A(_03409_),
    .B(_03413_),
    .C(_03414_),
    .X(_03415_));
 sky130_fd_sc_hd__maj3_1 _23114_ (.A(_03289_),
    .B(_03290_),
    .C(_03294_),
    .X(_03416_));
 sky130_fd_sc_hd__xnor2_1 _23115_ (.A(_03415_),
    .B(_03416_),
    .Y(_03417_));
 sky130_fd_sc_hd__xnor2_1 _23116_ (.A(_03404_),
    .B(_03417_),
    .Y(_03418_));
 sky130_fd_sc_hd__xnor2_1 _23117_ (.A(_03401_),
    .B(_03418_),
    .Y(_03419_));
 sky130_fd_sc_hd__xnor2_2 _23118_ (.A(_03359_),
    .B(_03419_),
    .Y(_03420_));
 sky130_fd_sc_hd__maj3_1 _23119_ (.A(_03297_),
    .B(_03296_),
    .C(_03298_),
    .X(_03421_));
 sky130_fd_sc_hd__o211ai_2 _23120_ (.A1(_03252_),
    .A2(_03257_),
    .B1(_03282_),
    .C1(_03263_),
    .Y(_03422_));
 sky130_fd_sc_hd__nand3_2 _23121_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .B(_08235_),
    .C(_08216_),
    .Y(_03423_));
 sky130_fd_sc_hd__nor3_4 _23122_ (.A(_08294_),
    .B(_13439_),
    .C(_03423_),
    .Y(_03424_));
 sky130_fd_sc_hd__a22o_1 _23123_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .A2(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ),
    .B1(_03424_),
    .B2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[48] ),
    .X(_03425_));
 sky130_fd_sc_hd__a221oi_2 _23124_ (.A1(net699),
    .A2(_01712_),
    .B1(_03271_),
    .B2(_03273_),
    .C1(net1268),
    .Y(_03426_));
 sky130_fd_sc_hd__nor4b_2 _23125_ (.A(_13439_),
    .B(_01968_),
    .C(_13440_),
    .D_N(_13357_),
    .Y(_03427_));
 sky130_fd_sc_hd__and4_4 _23126_ (.A(_10676_),
    .B(_10683_),
    .C(_10690_),
    .D(_03427_),
    .X(_03428_));
 sky130_fd_sc_hd__o221ai_4 _23127_ (.A1(_01711_),
    .A2(net320),
    .B1(_01715_),
    .B2(_01716_),
    .C1(_03428_),
    .Y(_03429_));
 sky130_fd_sc_hd__mux2i_1 _23128_ (.A0(_01982_),
    .A1(_03426_),
    .S(_03429_),
    .Y(_03430_));
 sky130_fd_sc_hd__xnor2_1 _23129_ (.A(_03425_),
    .B(_03430_),
    .Y(_03431_));
 sky130_fd_sc_hd__maj3_1 _23130_ (.A(_03266_),
    .B(_03269_),
    .C(_03275_),
    .X(_03432_));
 sky130_fd_sc_hd__maj3_1 _23131_ (.A(_03291_),
    .B(_03292_),
    .C(_03293_),
    .X(_03433_));
 sky130_fd_sc_hd__xnor3_4 _23132_ (.A(_03431_),
    .B(_03432_),
    .C(_03433_),
    .X(_03434_));
 sky130_fd_sc_hd__o21bai_1 _23133_ (.A1(_03276_),
    .A2(_03280_),
    .B1_N(_03279_),
    .Y(_03435_));
 sky130_fd_sc_hd__xor2_1 _23134_ (.A(_03434_),
    .B(_03435_),
    .X(_03436_));
 sky130_fd_sc_hd__xnor2_2 _23135_ (.A(_03436_),
    .B(_03370_),
    .Y(_03437_));
 sky130_fd_sc_hd__xnor2_1 _23136_ (.A(_03422_),
    .B(_03437_),
    .Y(_03438_));
 sky130_fd_sc_hd__xnor2_1 _23137_ (.A(_03421_),
    .B(_03438_),
    .Y(_03439_));
 sky130_fd_sc_hd__nand2_1 _23138_ (.A(_03300_),
    .B(_03323_),
    .Y(_03440_));
 sky130_fd_sc_hd__nor2_1 _23139_ (.A(_03300_),
    .B(_03323_),
    .Y(_03441_));
 sky130_fd_sc_hd__a21o_1 _23140_ (.A1(_03301_),
    .A2(_03440_),
    .B1(_03441_),
    .X(_03442_));
 sky130_fd_sc_hd__xnor2_1 _23141_ (.A(_03439_),
    .B(_03442_),
    .Y(_03443_));
 sky130_fd_sc_hd__xnor2_2 _23142_ (.A(_03420_),
    .B(_03443_),
    .Y(_03444_));
 sky130_fd_sc_hd__xnor2_1 _23143_ (.A(_03264_),
    .B(_03282_),
    .Y(_03445_));
 sky130_fd_sc_hd__nor2_1 _23144_ (.A(_03132_),
    .B(_03445_),
    .Y(_03446_));
 sky130_fd_sc_hd__nand2_1 _23145_ (.A(_03132_),
    .B(_03445_),
    .Y(_03447_));
 sky130_fd_sc_hd__o21a_1 _23146_ (.A1(_03283_),
    .A2(_03446_),
    .B1(_03447_),
    .X(_03448_));
 sky130_fd_sc_hd__nor2_1 _23147_ (.A(_03249_),
    .B(_03325_),
    .Y(_03449_));
 sky130_fd_sc_hd__nand2_1 _23148_ (.A(_03249_),
    .B(_03325_),
    .Y(_03450_));
 sky130_fd_sc_hd__o21ai_2 _23149_ (.A1(_03285_),
    .A2(_03449_),
    .B1(_03450_),
    .Y(_03451_));
 sky130_fd_sc_hd__xor2_2 _23150_ (.A(_03448_),
    .B(_03451_),
    .X(_03452_));
 sky130_fd_sc_hd__xnor2_4 _23151_ (.A(_03444_),
    .B(_03452_),
    .Y(_03453_));
 sky130_fd_sc_hd__a21oi_1 _23152_ (.A1(_03327_),
    .A2(_03337_),
    .B1(_03177_),
    .Y(_03454_));
 sky130_fd_sc_hd__o21a_1 _23153_ (.A1(_03177_),
    .A2(_03336_),
    .B1(_03337_),
    .X(_03455_));
 sky130_fd_sc_hd__a21oi_1 _23154_ (.A1(_03338_),
    .A2(_03455_),
    .B1(_03327_),
    .Y(_03456_));
 sky130_fd_sc_hd__o32ai_2 _23155_ (.A1(_03336_),
    .A2(_03335_),
    .A3(_03327_),
    .B1(_03455_),
    .B2(_03338_),
    .Y(_03457_));
 sky130_fd_sc_hd__a211o_2 _23156_ (.A1(_03454_),
    .A2(_03328_),
    .B1(_03457_),
    .C1(_03456_),
    .X(_03458_));
 sky130_fd_sc_hd__xnor2_4 _23157_ (.A(_03453_),
    .B(_03458_),
    .Y(_03459_));
 sky130_fd_sc_hd__xor2_4 _23158_ (.A(_03358_),
    .B(_03459_),
    .X(_03460_));
 sky130_fd_sc_hd__nor2_1 _23159_ (.A(_01698_),
    .B(_03460_),
    .Y(_03461_));
 sky130_fd_sc_hd__a21oi_2 _23160_ (.A1(_01698_),
    .A2(_01727_),
    .B1(_03461_),
    .Y(_03462_));
 sky130_fd_sc_hd__mux2i_2 _23161_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[48] ),
    .A1(_03462_),
    .S(_08100_),
    .Y(_03463_));
 sky130_fd_sc_hd__nor2_1 _23162_ (.A(net295),
    .B(_03234_),
    .Y(_03464_));
 sky130_fd_sc_hd__a211oi_2 _23163_ (.A1(net295),
    .A2(_03233_),
    .B1(_03464_),
    .C1(_01761_),
    .Y(_03465_));
 sky130_fd_sc_hd__nand3_1 _23164_ (.A(_09825_),
    .B(_09859_),
    .C(_02228_),
    .Y(_03466_));
 sky130_fd_sc_hd__o21ai_0 _23165_ (.A1(_09859_),
    .A2(_01902_),
    .B1(_03466_),
    .Y(_03467_));
 sky130_fd_sc_hd__a21oi_1 _23166_ (.A1(_09859_),
    .A2(_02233_),
    .B1(_09825_),
    .Y(_03468_));
 sky130_fd_sc_hd__a21oi_1 _23167_ (.A1(_02225_),
    .A2(_03467_),
    .B1(_03468_),
    .Y(_03469_));
 sky130_fd_sc_hd__a2111oi_0 _23168_ (.A1(net157),
    .A2(_01929_),
    .B1(_03465_),
    .C1(_03469_),
    .D1(net314),
    .Y(_03470_));
 sky130_fd_sc_hd__a21oi_1 _23169_ (.A1(net314),
    .A2(_03463_),
    .B1(_03470_),
    .Y(_03471_));
 sky130_fd_sc_hd__nand2_1 _23170_ (.A(_11503_),
    .B(net265),
    .Y(_03472_));
 sky130_fd_sc_hd__mux4_1 _23171_ (.A0(net34),
    .A1(net27),
    .A2(\load_store_unit_i.rdata_q[24] ),
    .A3(net57),
    .S0(\load_store_unit_i.rdata_offset_q[1] ),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .X(_03473_));
 sky130_fd_sc_hd__nand2_1 _23172_ (.A(\load_store_unit_i.rdata_offset_q[1] ),
    .B(net56),
    .Y(_03474_));
 sky130_fd_sc_hd__nand2_1 _23173_ (.A(_03220_),
    .B(_03474_),
    .Y(_03475_));
 sky130_fd_sc_hd__nand2_1 _23174_ (.A(\load_store_unit_i.rdata_offset_q[0] ),
    .B(_03475_),
    .Y(_03476_));
 sky130_fd_sc_hd__o21ai_1 _23175_ (.A1(\load_store_unit_i.rdata_offset_q[0] ),
    .A2(_02547_),
    .B1(_03476_),
    .Y(_03477_));
 sky130_fd_sc_hd__a31oi_4 _23176_ (.A1(\load_store_unit_i.data_type_q[2] ),
    .A2(\load_store_unit_i.data_sign_ext_q ),
    .A3(_03477_),
    .B1(_02549_),
    .Y(_03478_));
 sky130_fd_sc_hd__nand2_4 _23177_ (.A(_02646_),
    .B(_03478_),
    .Y(_03479_));
 sky130_fd_sc_hd__a21oi_2 _23178_ (.A1(_01674_),
    .A2(_03473_),
    .B1(_03479_),
    .Y(_03480_));
 sky130_fd_sc_hd__o21bai_4 _23179_ (.A1(_03471_),
    .A2(_03472_),
    .B1_N(_03480_),
    .Y(_03481_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_311 ();
 sky130_fd_sc_hd__nand2_1 _23181_ (.A(\gen_regfile_ff.register_file_i.rf_reg[144] ),
    .B(_02123_),
    .Y(_03483_));
 sky130_fd_sc_hd__o21ai_0 _23182_ (.A1(_02123_),
    .A2(_03481_),
    .B1(_03483_),
    .Y(_00528_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_310 ();
 sky130_fd_sc_hd__mux4_1 _23184_ (.A0(net35),
    .A1(net38),
    .A2(\load_store_unit_i.rdata_q[25] ),
    .A3(net58),
    .S0(\load_store_unit_i.rdata_offset_q[1] ),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .X(_03485_));
 sky130_fd_sc_hd__nand2_1 _23185_ (.A(_01674_),
    .B(_03485_),
    .Y(_03486_));
 sky130_fd_sc_hd__a21oi_1 _23186_ (.A1(net857),
    .A2(_02297_),
    .B1(_01984_),
    .Y(_03487_));
 sky130_fd_sc_hd__inv_1 _23187_ (.A(_01710_),
    .Y(_03488_));
 sky130_fd_sc_hd__o22ai_1 _23188_ (.A1(_01998_),
    .A2(net887),
    .B1(_03487_),
    .B2(_03488_),
    .Y(_03489_));
 sky130_fd_sc_hd__nor2_1 _23189_ (.A(net984),
    .B(_02034_),
    .Y(_03490_));
 sky130_fd_sc_hd__a21oi_1 _23190_ (.A1(net984),
    .A2(_02297_),
    .B1(_03490_),
    .Y(_03491_));
 sky130_fd_sc_hd__o22ai_1 _23191_ (.A1(_02032_),
    .A2(_02028_),
    .B1(_03491_),
    .B2(_01710_),
    .Y(_03492_));
 sky130_fd_sc_hd__a21oi_2 _23192_ (.A1(_02032_),
    .A2(_03489_),
    .B1(_03492_),
    .Y(_03493_));
 sky130_fd_sc_hd__xnor2_2 _23193_ (.A(_02018_),
    .B(_03493_),
    .Y(_03494_));
 sky130_fd_sc_hd__nand2b_1 _23194_ (.A_N(_03458_),
    .B(_03453_),
    .Y(_03495_));
 sky130_fd_sc_hd__nor2b_1 _23195_ (.A(_03453_),
    .B_N(_03458_),
    .Y(_03496_));
 sky130_fd_sc_hd__a21oi_2 _23196_ (.A1(_03354_),
    .A2(_03495_),
    .B1(_03496_),
    .Y(_03497_));
 sky130_fd_sc_hd__o2111ai_4 _23197_ (.A1(_03242_),
    .A2(_03245_),
    .B1(_03342_),
    .C1(_03459_),
    .D1(_03185_),
    .Y(_03498_));
 sky130_fd_sc_hd__nand2_1 _23198_ (.A(_03497_),
    .B(_03498_),
    .Y(_03499_));
 sky130_fd_sc_hd__inv_1 _23199_ (.A(_03448_),
    .Y(_03500_));
 sky130_fd_sc_hd__inv_1 _23200_ (.A(_03451_),
    .Y(_03501_));
 sky130_fd_sc_hd__maj3_1 _23201_ (.A(_03500_),
    .B(_03501_),
    .C(_03444_),
    .X(_03502_));
 sky130_fd_sc_hd__maj3_1 _23202_ (.A(_03420_),
    .B(_03439_),
    .C(_03442_),
    .X(_03503_));
 sky130_fd_sc_hd__nor2b_1 _23203_ (.A(_03264_),
    .B_N(_03282_),
    .Y(_03504_));
 sky130_fd_sc_hd__nor2_1 _23204_ (.A(_03504_),
    .B(_03437_),
    .Y(_03505_));
 sky130_fd_sc_hd__nand2_1 _23205_ (.A(_03504_),
    .B(_03437_),
    .Y(_03506_));
 sky130_fd_sc_hd__o21ai_1 _23206_ (.A1(_03421_),
    .A2(_03505_),
    .B1(_03506_),
    .Y(_03507_));
 sky130_fd_sc_hd__nand2_4 _23207_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ),
    .Y(_03508_));
 sky130_fd_sc_hd__nor3_4 _23208_ (.A(_08294_),
    .B(_13439_),
    .C(_03423_),
    .Y(_03509_));
 sky130_fd_sc_hd__nand2_1 _23209_ (.A(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[49] ),
    .B(_03509_),
    .Y(_03510_));
 sky130_fd_sc_hd__nand2_2 _23210_ (.A(_03508_),
    .B(_03510_),
    .Y(_03511_));
 sky130_fd_sc_hd__nand4_4 _23211_ (.A(net316),
    .B(_10691_),
    .C(_13357_),
    .D(_01720_),
    .Y(_03512_));
 sky130_fd_sc_hd__xnor2_1 _23212_ (.A(_08950_),
    .B(net699),
    .Y(_03513_));
 sky130_fd_sc_hd__xnor2_1 _23213_ (.A(_09784_),
    .B(_09856_),
    .Y(_03514_));
 sky130_fd_sc_hd__mux2i_4 _23214_ (.A0(_03513_),
    .A1(_03514_),
    .S(net322),
    .Y(_03515_));
 sky130_fd_sc_hd__nor2_8 _23215_ (.A(_03512_),
    .B(_03515_),
    .Y(_03516_));
 sky130_fd_sc_hd__xnor2_4 _23216_ (.A(_03511_),
    .B(_03516_),
    .Y(_03517_));
 sky130_fd_sc_hd__maj3_2 _23217_ (.A(_03410_),
    .B(_03411_),
    .C(_03412_),
    .X(_03518_));
 sky130_fd_sc_hd__nor2_1 _23218_ (.A(net904),
    .B(_03425_),
    .Y(_03519_));
 sky130_fd_sc_hd__nand2_1 _23219_ (.A(_03425_),
    .B(_03426_),
    .Y(_03520_));
 sky130_fd_sc_hd__o21ai_2 _23220_ (.A1(_03429_),
    .A2(_03519_),
    .B1(_03520_),
    .Y(_03521_));
 sky130_fd_sc_hd__xor2_2 _23221_ (.A(_03518_),
    .B(_03521_),
    .X(_03522_));
 sky130_fd_sc_hd__xnor2_4 _23222_ (.A(_03517_),
    .B(_03522_),
    .Y(_03523_));
 sky130_fd_sc_hd__inv_1 _23223_ (.A(_03432_),
    .Y(_03524_));
 sky130_fd_sc_hd__maj3_2 _23224_ (.A(_03431_),
    .B(_03524_),
    .C(_03433_),
    .X(_03525_));
 sky130_fd_sc_hd__xor2_4 _23225_ (.A(_03523_),
    .B(_03525_),
    .X(_03526_));
 sky130_fd_sc_hd__maj3_1 _23226_ (.A(_03404_),
    .B(_03415_),
    .C(_03416_),
    .X(_03527_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_309 ();
 sky130_fd_sc_hd__o21a_1 _23228_ (.A1(_03376_),
    .A2(_03434_),
    .B1(_03435_),
    .X(_03529_));
 sky130_fd_sc_hd__a21oi_4 _23229_ (.A1(_03376_),
    .A2(_03434_),
    .B1(_03529_),
    .Y(_03530_));
 sky130_fd_sc_hd__xnor2_1 _23230_ (.A(_03527_),
    .B(_03530_),
    .Y(_03531_));
 sky130_fd_sc_hd__xnor2_1 _23231_ (.A(_03526_),
    .B(_03531_),
    .Y(_03532_));
 sky130_fd_sc_hd__a211oi_1 _23232_ (.A1(_02160_),
    .A2(_03161_),
    .B1(_03373_),
    .C1(_02158_),
    .Y(_03533_));
 sky130_fd_sc_hd__nor4_1 _23233_ (.A(net781),
    .B(net939),
    .C(_03313_),
    .D(_03370_),
    .Y(_03534_));
 sky130_fd_sc_hd__o21ai_0 _23234_ (.A1(_03533_),
    .A2(_03534_),
    .B1(net1287),
    .Y(_03535_));
 sky130_fd_sc_hd__o21ai_0 _23235_ (.A1(net939),
    .A2(_03313_),
    .B1(_03384_),
    .Y(_03536_));
 sky130_fd_sc_hd__o311ai_0 _23236_ (.A1(net939),
    .A2(_03313_),
    .A3(_03380_),
    .B1(_03536_),
    .C1(net781),
    .Y(_03537_));
 sky130_fd_sc_hd__nor2_1 _23237_ (.A(net939),
    .B(_03313_),
    .Y(_03538_));
 sky130_fd_sc_hd__nor2_1 _23238_ (.A(net781),
    .B(_03373_),
    .Y(_03539_));
 sky130_fd_sc_hd__o21ai_0 _23239_ (.A1(net1287),
    .A2(_03379_),
    .B1(_03310_),
    .Y(_03540_));
 sky130_fd_sc_hd__a21oi_1 _23240_ (.A1(_02160_),
    .A2(_03161_),
    .B1(net781),
    .Y(_03541_));
 sky130_fd_sc_hd__a32oi_1 _23241_ (.A1(_03379_),
    .A2(_03538_),
    .A3(_03539_),
    .B1(_03540_),
    .B2(_03541_),
    .Y(_03542_));
 sky130_fd_sc_hd__nand3_1 _23242_ (.A(_03535_),
    .B(_03537_),
    .C(_03542_),
    .Y(_03543_));
 sky130_fd_sc_hd__nor2_1 _23243_ (.A(_02080_),
    .B(_03165_),
    .Y(_03544_));
 sky130_fd_sc_hd__a21oi_1 _23244_ (.A1(net882),
    .A2(_02931_),
    .B1(_02150_),
    .Y(_03545_));
 sky130_fd_sc_hd__a211oi_2 _23245_ (.A1(net307),
    .A2(_01712_),
    .B1(net1069),
    .C1(net1222),
    .Y(_03546_));
 sky130_fd_sc_hd__xnor2_1 _23246_ (.A(_03545_),
    .B(_03546_),
    .Y(_03547_));
 sky130_fd_sc_hd__xnor2_1 _23247_ (.A(_03544_),
    .B(_03547_),
    .Y(_03548_));
 sky130_fd_sc_hd__nor2_1 _23248_ (.A(net792),
    .B(_03373_),
    .Y(_03549_));
 sky130_fd_sc_hd__nor2_1 _23249_ (.A(_01998_),
    .B(_03379_),
    .Y(_03550_));
 sky130_fd_sc_hd__maj3_1 _23250_ (.A(_03549_),
    .B(_03364_),
    .C(_03550_),
    .X(_03551_));
 sky130_fd_sc_hd__xnor2_1 _23251_ (.A(_03548_),
    .B(_03551_),
    .Y(_03552_));
 sky130_fd_sc_hd__xnor2_1 _23252_ (.A(_03543_),
    .B(_03552_),
    .Y(_03553_));
 sky130_fd_sc_hd__maj3_1 _23253_ (.A(_03360_),
    .B(_03361_),
    .C(_03362_),
    .X(_03554_));
 sky130_fd_sc_hd__nor2_1 _23254_ (.A(net1228),
    .B(_02730_),
    .Y(_03555_));
 sky130_fd_sc_hd__nor2_1 _23255_ (.A(_02513_),
    .B(_03142_),
    .Y(_03556_));
 sky130_fd_sc_hd__nor2_1 _23256_ (.A(net1277),
    .B(net1192),
    .Y(_03557_));
 sky130_fd_sc_hd__xnor3_1 _23257_ (.A(_03555_),
    .B(_03556_),
    .C(_03557_),
    .X(_03558_));
 sky130_fd_sc_hd__maj3_1 _23258_ (.A(_03394_),
    .B(_03395_),
    .C(_03396_),
    .X(_03559_));
 sky130_fd_sc_hd__xnor3_1 _23259_ (.A(_03554_),
    .B(_03558_),
    .C(_03559_),
    .X(_03560_));
 sky130_fd_sc_hd__nand3_1 _23260_ (.A(net1287),
    .B(_03310_),
    .C(_03384_),
    .Y(_03561_));
 sky130_fd_sc_hd__o21ai_0 _23261_ (.A1(net781),
    .A2(_03313_),
    .B1(net1178),
    .Y(_03562_));
 sky130_fd_sc_hd__o32a_1 _23262_ (.A1(_03549_),
    .A2(_03364_),
    .A3(_03550_),
    .B1(_03561_),
    .B2(_03562_),
    .X(_03563_));
 sky130_fd_sc_hd__o211ai_1 _23263_ (.A1(_03377_),
    .A2(_03380_),
    .B1(net1179),
    .C1(_03364_),
    .Y(_03564_));
 sky130_fd_sc_hd__nor3_1 _23264_ (.A(_02158_),
    .B(_03162_),
    .C(_03383_),
    .Y(_03565_));
 sky130_fd_sc_hd__a31oi_2 _23265_ (.A1(_03363_),
    .A2(_03563_),
    .A3(_03564_),
    .B1(_03565_),
    .Y(_03566_));
 sky130_fd_sc_hd__xnor2_1 _23266_ (.A(_03560_),
    .B(_03566_),
    .Y(_03567_));
 sky130_fd_sc_hd__xnor2_2 _23267_ (.A(_03567_),
    .B(_03553_),
    .Y(_03568_));
 sky130_fd_sc_hd__nand2_1 _23268_ (.A(_02301_),
    .B(_02889_),
    .Y(_03569_));
 sky130_fd_sc_hd__nand2_1 _23269_ (.A(_02421_),
    .B(_03407_),
    .Y(_03570_));
 sky130_fd_sc_hd__nand2_1 _23270_ (.A(net1181),
    .B(_02897_),
    .Y(_03571_));
 sky130_fd_sc_hd__xor3_1 _23271_ (.A(_03569_),
    .B(_03570_),
    .C(_03571_),
    .X(_03572_));
 sky130_fd_sc_hd__maj3_1 _23272_ (.A(_03405_),
    .B(_03406_),
    .C(_03408_),
    .X(_03573_));
 sky130_fd_sc_hd__a221oi_4 _23273_ (.A1(net305),
    .A2(net322),
    .B1(_03271_),
    .B2(_03273_),
    .C1(net302),
    .Y(_03574_));
 sky130_fd_sc_hd__a221oi_4 _23274_ (.A1(net1186),
    .A2(_01712_),
    .B1(_03039_),
    .B2(_03040_),
    .C1(_02061_),
    .Y(_03575_));
 sky130_fd_sc_hd__a2111oi_4 _23275_ (.A1(net303),
    .A2(net322),
    .B1(net1055),
    .C1(_03113_),
    .D1(net1063),
    .Y(_03576_));
 sky130_fd_sc_hd__xnor2_1 _23276_ (.A(_03575_),
    .B(_03576_),
    .Y(_03577_));
 sky130_fd_sc_hd__xor2_2 _23277_ (.A(_03574_),
    .B(_03577_),
    .X(_03578_));
 sky130_fd_sc_hd__xor2_1 _23278_ (.A(_03573_),
    .B(_03578_),
    .X(_03579_));
 sky130_fd_sc_hd__xnor2_2 _23279_ (.A(_03572_),
    .B(_03579_),
    .Y(_03580_));
 sky130_fd_sc_hd__maj3_1 _23280_ (.A(_03409_),
    .B(_03413_),
    .C(_03414_),
    .X(_03581_));
 sky130_fd_sc_hd__maj3_2 _23281_ (.A(_03393_),
    .B(_03397_),
    .C(_03398_),
    .X(_03582_));
 sky130_fd_sc_hd__xor2_1 _23282_ (.A(_03581_),
    .B(_03582_),
    .X(_03583_));
 sky130_fd_sc_hd__xnor2_2 _23283_ (.A(_03583_),
    .B(_03580_),
    .Y(_03584_));
 sky130_fd_sc_hd__inv_1 _23284_ (.A(_03390_),
    .Y(_03585_));
 sky130_fd_sc_hd__maj3_2 _23285_ (.A(_03585_),
    .B(_03389_),
    .C(_03399_),
    .X(_03586_));
 sky130_fd_sc_hd__xnor3_2 _23286_ (.A(_03586_),
    .B(_03584_),
    .C(_03568_),
    .X(_03587_));
 sky130_fd_sc_hd__maj3_2 _23287_ (.A(_03359_),
    .B(_03401_),
    .C(_03418_),
    .X(_03588_));
 sky130_fd_sc_hd__xor2_2 _23288_ (.A(_03588_),
    .B(_03587_),
    .X(_03589_));
 sky130_fd_sc_hd__xnor2_2 _23289_ (.A(_03589_),
    .B(_03532_),
    .Y(_03590_));
 sky130_fd_sc_hd__xor2_1 _23290_ (.A(_03590_),
    .B(_03507_),
    .X(_03591_));
 sky130_fd_sc_hd__xnor2_1 _23291_ (.A(_03591_),
    .B(_03503_),
    .Y(_03592_));
 sky130_fd_sc_hd__nand2_1 _23292_ (.A(_03592_),
    .B(_03502_),
    .Y(_03593_));
 sky130_fd_sc_hd__or2_4 _23293_ (.A(_03592_),
    .B(_03502_),
    .X(_03594_));
 sky130_fd_sc_hd__nand2_1 _23294_ (.A(_03593_),
    .B(_03594_),
    .Y(_03595_));
 sky130_fd_sc_hd__xnor2_4 _23295_ (.A(_03499_),
    .B(_03595_),
    .Y(_03596_));
 sky130_fd_sc_hd__nand2_1 _23296_ (.A(_02169_),
    .B(_03596_),
    .Y(_03597_));
 sky130_fd_sc_hd__o21ai_2 _23297_ (.A1(_02169_),
    .A2(_03494_),
    .B1(_03597_),
    .Y(_03598_));
 sky130_fd_sc_hd__mux2i_1 _23298_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[49] ),
    .A1(_03598_),
    .S(_08100_),
    .Y(_03599_));
 sky130_fd_sc_hd__nor2_1 _23299_ (.A(net295),
    .B(_03207_),
    .Y(_03600_));
 sky130_fd_sc_hd__a21oi_1 _23300_ (.A1(net295),
    .A2(_03204_),
    .B1(_03600_),
    .Y(_03601_));
 sky130_fd_sc_hd__nor2_1 _23301_ (.A(_09754_),
    .B(_01898_),
    .Y(_03602_));
 sky130_fd_sc_hd__nor2_1 _23302_ (.A(_09789_),
    .B(_01902_),
    .Y(_03603_));
 sky130_fd_sc_hd__a21oi_1 _23303_ (.A1(_09789_),
    .A2(_03602_),
    .B1(_03603_),
    .Y(_03604_));
 sky130_fd_sc_hd__nand2_1 _23304_ (.A(_09789_),
    .B(_02233_),
    .Y(_03605_));
 sky130_fd_sc_hd__nand2_1 _23305_ (.A(_09754_),
    .B(_03605_),
    .Y(_03606_));
 sky130_fd_sc_hd__o21ai_0 _23306_ (.A1(_01893_),
    .A2(_03604_),
    .B1(_03606_),
    .Y(_03607_));
 sky130_fd_sc_hd__o21ai_0 _23307_ (.A1(_01761_),
    .A2(_03601_),
    .B1(_03607_),
    .Y(_03608_));
 sky130_fd_sc_hd__a211oi_1 _23308_ (.A1(net158),
    .A2(_01929_),
    .B1(_03608_),
    .C1(net314),
    .Y(_03609_));
 sky130_fd_sc_hd__a21oi_1 _23309_ (.A1(net312),
    .A2(_03599_),
    .B1(_03609_),
    .Y(_03610_));
 sky130_fd_sc_hd__nor2_1 _23310_ (.A(_08632_),
    .B(_03610_),
    .Y(_03611_));
 sky130_fd_sc_hd__a21oi_2 _23311_ (.A1(_08632_),
    .A2(_11521_),
    .B1(_03611_),
    .Y(_03612_));
 sky130_fd_sc_hd__nor2_4 _23312_ (.A(_02646_),
    .B(_03612_),
    .Y(_03613_));
 sky130_fd_sc_hd__a31oi_4 _23313_ (.A1(_02646_),
    .A2(_03478_),
    .A3(_03486_),
    .B1(_03613_),
    .Y(_03614_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_308 ();
 sky130_fd_sc_hd__nand2_1 _23315_ (.A(_02119_),
    .B(_03614_),
    .Y(_03616_));
 sky130_fd_sc_hd__nand2_1 _23316_ (.A(\gen_regfile_ff.register_file_i.rf_reg[145] ),
    .B(_02123_),
    .Y(_03617_));
 sky130_fd_sc_hd__nand2_1 _23317_ (.A(_03616_),
    .B(_03617_),
    .Y(_00529_));
 sky130_fd_sc_hd__xor2_1 _23318_ (.A(_02020_),
    .B(_02025_),
    .X(_03618_));
 sky130_fd_sc_hd__xnor2_2 _23319_ (.A(_02041_),
    .B(_03618_),
    .Y(_03619_));
 sky130_fd_sc_hd__o21ai_0 _23320_ (.A1(_03358_),
    .A2(_03496_),
    .B1(_03495_),
    .Y(_03620_));
 sky130_fd_sc_hd__inv_1 _23321_ (.A(_03594_),
    .Y(_03621_));
 sky130_fd_sc_hd__a21oi_2 _23322_ (.A1(_03593_),
    .A2(_03620_),
    .B1(_03621_),
    .Y(_03622_));
 sky130_fd_sc_hd__nand2b_1 _23323_ (.A_N(_03503_),
    .B(_03590_),
    .Y(_03623_));
 sky130_fd_sc_hd__nor2b_1 _23324_ (.A(_03590_),
    .B_N(_03503_),
    .Y(_03624_));
 sky130_fd_sc_hd__a21o_1 _23325_ (.A1(_03507_),
    .A2(_03623_),
    .B1(_03624_),
    .X(_03625_));
 sky130_fd_sc_hd__nor2_1 _23326_ (.A(_03526_),
    .B(_03527_),
    .Y(_03626_));
 sky130_fd_sc_hd__inv_1 _23327_ (.A(_03587_),
    .Y(_03627_));
 sky130_fd_sc_hd__inv_1 _23328_ (.A(_03530_),
    .Y(_03628_));
 sky130_fd_sc_hd__and2_0 _23329_ (.A(_03628_),
    .B(_03588_),
    .X(_03629_));
 sky130_fd_sc_hd__or2_1 _23330_ (.A(_03628_),
    .B(_03588_),
    .X(_03630_));
 sky130_fd_sc_hd__o21ai_0 _23331_ (.A1(_03627_),
    .A2(_03629_),
    .B1(_03630_),
    .Y(_03631_));
 sky130_fd_sc_hd__nand2_1 _23332_ (.A(_03526_),
    .B(_03527_),
    .Y(_03632_));
 sky130_fd_sc_hd__o21a_1 _23333_ (.A1(_03587_),
    .A2(_03626_),
    .B1(_03632_),
    .X(_03633_));
 sky130_fd_sc_hd__or2_0 _23334_ (.A(_03587_),
    .B(_03632_),
    .X(_03634_));
 sky130_fd_sc_hd__o21ai_1 _23335_ (.A1(_03530_),
    .A2(_03633_),
    .B1(_03634_),
    .Y(_03635_));
 sky130_fd_sc_hd__nand2_1 _23336_ (.A(_03587_),
    .B(_03632_),
    .Y(_03636_));
 sky130_fd_sc_hd__o22ai_1 _23337_ (.A1(_03530_),
    .A2(_03634_),
    .B1(_03630_),
    .B2(_03636_),
    .Y(_03637_));
 sky130_fd_sc_hd__a221oi_2 _23338_ (.A1(_03626_),
    .A2(_03631_),
    .B1(_03635_),
    .B2(_03588_),
    .C1(_03637_),
    .Y(_03638_));
 sky130_fd_sc_hd__nor2_1 _23339_ (.A(_03548_),
    .B(_03551_),
    .Y(_03639_));
 sky130_fd_sc_hd__nand2_1 _23340_ (.A(_03548_),
    .B(_03551_),
    .Y(_03640_));
 sky130_fd_sc_hd__o21ai_2 _23341_ (.A1(_03543_),
    .A2(_03639_),
    .B1(_03640_),
    .Y(_03641_));
 sky130_fd_sc_hd__maj3_1 _23342_ (.A(_03380_),
    .B(_03538_),
    .C(_03539_),
    .X(_03642_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_307 ();
 sky130_fd_sc_hd__nor2_1 _23344_ (.A(_02150_),
    .B(net1243),
    .Y(_03644_));
 sky130_fd_sc_hd__a21oi_2 _23345_ (.A1(net882),
    .A2(_02931_),
    .B1(net1069),
    .Y(_03645_));
 sky130_fd_sc_hd__a211oi_4 _23346_ (.A1(net307),
    .A2(_01712_),
    .B1(net1228),
    .C1(net1222),
    .Y(_03646_));
 sky130_fd_sc_hd__xnor2_1 _23347_ (.A(_03645_),
    .B(_03646_),
    .Y(_03647_));
 sky130_fd_sc_hd__xnor2_1 _23348_ (.A(_03644_),
    .B(_03647_),
    .Y(_03648_));
 sky130_fd_sc_hd__nor2_1 _23349_ (.A(_02080_),
    .B(_03313_),
    .Y(_03649_));
 sky130_fd_sc_hd__nor2_1 _23350_ (.A(net939),
    .B(_03373_),
    .Y(_03650_));
 sky130_fd_sc_hd__nor2_1 _23351_ (.A(_02158_),
    .B(_03370_),
    .Y(_03651_));
 sky130_fd_sc_hd__xor3_1 _23352_ (.A(_03649_),
    .B(_03650_),
    .C(_03651_),
    .X(_03652_));
 sky130_fd_sc_hd__xor3_1 _23353_ (.A(_03642_),
    .B(_03648_),
    .C(_03652_),
    .X(_03653_));
 sky130_fd_sc_hd__maj3_1 _23354_ (.A(_03545_),
    .B(_03544_),
    .C(_03546_),
    .X(_03654_));
 sky130_fd_sc_hd__nor2_1 _23355_ (.A(net1161),
    .B(net1413),
    .Y(_03655_));
 sky130_fd_sc_hd__nor2_1 _23356_ (.A(_03142_),
    .B(net1173),
    .Y(_03656_));
 sky130_fd_sc_hd__nor2_1 _23357_ (.A(net1004),
    .B(_02730_),
    .Y(_03657_));
 sky130_fd_sc_hd__xor3_1 _23358_ (.A(_03655_),
    .B(_03656_),
    .C(_03657_),
    .X(_03658_));
 sky130_fd_sc_hd__maj3_1 _23359_ (.A(_03555_),
    .B(_03556_),
    .C(_03557_),
    .X(_03659_));
 sky130_fd_sc_hd__xnor3_1 _23360_ (.A(_03654_),
    .B(_03658_),
    .C(_03659_),
    .X(_03660_));
 sky130_fd_sc_hd__xnor2_1 _23361_ (.A(_03653_),
    .B(_03660_),
    .Y(_03661_));
 sky130_fd_sc_hd__xnor2_2 _23362_ (.A(_03641_),
    .B(_03661_),
    .Y(_03662_));
 sky130_fd_sc_hd__maj3_1 _23363_ (.A(_03569_),
    .B(_03570_),
    .C(_03571_),
    .X(_03663_));
 sky130_fd_sc_hd__nand2_1 _23364_ (.A(net898),
    .B(_02897_),
    .Y(_03664_));
 sky130_fd_sc_hd__nand2_1 _23365_ (.A(net1181),
    .B(_03041_),
    .Y(_03665_));
 sky130_fd_sc_hd__nand2_1 _23366_ (.A(_02421_),
    .B(_02889_),
    .Y(_03666_));
 sky130_fd_sc_hd__xor3_1 _23367_ (.A(_03664_),
    .B(_03665_),
    .C(_03666_),
    .X(_03667_));
 sky130_fd_sc_hd__a2111oi_4 _23368_ (.A1(net1186),
    .A2(_01712_),
    .B1(_02061_),
    .C1(_03113_),
    .D1(net1063),
    .Y(_03668_));
 sky130_fd_sc_hd__a221oi_4 _23369_ (.A1(net303),
    .A2(net322),
    .B1(_03271_),
    .B2(_03273_),
    .C1(net1054),
    .Y(_03669_));
 sky130_fd_sc_hd__nand4_4 _23370_ (.A(_10676_),
    .B(_10683_),
    .C(_10690_),
    .D(_03427_),
    .Y(_03670_));
 sky130_fd_sc_hd__a211oi_2 _23371_ (.A1(net305),
    .A2(net322),
    .B1(net302),
    .C1(_03670_),
    .Y(_03671_));
 sky130_fd_sc_hd__xnor2_1 _23372_ (.A(_03669_),
    .B(_03671_),
    .Y(_03672_));
 sky130_fd_sc_hd__xor2_2 _23373_ (.A(_03668_),
    .B(_03672_),
    .X(_03673_));
 sky130_fd_sc_hd__xor3_1 _23374_ (.A(_03663_),
    .B(_03667_),
    .C(_03673_),
    .X(_03674_));
 sky130_fd_sc_hd__maj3_2 _23375_ (.A(_03554_),
    .B(_03558_),
    .C(_03559_),
    .X(_03675_));
 sky130_fd_sc_hd__maj3_1 _23376_ (.A(_03572_),
    .B(_03573_),
    .C(_03578_),
    .X(_03676_));
 sky130_fd_sc_hd__xnor2_1 _23377_ (.A(_03675_),
    .B(_03676_),
    .Y(_03677_));
 sky130_fd_sc_hd__xnor2_1 _23378_ (.A(_03674_),
    .B(_03677_),
    .Y(_03678_));
 sky130_fd_sc_hd__inv_1 _23379_ (.A(_03560_),
    .Y(_03679_));
 sky130_fd_sc_hd__maj3_1 _23380_ (.A(_03679_),
    .B(_03553_),
    .C(_03566_),
    .X(_03680_));
 sky130_fd_sc_hd__xor2_1 _23381_ (.A(_03678_),
    .B(_03680_),
    .X(_03681_));
 sky130_fd_sc_hd__xnor2_2 _23382_ (.A(_03662_),
    .B(_03681_),
    .Y(_03682_));
 sky130_fd_sc_hd__maj3_2 _23383_ (.A(_03574_),
    .B(_03575_),
    .C(_03576_),
    .X(_03683_));
 sky130_fd_sc_hd__nor4b_4 _23384_ (.A(_13439_),
    .B(_13440_),
    .C(_03508_),
    .D_N(_13357_),
    .Y(_03684_));
 sky130_fd_sc_hd__a21oi_4 _23385_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[50] ),
    .A2(_03509_),
    .B1(_03684_),
    .Y(_03685_));
 sky130_fd_sc_hd__xnor2_2 _23386_ (.A(_03683_),
    .B(_03685_),
    .Y(_03686_));
 sky130_fd_sc_hd__nor2_1 _23387_ (.A(_03511_),
    .B(_03518_),
    .Y(_03687_));
 sky130_fd_sc_hd__nand2_2 _23388_ (.A(net316),
    .B(_13357_),
    .Y(_03688_));
 sky130_fd_sc_hd__nor3b_4 _23389_ (.A(_01968_),
    .B(_03688_),
    .C_N(_10691_),
    .Y(_03689_));
 sky130_fd_sc_hd__nand2b_4 _23390_ (.A_N(_03515_),
    .B(_03689_),
    .Y(_03690_));
 sky130_fd_sc_hd__and3_1 _23391_ (.A(_03511_),
    .B(_03690_),
    .C(_03518_),
    .X(_03691_));
 sky130_fd_sc_hd__and2_1 _23392_ (.A(_03508_),
    .B(_03510_),
    .X(_03692_));
 sky130_fd_sc_hd__xnor2_1 _23393_ (.A(_03692_),
    .B(_03516_),
    .Y(_03693_));
 sky130_fd_sc_hd__o32ai_1 _23394_ (.A1(_03521_),
    .A2(_03687_),
    .A3(_03691_),
    .B1(_03518_),
    .B2(_03693_),
    .Y(_03694_));
 sky130_fd_sc_hd__nand3_4 _23395_ (.A(_02032_),
    .B(net905),
    .C(_03689_),
    .Y(_03695_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_305 ();
 sky130_fd_sc_hd__nor3_4 _23398_ (.A(net947),
    .B(net857),
    .C(_03512_),
    .Y(_03698_));
 sky130_fd_sc_hd__nand3_1 _23399_ (.A(_03511_),
    .B(_03690_),
    .C(_03698_),
    .Y(_03699_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_304 ();
 sky130_fd_sc_hd__nand2_1 _23401_ (.A(_03692_),
    .B(_03516_),
    .Y(_03701_));
 sky130_fd_sc_hd__nor2_1 _23402_ (.A(_03518_),
    .B(_03521_),
    .Y(_03702_));
 sky130_fd_sc_hd__a21oi_1 _23403_ (.A1(_03699_),
    .A2(_03701_),
    .B1(_03702_),
    .Y(_03703_));
 sky130_fd_sc_hd__nand2_1 _23404_ (.A(_03518_),
    .B(_03521_),
    .Y(_03704_));
 sky130_fd_sc_hd__nor2_1 _23405_ (.A(_03704_),
    .B(_03695_),
    .Y(_03705_));
 sky130_fd_sc_hd__a211oi_2 _23406_ (.A1(_03694_),
    .A2(_03695_),
    .B1(_03703_),
    .C1(_03705_),
    .Y(_03706_));
 sky130_fd_sc_hd__xnor2_2 _23407_ (.A(_03686_),
    .B(_03706_),
    .Y(_03707_));
 sky130_fd_sc_hd__nand2_1 _23408_ (.A(_03523_),
    .B(_03525_),
    .Y(_03708_));
 sky130_fd_sc_hd__inv_1 _23409_ (.A(_03582_),
    .Y(_03709_));
 sky130_fd_sc_hd__maj3_1 _23410_ (.A(_03580_),
    .B(_03581_),
    .C(_03709_),
    .X(_03710_));
 sky130_fd_sc_hd__xnor2_1 _23411_ (.A(_03708_),
    .B(_03710_),
    .Y(_03711_));
 sky130_fd_sc_hd__xnor2_2 _23412_ (.A(_03707_),
    .B(_03711_),
    .Y(_03712_));
 sky130_fd_sc_hd__o21a_1 _23413_ (.A1(_03568_),
    .A2(net1511),
    .B1(_03586_),
    .X(_03713_));
 sky130_fd_sc_hd__a21oi_2 _23414_ (.A1(_03568_),
    .A2(_03584_),
    .B1(_03713_),
    .Y(_03714_));
 sky130_fd_sc_hd__xnor2_2 _23415_ (.A(_03712_),
    .B(_03714_),
    .Y(_03715_));
 sky130_fd_sc_hd__xnor2_4 _23416_ (.A(_03682_),
    .B(_03715_),
    .Y(_03716_));
 sky130_fd_sc_hd__xnor2_1 _23417_ (.A(_03716_),
    .B(_03638_),
    .Y(_03717_));
 sky130_fd_sc_hd__nand2_1 _23418_ (.A(_03625_),
    .B(_03717_),
    .Y(_03718_));
 sky130_fd_sc_hd__or2_4 _23419_ (.A(_03625_),
    .B(_03717_),
    .X(_03719_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_303 ();
 sky130_fd_sc_hd__nand2_1 _23421_ (.A(_03718_),
    .B(_03719_),
    .Y(_03721_));
 sky130_fd_sc_hd__xor2_4 _23422_ (.A(_03622_),
    .B(_03721_),
    .X(_03722_));
 sky130_fd_sc_hd__nand2_1 _23423_ (.A(_02169_),
    .B(_03722_),
    .Y(_03723_));
 sky130_fd_sc_hd__nand2_8 _23424_ (.A(net443),
    .B(net312),
    .Y(_03724_));
 sky130_fd_sc_hd__o211ai_4 _23425_ (.A1(_02169_),
    .A2(_03619_),
    .B1(_03723_),
    .C1(_03724_),
    .Y(_03725_));
 sky130_fd_sc_hd__a21oi_1 _23426_ (.A1(net443),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[50] ),
    .B1(net739),
    .Y(_03726_));
 sky130_fd_sc_hd__nand3_1 _23427_ (.A(_09898_),
    .B(_09932_),
    .C(_02228_),
    .Y(_03727_));
 sky130_fd_sc_hd__o21ai_0 _23428_ (.A1(_09932_),
    .A2(_01902_),
    .B1(_03727_),
    .Y(_03728_));
 sky130_fd_sc_hd__a21oi_1 _23429_ (.A1(_09932_),
    .A2(_02233_),
    .B1(_09898_),
    .Y(_03729_));
 sky130_fd_sc_hd__a21oi_1 _23430_ (.A1(_02225_),
    .A2(_03728_),
    .B1(_03729_),
    .Y(_03730_));
 sky130_fd_sc_hd__nor2_1 _23431_ (.A(net295),
    .B(_02987_),
    .Y(_03731_));
 sky130_fd_sc_hd__a211oi_2 _23432_ (.A1(net295),
    .A2(_02985_),
    .B1(_03731_),
    .C1(_01761_),
    .Y(_03732_));
 sky130_fd_sc_hd__a2111oi_0 _23433_ (.A1(net159),
    .A2(_01929_),
    .B1(_03730_),
    .C1(_03732_),
    .D1(net312),
    .Y(_03733_));
 sky130_fd_sc_hd__a21oi_1 _23434_ (.A1(_03725_),
    .A2(_03726_),
    .B1(_03733_),
    .Y(_03734_));
 sky130_fd_sc_hd__nand2_1 _23435_ (.A(_08632_),
    .B(_11543_),
    .Y(_03735_));
 sky130_fd_sc_hd__o21ai_4 _23436_ (.A1(_03734_),
    .A2(_08632_),
    .B1(_03735_),
    .Y(_03736_));
 sky130_fd_sc_hd__mux4_1 _23437_ (.A0(net36),
    .A1(net49),
    .A2(\load_store_unit_i.rdata_q[26] ),
    .A3(net28),
    .S0(\load_store_unit_i.rdata_offset_q[1] ),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .X(_03737_));
 sky130_fd_sc_hd__a21oi_1 _23438_ (.A1(_01674_),
    .A2(_03737_),
    .B1(_03479_),
    .Y(_03738_));
 sky130_fd_sc_hd__a21oi_4 _23439_ (.A1(_03736_),
    .A2(net266),
    .B1(_03738_),
    .Y(_03739_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_302 ();
 sky130_fd_sc_hd__nand2_1 _23441_ (.A(_02119_),
    .B(_03739_),
    .Y(_03741_));
 sky130_fd_sc_hd__nand2_1 _23442_ (.A(\gen_regfile_ff.register_file_i.rf_reg[146] ),
    .B(_02123_),
    .Y(_03742_));
 sky130_fd_sc_hd__nand2_1 _23443_ (.A(_03741_),
    .B(_03742_),
    .Y(_00530_));
 sky130_fd_sc_hd__mux4_1 _23444_ (.A0(net37),
    .A1(net52),
    .A2(\load_store_unit_i.rdata_q[27] ),
    .A3(net29),
    .S0(\load_store_unit_i.rdata_offset_q[1] ),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .X(_03743_));
 sky130_fd_sc_hd__nand2_1 _23445_ (.A(_01674_),
    .B(_03743_),
    .Y(_03744_));
 sky130_fd_sc_hd__nand2_1 _23446_ (.A(_08632_),
    .B(_11560_),
    .Y(_03745_));
 sky130_fd_sc_hd__nand2b_1 _23447_ (.A_N(_02020_),
    .B(_02025_),
    .Y(_03746_));
 sky130_fd_sc_hd__nand2b_1 _23448_ (.A_N(_02038_),
    .B(_02049_),
    .Y(_03747_));
 sky130_fd_sc_hd__a21oi_1 _23449_ (.A1(_03746_),
    .A2(_03747_),
    .B1(_02036_),
    .Y(_03748_));
 sky130_fd_sc_hd__o22ai_1 _23450_ (.A1(_02040_),
    .A2(_02049_),
    .B1(_03746_),
    .B2(_02038_),
    .Y(_03749_));
 sky130_fd_sc_hd__nor2_1 _23451_ (.A(_03748_),
    .B(_03749_),
    .Y(_03750_));
 sky130_fd_sc_hd__xnor2_2 _23452_ (.A(_02013_),
    .B(_03750_),
    .Y(_03751_));
 sky130_fd_sc_hd__nand2_1 _23453_ (.A(_01698_),
    .B(_03751_),
    .Y(_03752_));
 sky130_fd_sc_hd__and2_4 _23454_ (.A(_03593_),
    .B(_03718_),
    .X(_03753_));
 sky130_fd_sc_hd__a32oi_4 _23455_ (.A1(_03753_),
    .A2(_03497_),
    .A3(_03498_),
    .B1(_03718_),
    .B2(_03621_),
    .Y(_03754_));
 sky130_fd_sc_hd__nand2_1 _23456_ (.A(_03708_),
    .B(_03707_),
    .Y(_03755_));
 sky130_fd_sc_hd__nor2_1 _23457_ (.A(_03708_),
    .B(_03707_),
    .Y(_03756_));
 sky130_fd_sc_hd__a21oi_2 _23458_ (.A1(_03710_),
    .A2(_03755_),
    .B1(_03756_),
    .Y(_03757_));
 sky130_fd_sc_hd__inv_1 _23459_ (.A(_03682_),
    .Y(_03758_));
 sky130_fd_sc_hd__inv_1 _23460_ (.A(_03712_),
    .Y(_03759_));
 sky130_fd_sc_hd__maj3_1 _23461_ (.A(_03758_),
    .B(_03759_),
    .C(_03714_),
    .X(_03760_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_301 ();
 sky130_fd_sc_hd__o21ai_0 _23463_ (.A1(_03668_),
    .A2(_03669_),
    .B1(_02024_),
    .Y(_03762_));
 sky130_fd_sc_hd__maj3_1 _23464_ (.A(_02024_),
    .B(_03668_),
    .C(_03669_),
    .X(_03763_));
 sky130_fd_sc_hd__maj3_1 _23465_ (.A(_09784_),
    .B(net1190),
    .C(_03685_),
    .X(_03764_));
 sky130_fd_sc_hd__nand4_2 _23466_ (.A(_08967_),
    .B(_08978_),
    .C(_08986_),
    .D(_08994_),
    .Y(_03765_));
 sky130_fd_sc_hd__maj3_1 _23467_ (.A(_08950_),
    .B(_03765_),
    .C(_03685_),
    .X(_03766_));
 sky130_fd_sc_hd__mux2_1 _23468_ (.A0(_03764_),
    .A1(_03766_),
    .S(net320),
    .X(_03767_));
 sky130_fd_sc_hd__mux2i_1 _23469_ (.A0(_03762_),
    .A1(_03763_),
    .S(_03767_),
    .Y(_03768_));
 sky130_fd_sc_hd__nand2_1 _23470_ (.A(_03668_),
    .B(_03669_),
    .Y(_03769_));
 sky130_fd_sc_hd__a21oi_1 _23471_ (.A1(_03689_),
    .A2(_03767_),
    .B1(_03769_),
    .Y(_03770_));
 sky130_fd_sc_hd__a21oi_2 _23472_ (.A1(_03689_),
    .A2(_03768_),
    .B1(_03770_),
    .Y(_03771_));
 sky130_fd_sc_hd__nor2_8 _23473_ (.A(_13442_),
    .B(_03508_),
    .Y(_03772_));
 sky130_fd_sc_hd__a21oi_4 _23474_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[51] ),
    .A2(_03424_),
    .B1(_03772_),
    .Y(_03773_));
 sky130_fd_sc_hd__xnor2_2 _23475_ (.A(_03771_),
    .B(_03773_),
    .Y(_03774_));
 sky130_fd_sc_hd__o21ai_0 _23476_ (.A1(_03575_),
    .A2(_03576_),
    .B1(_03574_),
    .Y(_03775_));
 sky130_fd_sc_hd__a21boi_2 _23477_ (.A1(_03575_),
    .A2(_03576_),
    .B1_N(_03775_),
    .Y(_03776_));
 sky130_fd_sc_hd__xnor2_1 _23478_ (.A(_03690_),
    .B(_03685_),
    .Y(_03777_));
 sky130_fd_sc_hd__nor2_4 _23479_ (.A(_03688_),
    .B(_03508_),
    .Y(_03778_));
 sky130_fd_sc_hd__a21o_1 _23480_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[50] ),
    .A2(_08292_),
    .B1(_03778_),
    .X(_03779_));
 sky130_fd_sc_hd__nand2_1 _23481_ (.A(_03683_),
    .B(_03779_),
    .Y(_03780_));
 sky130_fd_sc_hd__o31ai_1 _23482_ (.A1(_03512_),
    .A2(_03515_),
    .A3(_03685_),
    .B1(_03683_),
    .Y(_03781_));
 sky130_fd_sc_hd__a22o_1 _23483_ (.A1(_03690_),
    .A2(_03780_),
    .B1(_03781_),
    .B2(_03692_),
    .X(_03782_));
 sky130_fd_sc_hd__a22oi_1 _23484_ (.A1(_03776_),
    .A2(_03777_),
    .B1(_03782_),
    .B2(_03695_),
    .Y(_03783_));
 sky130_fd_sc_hd__xnor2_1 _23485_ (.A(_03774_),
    .B(_03783_),
    .Y(_03784_));
 sky130_fd_sc_hd__maj3_1 _23486_ (.A(_03675_),
    .B(_03674_),
    .C(_03676_),
    .X(_03785_));
 sky130_fd_sc_hd__o31ai_1 _23487_ (.A1(_03512_),
    .A2(_03511_),
    .A3(_03515_),
    .B1(_03695_),
    .Y(_03786_));
 sky130_fd_sc_hd__xnor2_1 _23488_ (.A(_03686_),
    .B(_03786_),
    .Y(_03787_));
 sky130_fd_sc_hd__a211oi_2 _23489_ (.A1(_03517_),
    .A2(_03704_),
    .B1(_03787_),
    .C1(_03702_),
    .Y(_03788_));
 sky130_fd_sc_hd__xnor2_1 _23490_ (.A(_03785_),
    .B(_03788_),
    .Y(_03789_));
 sky130_fd_sc_hd__xnor2_1 _23491_ (.A(_03784_),
    .B(_03789_),
    .Y(_03790_));
 sky130_fd_sc_hd__maj3_1 _23492_ (.A(_03662_),
    .B(_03678_),
    .C(_03680_),
    .X(_03791_));
 sky130_fd_sc_hd__nor2_1 _23493_ (.A(_03790_),
    .B(_03791_),
    .Y(_03792_));
 sky130_fd_sc_hd__and2_0 _23494_ (.A(_03790_),
    .B(_03791_),
    .X(_03793_));
 sky130_fd_sc_hd__nor2_1 _23495_ (.A(_03792_),
    .B(_03793_),
    .Y(_03794_));
 sky130_fd_sc_hd__nor2_1 _23496_ (.A(net1228),
    .B(_02932_),
    .Y(_03795_));
 sky130_fd_sc_hd__nor2_1 _23497_ (.A(net1069),
    .B(net1243),
    .Y(_03796_));
 sky130_fd_sc_hd__nand2_1 _23498_ (.A(_03004_),
    .B(_02774_),
    .Y(_03797_));
 sky130_fd_sc_hd__xnor3_1 _23499_ (.A(_03795_),
    .B(_03796_),
    .C(_03797_),
    .X(_03798_));
 sky130_fd_sc_hd__nand2_1 _23500_ (.A(_02436_),
    .B(_03161_),
    .Y(_03799_));
 sky130_fd_sc_hd__o211ai_2 _23501_ (.A1(_09707_),
    .A2(net322),
    .B1(_02440_),
    .C1(_03309_),
    .Y(_03800_));
 sky130_fd_sc_hd__nand3_2 _23502_ (.A(_02083_),
    .B(_02085_),
    .C(_03384_),
    .Y(_03801_));
 sky130_fd_sc_hd__xor2_1 _23503_ (.A(_03800_),
    .B(_03801_),
    .X(_03802_));
 sky130_fd_sc_hd__xnor2_1 _23504_ (.A(_03799_),
    .B(_03802_),
    .Y(_03803_));
 sky130_fd_sc_hd__maj3_1 _23505_ (.A(_03649_),
    .B(_03650_),
    .C(_03651_),
    .X(_03804_));
 sky130_fd_sc_hd__xor3_1 _23506_ (.A(_03798_),
    .B(_03803_),
    .C(_03804_),
    .X(_03805_));
 sky130_fd_sc_hd__maj3_1 _23507_ (.A(_03642_),
    .B(_03648_),
    .C(_03652_),
    .X(_03806_));
 sky130_fd_sc_hd__maj3_1 _23508_ (.A(_03645_),
    .B(_03644_),
    .C(_03646_),
    .X(_03807_));
 sky130_fd_sc_hd__nand2b_1 _23509_ (.A_N(_02513_),
    .B(_02889_),
    .Y(_03808_));
 sky130_fd_sc_hd__nand2_1 _23510_ (.A(_02589_),
    .B(_02727_),
    .Y(_03809_));
 sky130_fd_sc_hd__nand2b_1 _23511_ (.A_N(net1192),
    .B(_03407_),
    .Y(_03810_));
 sky130_fd_sc_hd__xor3_1 _23512_ (.A(_03808_),
    .B(_03809_),
    .C(_03810_),
    .X(_03811_));
 sky130_fd_sc_hd__maj3_1 _23513_ (.A(_03655_),
    .B(_03656_),
    .C(_03657_),
    .X(_03812_));
 sky130_fd_sc_hd__xnor3_1 _23514_ (.A(_03807_),
    .B(_03811_),
    .C(_03812_),
    .X(_03813_));
 sky130_fd_sc_hd__xor2_1 _23515_ (.A(_03806_),
    .B(_03813_),
    .X(_03814_));
 sky130_fd_sc_hd__xnor2_2 _23516_ (.A(_03805_),
    .B(_03814_),
    .Y(_03815_));
 sky130_fd_sc_hd__nor2b_1 _23517_ (.A(_03660_),
    .B_N(_03653_),
    .Y(_03816_));
 sky130_fd_sc_hd__nand2b_1 _23518_ (.A_N(_03653_),
    .B(_03660_),
    .Y(_03817_));
 sky130_fd_sc_hd__o21ai_2 _23519_ (.A1(_03641_),
    .A2(_03816_),
    .B1(_03817_),
    .Y(_03818_));
 sky130_fd_sc_hd__maj3_1 _23520_ (.A(_03664_),
    .B(_03665_),
    .C(_03666_),
    .X(_03819_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_300 ();
 sky130_fd_sc_hd__nor2_1 _23522_ (.A(net909),
    .B(_03119_),
    .Y(_03821_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_299 ();
 sky130_fd_sc_hd__nor2_1 _23524_ (.A(net1216),
    .B(_03097_),
    .Y(_03823_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_298 ();
 sky130_fd_sc_hd__nor2_1 _23526_ (.A(_02289_),
    .B(_03100_),
    .Y(_03825_));
 sky130_fd_sc_hd__xnor2_1 _23527_ (.A(_03823_),
    .B(_03825_),
    .Y(_03826_));
 sky130_fd_sc_hd__xnor2_1 _23528_ (.A(_03821_),
    .B(_03826_),
    .Y(_03827_));
 sky130_fd_sc_hd__a221oi_4 _23529_ (.A1(net1186),
    .A2(_01712_),
    .B1(_03271_),
    .B2(_03273_),
    .C1(_02061_),
    .Y(_03828_));
 sky130_fd_sc_hd__nor2_1 _23530_ (.A(_02010_),
    .B(_02005_),
    .Y(_03829_));
 sky130_fd_sc_hd__nor2_1 _23531_ (.A(_02024_),
    .B(_02088_),
    .Y(_03830_));
 sky130_fd_sc_hd__o21ai_1 _23532_ (.A1(_03829_),
    .A2(_03830_),
    .B1(_03689_),
    .Y(_03831_));
 sky130_fd_sc_hd__xnor2_2 _23533_ (.A(_03828_),
    .B(_03831_),
    .Y(_03832_));
 sky130_fd_sc_hd__xnor3_1 _23534_ (.A(_03819_),
    .B(_03827_),
    .C(_03832_),
    .X(_03833_));
 sky130_fd_sc_hd__maj3_1 _23535_ (.A(_03654_),
    .B(_03658_),
    .C(_03659_),
    .X(_03834_));
 sky130_fd_sc_hd__maj3_1 _23536_ (.A(_03663_),
    .B(_03667_),
    .C(_03673_),
    .X(_03835_));
 sky130_fd_sc_hd__xnor2_1 _23537_ (.A(_03834_),
    .B(_03835_),
    .Y(_03836_));
 sky130_fd_sc_hd__xnor2_1 _23538_ (.A(_03833_),
    .B(_03836_),
    .Y(_03837_));
 sky130_fd_sc_hd__xnor2_1 _23539_ (.A(_03818_),
    .B(_03837_),
    .Y(_03838_));
 sky130_fd_sc_hd__xnor2_1 _23540_ (.A(_03815_),
    .B(_03838_),
    .Y(_03839_));
 sky130_fd_sc_hd__xnor2_1 _23541_ (.A(_03794_),
    .B(_03839_),
    .Y(_03840_));
 sky130_fd_sc_hd__xnor2_1 _23542_ (.A(_03760_),
    .B(_03840_),
    .Y(_03841_));
 sky130_fd_sc_hd__xnor2_2 _23543_ (.A(_03757_),
    .B(_03841_),
    .Y(_03842_));
 sky130_fd_sc_hd__o21bai_1 _23544_ (.A1(_03633_),
    .A2(_03716_),
    .B1_N(_03629_),
    .Y(_03843_));
 sky130_fd_sc_hd__nand2_1 _23545_ (.A(_03633_),
    .B(_03716_),
    .Y(_03844_));
 sky130_fd_sc_hd__nand2_1 _23546_ (.A(_03627_),
    .B(_03630_),
    .Y(_03845_));
 sky130_fd_sc_hd__a21oi_1 _23547_ (.A1(_03632_),
    .A2(_03716_),
    .B1(_03845_),
    .Y(_03846_));
 sky130_fd_sc_hd__nor3b_1 _23548_ (.A(_03716_),
    .B(_03626_),
    .C_N(_03630_),
    .Y(_03847_));
 sky130_fd_sc_hd__a211o_4 _23549_ (.A1(_03843_),
    .A2(_03844_),
    .B1(_03846_),
    .C1(_03847_),
    .X(_03848_));
 sky130_fd_sc_hd__xor2_1 _23550_ (.A(_03842_),
    .B(_03848_),
    .X(_03849_));
 sky130_fd_sc_hd__a21oi_1 _23551_ (.A1(_03719_),
    .A2(_03754_),
    .B1(_03849_),
    .Y(_03850_));
 sky130_fd_sc_hd__and3_1 _23552_ (.A(_03719_),
    .B(_03754_),
    .C(_03849_),
    .X(_03851_));
 sky130_fd_sc_hd__o21ai_1 _23553_ (.A1(_03850_),
    .A2(_03851_),
    .B1(_02169_),
    .Y(_03852_));
 sky130_fd_sc_hd__nand2_1 _23554_ (.A(_03752_),
    .B(_03852_),
    .Y(_03853_));
 sky130_fd_sc_hd__nor2_1 _23555_ (.A(net441),
    .B(_03853_),
    .Y(_03854_));
 sky130_fd_sc_hd__a211oi_4 _23556_ (.A1(net441),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[51] ),
    .B1(net739),
    .C1(_03854_),
    .Y(_03855_));
 sky130_fd_sc_hd__nor2_1 _23557_ (.A(net295),
    .B(_02864_),
    .Y(_03856_));
 sky130_fd_sc_hd__a21oi_1 _23558_ (.A1(net295),
    .A2(_02870_),
    .B1(_03856_),
    .Y(_03857_));
 sky130_fd_sc_hd__nor2_1 _23559_ (.A(_10001_),
    .B(_01902_),
    .Y(_03858_));
 sky130_fd_sc_hd__a31oi_1 _23560_ (.A1(_10001_),
    .A2(_10008_),
    .A3(_02228_),
    .B1(_03858_),
    .Y(_03859_));
 sky130_fd_sc_hd__a21o_1 _23561_ (.A1(_10001_),
    .A2(_02233_),
    .B1(_10008_),
    .X(_03860_));
 sky130_fd_sc_hd__o21ai_0 _23562_ (.A1(_01893_),
    .A2(_03859_),
    .B1(_03860_),
    .Y(_03861_));
 sky130_fd_sc_hd__o21ai_0 _23563_ (.A1(_01761_),
    .A2(_03857_),
    .B1(_03861_),
    .Y(_03862_));
 sky130_fd_sc_hd__a211oi_1 _23564_ (.A1(net160),
    .A2(_01929_),
    .B1(_03862_),
    .C1(net314),
    .Y(_03863_));
 sky130_fd_sc_hd__o21ai_1 _23565_ (.A1(_03855_),
    .A2(_03863_),
    .B1(_08581_),
    .Y(_03864_));
 sky130_fd_sc_hd__a21oi_4 _23566_ (.A1(_03864_),
    .A2(_03745_),
    .B1(_02646_),
    .Y(_03865_));
 sky130_fd_sc_hd__a31oi_4 _23567_ (.A1(_02646_),
    .A2(_03478_),
    .A3(_03744_),
    .B1(net1553),
    .Y(_03866_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_297 ();
 sky130_fd_sc_hd__nand2_1 _23569_ (.A(_02119_),
    .B(_03866_),
    .Y(_03868_));
 sky130_fd_sc_hd__nand2_1 _23570_ (.A(\gen_regfile_ff.register_file_i.rf_reg[147] ),
    .B(_02123_),
    .Y(_03869_));
 sky130_fd_sc_hd__nand2_1 _23571_ (.A(_03868_),
    .B(_03869_),
    .Y(_00531_));
 sky130_fd_sc_hd__mux4_1 _23572_ (.A0(net39),
    .A1(net53),
    .A2(\load_store_unit_i.rdata_q[28] ),
    .A3(net30),
    .S0(\load_store_unit_i.rdata_offset_q[1] ),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .X(_03870_));
 sky130_fd_sc_hd__nand2_1 _23573_ (.A(_01674_),
    .B(_03870_),
    .Y(_03871_));
 sky130_fd_sc_hd__nor2b_1 _23574_ (.A(_03757_),
    .B_N(_03840_),
    .Y(_03872_));
 sky130_fd_sc_hd__nor2b_1 _23575_ (.A(_03840_),
    .B_N(_03757_),
    .Y(_03873_));
 sky130_fd_sc_hd__nor2_1 _23576_ (.A(_03760_),
    .B(_03873_),
    .Y(_03874_));
 sky130_fd_sc_hd__nor2_1 _23577_ (.A(_03793_),
    .B(_03839_),
    .Y(_03875_));
 sky130_fd_sc_hd__nor2_1 _23578_ (.A(_03792_),
    .B(_03875_),
    .Y(_03876_));
 sky130_fd_sc_hd__inv_1 _23579_ (.A(_03785_),
    .Y(_03877_));
 sky130_fd_sc_hd__maj3_1 _23580_ (.A(_03877_),
    .B(_03788_),
    .C(_03784_),
    .X(_03878_));
 sky130_fd_sc_hd__maj3_1 _23581_ (.A(_03815_),
    .B(_03818_),
    .C(_03837_),
    .X(_03879_));
 sky130_fd_sc_hd__nand2_1 _23582_ (.A(_03807_),
    .B(_03812_),
    .Y(_03880_));
 sky130_fd_sc_hd__nor2_1 _23583_ (.A(_03807_),
    .B(_03812_),
    .Y(_03881_));
 sky130_fd_sc_hd__a21oi_2 _23584_ (.A1(_03811_),
    .A2(_03880_),
    .B1(_03881_),
    .Y(_03882_));
 sky130_fd_sc_hd__nor3_1 _23585_ (.A(_02010_),
    .B(_02005_),
    .C(_03828_),
    .Y(_03883_));
 sky130_fd_sc_hd__and3_1 _23586_ (.A(_02024_),
    .B(_02005_),
    .C(_03828_),
    .X(_03884_));
 sky130_fd_sc_hd__nor3_2 _23587_ (.A(_02024_),
    .B(_02088_),
    .C(_02286_),
    .Y(_03885_));
 sky130_fd_sc_hd__nor3_1 _23588_ (.A(_02024_),
    .B(_02005_),
    .C(_02292_),
    .Y(_03886_));
 sky130_fd_sc_hd__or4_4 _23589_ (.A(_03883_),
    .B(_03884_),
    .C(_03885_),
    .D(_03886_),
    .X(_03887_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_296 ();
 sky130_fd_sc_hd__nand2_1 _23591_ (.A(_03689_),
    .B(_03887_),
    .Y(_03889_));
 sky130_fd_sc_hd__nand2_1 _23592_ (.A(net1181),
    .B(_03274_),
    .Y(_03890_));
 sky130_fd_sc_hd__nand2_1 _23593_ (.A(_02421_),
    .B(_03041_),
    .Y(_03891_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_295 ();
 sky130_fd_sc_hd__nand2_1 _23595_ (.A(net898),
    .B(_03265_),
    .Y(_03893_));
 sky130_fd_sc_hd__xnor3_1 _23596_ (.A(_03890_),
    .B(_03891_),
    .C(_03893_),
    .X(_03894_));
 sky130_fd_sc_hd__maj3_1 _23597_ (.A(_03823_),
    .B(_03821_),
    .C(_03825_),
    .X(_03895_));
 sky130_fd_sc_hd__xnor2_1 _23598_ (.A(_03894_),
    .B(_03895_),
    .Y(_03896_));
 sky130_fd_sc_hd__xnor2_1 _23599_ (.A(_03889_),
    .B(_03896_),
    .Y(_03897_));
 sky130_fd_sc_hd__inv_1 _23600_ (.A(_03819_),
    .Y(_03898_));
 sky130_fd_sc_hd__maj3_1 _23601_ (.A(_03898_),
    .B(_03827_),
    .C(_03832_),
    .X(_03899_));
 sky130_fd_sc_hd__xnor3_1 _23602_ (.A(_03882_),
    .B(_03897_),
    .C(_03899_),
    .X(_03900_));
 sky130_fd_sc_hd__nor2_1 _23603_ (.A(net1277),
    .B(_02932_),
    .Y(_03901_));
 sky130_fd_sc_hd__nor2_1 _23604_ (.A(net1228),
    .B(net1243),
    .Y(_03902_));
 sky130_fd_sc_hd__nor2_1 _23605_ (.A(_03142_),
    .B(_02936_),
    .Y(_03903_));
 sky130_fd_sc_hd__xnor3_1 _23606_ (.A(_03901_),
    .B(_03902_),
    .C(_03903_),
    .X(_03904_));
 sky130_fd_sc_hd__nand2b_1 _23607_ (.A_N(net1069),
    .B(_03161_),
    .Y(_03905_));
 sky130_fd_sc_hd__nand2_1 _23608_ (.A(_02436_),
    .B(_03310_),
    .Y(_03906_));
 sky130_fd_sc_hd__nand2_1 _23609_ (.A(_02080_),
    .B(_03376_),
    .Y(_03907_));
 sky130_fd_sc_hd__xor3_4 _23610_ (.A(_03905_),
    .B(_03906_),
    .C(_03907_),
    .X(_03908_));
 sky130_fd_sc_hd__maj3_1 _23611_ (.A(_03799_),
    .B(_03800_),
    .C(_03801_),
    .X(_03909_));
 sky130_fd_sc_hd__xnor3_1 _23612_ (.A(_03904_),
    .B(_03908_),
    .C(_03909_),
    .X(_03910_));
 sky130_fd_sc_hd__maj3_1 _23613_ (.A(_03798_),
    .B(_03803_),
    .C(_03804_),
    .X(_03911_));
 sky130_fd_sc_hd__o22ai_1 _23614_ (.A1(net1004),
    .A2(_02936_),
    .B1(_02932_),
    .B2(net1228),
    .Y(_03912_));
 sky130_fd_sc_hd__nor4_1 _23615_ (.A(net1228),
    .B(net1004),
    .C(_02936_),
    .D(net899),
    .Y(_03913_));
 sky130_fd_sc_hd__a21oi_1 _23616_ (.A1(_03796_),
    .A2(_03912_),
    .B1(_03913_),
    .Y(_03914_));
 sky130_fd_sc_hd__nor2_1 _23617_ (.A(net1192),
    .B(net1239),
    .Y(_03915_));
 sky130_fd_sc_hd__nor2_1 _23618_ (.A(_02730_),
    .B(net1413),
    .Y(_03916_));
 sky130_fd_sc_hd__nor2_1 _23619_ (.A(net1161),
    .B(_03097_),
    .Y(_03917_));
 sky130_fd_sc_hd__xnor3_1 _23620_ (.A(_03915_),
    .B(_03916_),
    .C(_03917_),
    .X(_03918_));
 sky130_fd_sc_hd__maj3_1 _23621_ (.A(_03808_),
    .B(_03809_),
    .C(_03810_),
    .X(_03919_));
 sky130_fd_sc_hd__xor3_1 _23622_ (.A(_03914_),
    .B(_03918_),
    .C(_03919_),
    .X(_03920_));
 sky130_fd_sc_hd__xnor3_1 _23623_ (.A(_03910_),
    .B(_03911_),
    .C(_03920_),
    .X(_03921_));
 sky130_fd_sc_hd__maj3_1 _23624_ (.A(_03805_),
    .B(_03806_),
    .C(_03813_),
    .X(_03922_));
 sky130_fd_sc_hd__xor2_1 _23625_ (.A(_03921_),
    .B(_03922_),
    .X(_03923_));
 sky130_fd_sc_hd__xnor2_2 _23626_ (.A(_03900_),
    .B(_03923_),
    .Y(_03924_));
 sky130_fd_sc_hd__inv_1 _23627_ (.A(_03835_),
    .Y(_03925_));
 sky130_fd_sc_hd__maj3_2 _23628_ (.A(_03834_),
    .B(_03833_),
    .C(_03925_),
    .X(_03926_));
 sky130_fd_sc_hd__nor2_8 _23629_ (.A(_03670_),
    .B(_03515_),
    .Y(_03927_));
 sky130_fd_sc_hd__a21oi_2 _23630_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[50] ),
    .A2(_03424_),
    .B1(_03772_),
    .Y(_03928_));
 sky130_fd_sc_hd__nor2_1 _23631_ (.A(_03776_),
    .B(_03928_),
    .Y(_03929_));
 sky130_fd_sc_hd__nand2_1 _23632_ (.A(_03692_),
    .B(_03781_),
    .Y(_03930_));
 sky130_fd_sc_hd__o21ai_0 _23633_ (.A1(_03927_),
    .A2(_03929_),
    .B1(_03930_),
    .Y(_03931_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_294 ();
 sky130_fd_sc_hd__nand3_4 _23635_ (.A(_02032_),
    .B(net904),
    .C(_03428_),
    .Y(_03933_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_293 ();
 sky130_fd_sc_hd__a221oi_2 _23637_ (.A1(_03776_),
    .A2(_03777_),
    .B1(_03931_),
    .B2(_03933_),
    .C1(_03774_),
    .Y(_03935_));
 sky130_fd_sc_hd__maj3_4 _23638_ (.A(_02024_),
    .B(_02005_),
    .C(_03828_),
    .X(_03936_));
 sky130_fd_sc_hd__and2_4 _23639_ (.A(_03428_),
    .B(_03936_),
    .X(_03937_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_292 ();
 sky130_fd_sc_hd__a21oi_4 _23641_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[52] ),
    .A2(_03424_),
    .B1(_03772_),
    .Y(_03939_));
 sky130_fd_sc_hd__xnor2_2 _23642_ (.A(_03937_),
    .B(_03939_),
    .Y(_03940_));
 sky130_fd_sc_hd__nor2_8 _23643_ (.A(net857),
    .B(_03429_),
    .Y(_03941_));
 sky130_fd_sc_hd__a21o_1 _23644_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[51] ),
    .A2(_03424_),
    .B1(_03772_),
    .X(_03942_));
 sky130_fd_sc_hd__nor3_1 _23645_ (.A(_03928_),
    .B(_03941_),
    .C(_03942_),
    .Y(_03943_));
 sky130_fd_sc_hd__maj3_4 _23646_ (.A(_03668_),
    .B(_03669_),
    .C(_03671_),
    .X(_03944_));
 sky130_fd_sc_hd__nor2_1 _23647_ (.A(_03773_),
    .B(_03944_),
    .Y(_03945_));
 sky130_fd_sc_hd__and3_1 _23648_ (.A(_03927_),
    .B(_03928_),
    .C(_03944_),
    .X(_03946_));
 sky130_fd_sc_hd__nand2_1 _23649_ (.A(_03941_),
    .B(_03944_),
    .Y(_03947_));
 sky130_fd_sc_hd__nand2_1 _23650_ (.A(_03933_),
    .B(_03773_),
    .Y(_03948_));
 sky130_fd_sc_hd__a21oi_1 _23651_ (.A1(_03947_),
    .A2(_03948_),
    .B1(_03927_),
    .Y(_03949_));
 sky130_fd_sc_hd__nor4_1 _23652_ (.A(_03943_),
    .B(_03945_),
    .C(_03946_),
    .D(_03949_),
    .Y(_03950_));
 sky130_fd_sc_hd__xnor2_2 _23653_ (.A(_03940_),
    .B(_03950_),
    .Y(_03951_));
 sky130_fd_sc_hd__xor2_1 _23654_ (.A(_03935_),
    .B(_03951_),
    .X(_03952_));
 sky130_fd_sc_hd__xnor2_1 _23655_ (.A(_03926_),
    .B(_03952_),
    .Y(_03953_));
 sky130_fd_sc_hd__xnor2_1 _23656_ (.A(_03924_),
    .B(_03953_),
    .Y(_03954_));
 sky130_fd_sc_hd__xnor2_1 _23657_ (.A(_03879_),
    .B(_03954_),
    .Y(_03955_));
 sky130_fd_sc_hd__xor2_1 _23658_ (.A(_03878_),
    .B(_03955_),
    .X(_03956_));
 sky130_fd_sc_hd__xnor2_1 _23659_ (.A(_03876_),
    .B(_03956_),
    .Y(_03957_));
 sky130_fd_sc_hd__o21ai_2 _23660_ (.A1(_03872_),
    .A2(_03874_),
    .B1(_03957_),
    .Y(_03958_));
 sky130_fd_sc_hd__or3_2 _23661_ (.A(_03872_),
    .B(_03874_),
    .C(_03957_),
    .X(_03959_));
 sky130_fd_sc_hd__nand2_1 _23662_ (.A(_03958_),
    .B(_03959_),
    .Y(_03960_));
 sky130_fd_sc_hd__nor2b_4 _23663_ (.A(_03458_),
    .B_N(_03453_),
    .Y(_03961_));
 sky130_fd_sc_hd__a311oi_2 _23664_ (.A1(_03187_),
    .A2(_03190_),
    .A3(_03355_),
    .B1(_03357_),
    .C1(_03961_),
    .Y(_03962_));
 sky130_fd_sc_hd__o21ai_2 _23665_ (.A1(_03496_),
    .A2(_03962_),
    .B1(_03594_),
    .Y(_03963_));
 sky130_fd_sc_hd__a21boi_4 _23666_ (.A1(_03753_),
    .A2(net1522),
    .B1_N(_03719_),
    .Y(_03964_));
 sky130_fd_sc_hd__maj3_2 _23667_ (.A(_03842_),
    .B(_03964_),
    .C(_03848_),
    .X(_03965_));
 sky130_fd_sc_hd__xnor2_2 _23668_ (.A(_03960_),
    .B(_03965_),
    .Y(_03966_));
 sky130_fd_sc_hd__nand2_2 _23669_ (.A(_02169_),
    .B(_03966_),
    .Y(_03967_));
 sky130_fd_sc_hd__o21ai_4 _23670_ (.A1(_02169_),
    .A2(_02097_),
    .B1(_03967_),
    .Y(_03968_));
 sky130_fd_sc_hd__mux2i_4 _23671_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[52] ),
    .A1(_03968_),
    .S(_08100_),
    .Y(_03969_));
 sky130_fd_sc_hd__nor2_1 _23672_ (.A(_01773_),
    .B(_02838_),
    .Y(_03970_));
 sky130_fd_sc_hd__a21oi_1 _23673_ (.A1(_01773_),
    .A2(_02832_),
    .B1(_03970_),
    .Y(_03971_));
 sky130_fd_sc_hd__nor2_1 _23674_ (.A(_10044_),
    .B(_01898_),
    .Y(_03972_));
 sky130_fd_sc_hd__nor2_1 _23675_ (.A(_10070_),
    .B(_01902_),
    .Y(_03973_));
 sky130_fd_sc_hd__a21oi_1 _23676_ (.A1(_10070_),
    .A2(_03972_),
    .B1(_03973_),
    .Y(_03974_));
 sky130_fd_sc_hd__nand2_1 _23677_ (.A(_10070_),
    .B(_02233_),
    .Y(_03975_));
 sky130_fd_sc_hd__nand2_1 _23678_ (.A(_10044_),
    .B(_03975_),
    .Y(_03976_));
 sky130_fd_sc_hd__o21ai_0 _23679_ (.A1(_01893_),
    .A2(_03974_),
    .B1(_03976_),
    .Y(_03977_));
 sky130_fd_sc_hd__o21ai_0 _23680_ (.A1(_01761_),
    .A2(_03971_),
    .B1(_03977_),
    .Y(_03978_));
 sky130_fd_sc_hd__a211oi_1 _23681_ (.A1(net1007),
    .A2(_01929_),
    .B1(_03978_),
    .C1(net314),
    .Y(_03979_));
 sky130_fd_sc_hd__a21oi_4 _23682_ (.A1(_03969_),
    .A2(net314),
    .B1(_03979_),
    .Y(_03980_));
 sky130_fd_sc_hd__nor3_4 _23683_ (.A(_03980_),
    .B(_02646_),
    .C(_11597_),
    .Y(_03981_));
 sky130_fd_sc_hd__a31oi_4 _23684_ (.A1(_02646_),
    .A2(_03478_),
    .A3(_03871_),
    .B1(_03981_),
    .Y(_03982_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_291 ();
 sky130_fd_sc_hd__nand2_1 _23686_ (.A(_02119_),
    .B(_03982_),
    .Y(_03984_));
 sky130_fd_sc_hd__nand2_1 _23687_ (.A(\gen_regfile_ff.register_file_i.rf_reg[148] ),
    .B(_02123_),
    .Y(_03985_));
 sky130_fd_sc_hd__nand2_1 _23688_ (.A(_03984_),
    .B(_03985_),
    .Y(_00532_));
 sky130_fd_sc_hd__mux4_1 _23689_ (.A0(net40),
    .A1(net54),
    .A2(\load_store_unit_i.rdata_q[29] ),
    .A3(net31),
    .S0(\load_store_unit_i.rdata_offset_q[1] ),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .X(_03986_));
 sky130_fd_sc_hd__nand2_1 _23690_ (.A(_01674_),
    .B(_03986_),
    .Y(_03987_));
 sky130_fd_sc_hd__maj3_1 _23691_ (.A(_03719_),
    .B(_03842_),
    .C(_03848_),
    .X(_03988_));
 sky130_fd_sc_hd__nand2_1 _23692_ (.A(_03959_),
    .B(_03988_),
    .Y(_03989_));
 sky130_fd_sc_hd__nand2_1 _23693_ (.A(_03842_),
    .B(_03848_),
    .Y(_03990_));
 sky130_fd_sc_hd__a21boi_0 _23694_ (.A1(_03990_),
    .A2(_03958_),
    .B1_N(_03959_),
    .Y(_03991_));
 sky130_fd_sc_hd__o2bb2a_4 _23695_ (.A1_N(_03958_),
    .A2_N(_03989_),
    .B1(_03991_),
    .B2(_03754_),
    .X(_03992_));
 sky130_fd_sc_hd__nand2_1 _23696_ (.A(_02150_),
    .B(_03376_),
    .Y(_03993_));
 sky130_fd_sc_hd__nand2_1 _23697_ (.A(_02918_),
    .B(_03161_),
    .Y(_03994_));
 sky130_fd_sc_hd__nand2b_1 _23698_ (.A_N(net1069),
    .B(_03310_),
    .Y(_03995_));
 sky130_fd_sc_hd__xor2_1 _23699_ (.A(_03994_),
    .B(_03995_),
    .X(_03996_));
 sky130_fd_sc_hd__xor2_2 _23700_ (.A(_03993_),
    .B(_03996_),
    .X(_03997_));
 sky130_fd_sc_hd__nor2_1 _23701_ (.A(_03142_),
    .B(_02932_),
    .Y(_03998_));
 sky130_fd_sc_hd__nor2_1 _23702_ (.A(net1413),
    .B(_02936_),
    .Y(_03999_));
 sky130_fd_sc_hd__nor2_1 _23703_ (.A(net1004),
    .B(net1243),
    .Y(_04000_));
 sky130_fd_sc_hd__xnor3_1 _23704_ (.A(_03998_),
    .B(_03999_),
    .C(_04000_),
    .X(_04001_));
 sky130_fd_sc_hd__maj3_1 _23705_ (.A(_03905_),
    .B(_03906_),
    .C(_03907_),
    .X(_04002_));
 sky130_fd_sc_hd__xnor2_1 _23706_ (.A(_04001_),
    .B(_04002_),
    .Y(_04003_));
 sky130_fd_sc_hd__xnor2_2 _23707_ (.A(_03997_),
    .B(_04003_),
    .Y(_04004_));
 sky130_fd_sc_hd__nor2_1 _23708_ (.A(net1161),
    .B(_03100_),
    .Y(_04005_));
 sky130_fd_sc_hd__a221oi_4 _23709_ (.A1(_02619_),
    .A2(_01712_),
    .B1(_02895_),
    .B2(_02896_),
    .C1(net855),
    .Y(_04006_));
 sky130_fd_sc_hd__nor3_1 _23710_ (.A(_02723_),
    .B(_02725_),
    .C(net1239),
    .Y(_04007_));
 sky130_fd_sc_hd__xnor2_1 _23711_ (.A(_04006_),
    .B(_04007_),
    .Y(_04008_));
 sky130_fd_sc_hd__xnor2_2 _23712_ (.A(_04005_),
    .B(_04008_),
    .Y(_04009_));
 sky130_fd_sc_hd__maj3_1 _23713_ (.A(_03901_),
    .B(_03902_),
    .C(_03903_),
    .X(_04010_));
 sky130_fd_sc_hd__maj3_1 _23714_ (.A(_03915_),
    .B(_03916_),
    .C(_03917_),
    .X(_04011_));
 sky130_fd_sc_hd__xnor2_1 _23715_ (.A(_04010_),
    .B(_04011_),
    .Y(_04012_));
 sky130_fd_sc_hd__xor2_1 _23716_ (.A(_04009_),
    .B(_04012_),
    .X(_04013_));
 sky130_fd_sc_hd__maj3_1 _23717_ (.A(_03904_),
    .B(_03908_),
    .C(_03909_),
    .X(_04014_));
 sky130_fd_sc_hd__xor3_1 _23718_ (.A(_04004_),
    .B(_04013_),
    .C(_04014_),
    .X(_04015_));
 sky130_fd_sc_hd__xnor2_1 _23719_ (.A(_03904_),
    .B(_03909_),
    .Y(_04016_));
 sky130_fd_sc_hd__xnor2_1 _23720_ (.A(_03908_),
    .B(_04016_),
    .Y(_04017_));
 sky130_fd_sc_hd__inv_1 _23721_ (.A(_03911_),
    .Y(_04018_));
 sky130_fd_sc_hd__maj3_1 _23722_ (.A(_04017_),
    .B(_04018_),
    .C(_03920_),
    .X(_04019_));
 sky130_fd_sc_hd__and2_4 _23723_ (.A(_03271_),
    .B(_03273_),
    .X(_04020_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_290 ();
 sky130_fd_sc_hd__nand2_1 _23725_ (.A(net898),
    .B(_04020_),
    .Y(_04022_));
 sky130_fd_sc_hd__nor2_1 _23726_ (.A(_03119_),
    .B(_04020_),
    .Y(_04023_));
 sky130_fd_sc_hd__nor4_1 _23727_ (.A(net910),
    .B(_02289_),
    .C(net1010),
    .D(_03265_),
    .Y(_04024_));
 sky130_fd_sc_hd__a31oi_1 _23728_ (.A1(net1167),
    .A2(_02289_),
    .A3(_04023_),
    .B1(_04024_),
    .Y(_04025_));
 sky130_fd_sc_hd__a21oi_1 _23729_ (.A1(_04022_),
    .A2(_04025_),
    .B1(_03100_),
    .Y(_04026_));
 sky130_fd_sc_hd__nor2_1 _23730_ (.A(_02289_),
    .B(net1216),
    .Y(_04027_));
 sky130_fd_sc_hd__a32oi_1 _23731_ (.A1(_03100_),
    .A2(_04023_),
    .A3(_04027_),
    .B1(_03119_),
    .B2(_02289_),
    .Y(_04028_));
 sky130_fd_sc_hd__nor2_1 _23732_ (.A(net1168),
    .B(_04028_),
    .Y(_04029_));
 sky130_fd_sc_hd__a21oi_1 _23733_ (.A1(_03100_),
    .A2(_03119_),
    .B1(net1010),
    .Y(_04030_));
 sky130_fd_sc_hd__o21ai_0 _23734_ (.A1(_04020_),
    .A2(_03821_),
    .B1(net1010),
    .Y(_04031_));
 sky130_fd_sc_hd__o221ai_1 _23735_ (.A1(_03265_),
    .A2(_03274_),
    .B1(_04030_),
    .B2(net898),
    .C1(_04031_),
    .Y(_04032_));
 sky130_fd_sc_hd__nor3_1 _23736_ (.A(_04026_),
    .B(_04029_),
    .C(_04032_),
    .Y(_04033_));
 sky130_fd_sc_hd__xnor2_1 _23737_ (.A(net1168),
    .B(_03887_),
    .Y(_04034_));
 sky130_fd_sc_hd__nor2_2 _23738_ (.A(_03512_),
    .B(_04034_),
    .Y(_04035_));
 sky130_fd_sc_hd__maj3_1 _23739_ (.A(_03914_),
    .B(_03918_),
    .C(_03919_),
    .X(_04036_));
 sky130_fd_sc_hd__o41a_1 _23740_ (.A1(_03883_),
    .A2(_03884_),
    .A3(_03885_),
    .A4(_03886_),
    .B1(_03428_),
    .X(_04037_));
 sky130_fd_sc_hd__maj3_1 _23741_ (.A(_03894_),
    .B(_03895_),
    .C(_04037_),
    .X(_04038_));
 sky130_fd_sc_hd__xnor2_1 _23742_ (.A(_04036_),
    .B(_04038_),
    .Y(_04039_));
 sky130_fd_sc_hd__xnor3_1 _23743_ (.A(_04033_),
    .B(_04035_),
    .C(_04039_),
    .X(_04040_));
 sky130_fd_sc_hd__xnor3_2 _23744_ (.A(_04015_),
    .B(_04019_),
    .C(_04040_),
    .X(_04041_));
 sky130_fd_sc_hd__inv_1 _23745_ (.A(_03897_),
    .Y(_04042_));
 sky130_fd_sc_hd__maj3_1 _23746_ (.A(_03882_),
    .B(_04042_),
    .C(_03899_),
    .X(_04043_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_288 ();
 sky130_fd_sc_hd__a21oi_4 _23749_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[53] ),
    .A2(_03424_),
    .B1(_03772_),
    .Y(_04046_));
 sky130_fd_sc_hd__a21oi_1 _23750_ (.A1(_03933_),
    .A2(_03939_),
    .B1(_03937_),
    .Y(_04047_));
 sky130_fd_sc_hd__o22ai_2 _23751_ (.A1(_03933_),
    .A2(_03939_),
    .B1(_04047_),
    .B2(_03942_),
    .Y(_04048_));
 sky130_fd_sc_hd__nand2_8 _23752_ (.A(_03428_),
    .B(_03936_),
    .Y(_04049_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_287 ();
 sky130_fd_sc_hd__o21ai_0 _23754_ (.A1(_03670_),
    .A2(_03515_),
    .B1(_03939_),
    .Y(_04051_));
 sky130_fd_sc_hd__a21oi_1 _23755_ (.A1(_04049_),
    .A2(_04051_),
    .B1(_03933_),
    .Y(_04052_));
 sky130_fd_sc_hd__a221oi_4 _23756_ (.A1(_03937_),
    .A2(_03939_),
    .B1(_04048_),
    .B2(_03927_),
    .C1(_04052_),
    .Y(_04053_));
 sky130_fd_sc_hd__xor2_4 _23757_ (.A(_04046_),
    .B(_04053_),
    .X(_04054_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_285 ();
 sky130_fd_sc_hd__nand2_1 _23760_ (.A(_03773_),
    .B(_03944_),
    .Y(_04057_));
 sky130_fd_sc_hd__nor4_1 _23761_ (.A(_03670_),
    .B(_03515_),
    .C(_03942_),
    .D(_03940_),
    .Y(_04058_));
 sky130_fd_sc_hd__a31oi_1 _23762_ (.A1(_03942_),
    .A2(_03940_),
    .A3(_03944_),
    .B1(_04058_),
    .Y(_04059_));
 sky130_fd_sc_hd__a31oi_1 _23763_ (.A1(_03927_),
    .A2(_03928_),
    .A3(_04057_),
    .B1(_04059_),
    .Y(_04060_));
 sky130_fd_sc_hd__and2_4 _23764_ (.A(_03689_),
    .B(_03936_),
    .X(_04061_));
 sky130_fd_sc_hd__a21oi_1 _23765_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[52] ),
    .A2(_03509_),
    .B1(_03684_),
    .Y(_04062_));
 sky130_fd_sc_hd__xnor2_1 _23766_ (.A(_04061_),
    .B(_04062_),
    .Y(_04063_));
 sky130_fd_sc_hd__a21oi_1 _23767_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[51] ),
    .A2(_03509_),
    .B1(_03684_),
    .Y(_04064_));
 sky130_fd_sc_hd__or2_0 _23768_ (.A(_04064_),
    .B(_03944_),
    .X(_04065_));
 sky130_fd_sc_hd__nor2_1 _23769_ (.A(_03942_),
    .B(_03944_),
    .Y(_04066_));
 sky130_fd_sc_hd__nor3_1 _23770_ (.A(_03516_),
    .B(_03940_),
    .C(_04066_),
    .Y(_04067_));
 sky130_fd_sc_hd__a31oi_1 _23771_ (.A1(_03516_),
    .A2(_04063_),
    .A3(_04065_),
    .B1(_04067_),
    .Y(_04068_));
 sky130_fd_sc_hd__nor2_1 _23772_ (.A(_03933_),
    .B(_04068_),
    .Y(_04069_));
 sky130_fd_sc_hd__a21oi_1 _23773_ (.A1(_03933_),
    .A2(_04060_),
    .B1(_04069_),
    .Y(_04070_));
 sky130_fd_sc_hd__xnor3_1 _23774_ (.A(_04043_),
    .B(_04054_),
    .C(_04070_),
    .X(_04071_));
 sky130_fd_sc_hd__maj3_1 _23775_ (.A(_03921_),
    .B(_03900_),
    .C(_03922_),
    .X(_04072_));
 sky130_fd_sc_hd__xnor2_1 _23776_ (.A(_04071_),
    .B(_04072_),
    .Y(_04073_));
 sky130_fd_sc_hd__xnor2_2 _23777_ (.A(_04041_),
    .B(_04073_),
    .Y(_04074_));
 sky130_fd_sc_hd__inv_1 _23778_ (.A(_03935_),
    .Y(_04075_));
 sky130_fd_sc_hd__and2_1 _23779_ (.A(_03879_),
    .B(_03924_),
    .X(_04076_));
 sky130_fd_sc_hd__nor2_1 _23780_ (.A(_03879_),
    .B(_03924_),
    .Y(_04077_));
 sky130_fd_sc_hd__nor2_1 _23781_ (.A(_03926_),
    .B(_04077_),
    .Y(_04078_));
 sky130_fd_sc_hd__nand2_1 _23782_ (.A(_03926_),
    .B(_04077_),
    .Y(_04079_));
 sky130_fd_sc_hd__o31a_1 _23783_ (.A1(_03951_),
    .A2(_04076_),
    .A3(_04078_),
    .B1(_04079_),
    .X(_04080_));
 sky130_fd_sc_hd__nor2b_1 _23784_ (.A(_03774_),
    .B_N(_03783_),
    .Y(_04081_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_284 ();
 sky130_fd_sc_hd__nand2_1 _23786_ (.A(_03698_),
    .B(_03944_),
    .Y(_04083_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_283 ();
 sky130_fd_sc_hd__nand2_1 _23788_ (.A(_03695_),
    .B(_04064_),
    .Y(_04085_));
 sky130_fd_sc_hd__a21oi_1 _23789_ (.A1(_04083_),
    .A2(_04085_),
    .B1(_03516_),
    .Y(_04086_));
 sky130_fd_sc_hd__o21ai_0 _23790_ (.A1(_03685_),
    .A2(_04085_),
    .B1(_04065_),
    .Y(_04087_));
 sky130_fd_sc_hd__a311oi_1 _23791_ (.A1(_03516_),
    .A2(_03685_),
    .A3(_03944_),
    .B1(_04086_),
    .C1(_04087_),
    .Y(_04088_));
 sky130_fd_sc_hd__xor2_1 _23792_ (.A(_04063_),
    .B(_04088_),
    .X(_04089_));
 sky130_fd_sc_hd__inv_1 _23793_ (.A(_04076_),
    .Y(_04090_));
 sky130_fd_sc_hd__a211o_1 _23794_ (.A1(_04081_),
    .A2(_04089_),
    .B1(_04090_),
    .C1(_03926_),
    .X(_04091_));
 sky130_fd_sc_hd__o211ai_1 _23795_ (.A1(_04076_),
    .A2(_04078_),
    .B1(_04075_),
    .C1(_03951_),
    .Y(_04092_));
 sky130_fd_sc_hd__o211a_1 _23796_ (.A1(_03951_),
    .A2(_04079_),
    .B1(_04091_),
    .C1(_04092_),
    .X(_04093_));
 sky130_fd_sc_hd__o21ai_1 _23797_ (.A1(_04075_),
    .A2(_04080_),
    .B1(_04093_),
    .Y(_04094_));
 sky130_fd_sc_hd__xnor2_1 _23798_ (.A(_04074_),
    .B(_04094_),
    .Y(_04095_));
 sky130_fd_sc_hd__nor2_1 _23799_ (.A(_03878_),
    .B(_03955_),
    .Y(_04096_));
 sky130_fd_sc_hd__nand2_1 _23800_ (.A(_03878_),
    .B(_03955_),
    .Y(_04097_));
 sky130_fd_sc_hd__o21ai_0 _23801_ (.A1(_03876_),
    .A2(_04096_),
    .B1(_04097_),
    .Y(_04098_));
 sky130_fd_sc_hd__or2_1 _23802_ (.A(_04095_),
    .B(_04098_),
    .X(_04099_));
 sky130_fd_sc_hd__inv_1 _23803_ (.A(_04099_),
    .Y(_04100_));
 sky130_fd_sc_hd__and2_1 _23804_ (.A(_04095_),
    .B(_04098_),
    .X(_04101_));
 sky130_fd_sc_hd__nor2_1 _23805_ (.A(_04100_),
    .B(_04101_),
    .Y(_04102_));
 sky130_fd_sc_hd__xnor2_1 _23806_ (.A(_03992_),
    .B(_04102_),
    .Y(_04103_));
 sky130_fd_sc_hd__nor2_1 _23807_ (.A(_02169_),
    .B(_02168_),
    .Y(_04104_));
 sky130_fd_sc_hd__a21oi_2 _23808_ (.A1(_02169_),
    .A2(_04103_),
    .B1(_04104_),
    .Y(_04105_));
 sky130_fd_sc_hd__mux2i_1 _23809_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[53] ),
    .A1(_04105_),
    .S(_08100_),
    .Y(_04106_));
 sky130_fd_sc_hd__nand2_2 _23810_ (.A(net312),
    .B(_04106_),
    .Y(_04107_));
 sky130_fd_sc_hd__nand2_1 _23811_ (.A(net295),
    .B(_02662_),
    .Y(_04108_));
 sky130_fd_sc_hd__o21ai_2 _23812_ (.A1(net295),
    .A2(_02659_),
    .B1(_04108_),
    .Y(_04109_));
 sky130_fd_sc_hd__nand3_1 _23813_ (.A(_10112_),
    .B(_10145_),
    .C(_02228_),
    .Y(_04110_));
 sky130_fd_sc_hd__o21ai_0 _23814_ (.A1(_10145_),
    .A2(_01902_),
    .B1(_04110_),
    .Y(_04111_));
 sky130_fd_sc_hd__a21oi_1 _23815_ (.A1(_10145_),
    .A2(_02233_),
    .B1(_10112_),
    .Y(_04112_));
 sky130_fd_sc_hd__a21oi_1 _23816_ (.A1(_02225_),
    .A2(_04111_),
    .B1(_04112_),
    .Y(_04113_));
 sky130_fd_sc_hd__a221oi_1 _23817_ (.A1(net1259),
    .A2(_01929_),
    .B1(_04109_),
    .B2(_01734_),
    .C1(_04113_),
    .Y(_04114_));
 sky130_fd_sc_hd__nand2_1 _23818_ (.A(net739),
    .B(_04114_),
    .Y(_04115_));
 sky130_fd_sc_hd__a21oi_4 _23819_ (.A1(_04107_),
    .A2(_04115_),
    .B1(_08632_),
    .Y(_04116_));
 sky130_fd_sc_hd__a21oi_4 _23820_ (.A1(_08632_),
    .A2(_11621_),
    .B1(_04116_),
    .Y(_04117_));
 sky130_fd_sc_hd__nor2_2 _23821_ (.A(_02646_),
    .B(_04117_),
    .Y(_04118_));
 sky130_fd_sc_hd__a31oi_4 _23822_ (.A1(_02646_),
    .A2(_03478_),
    .A3(_03987_),
    .B1(_04118_),
    .Y(_04119_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_282 ();
 sky130_fd_sc_hd__nand2_1 _23824_ (.A(_02119_),
    .B(net1585),
    .Y(_04121_));
 sky130_fd_sc_hd__nand2_1 _23825_ (.A(\gen_regfile_ff.register_file_i.rf_reg[149] ),
    .B(_02123_),
    .Y(_04122_));
 sky130_fd_sc_hd__nand2_1 _23826_ (.A(_04121_),
    .B(_04122_),
    .Y(_00533_));
 sky130_fd_sc_hd__nand2_1 _23827_ (.A(_03719_),
    .B(_03848_),
    .Y(_04123_));
 sky130_fd_sc_hd__a21oi_4 _23828_ (.A1(net858),
    .A2(_03753_),
    .B1(_04123_),
    .Y(_04124_));
 sky130_fd_sc_hd__o22ai_4 _23829_ (.A1(_03848_),
    .A2(_03964_),
    .B1(_03842_),
    .B2(_04124_),
    .Y(_04125_));
 sky130_fd_sc_hd__a21boi_2 _23830_ (.A1(_04125_),
    .A2(_03958_),
    .B1_N(_03959_),
    .Y(_04126_));
 sky130_fd_sc_hd__o21ai_1 _23831_ (.A1(_04101_),
    .A2(_04126_),
    .B1(_04099_),
    .Y(_04127_));
 sky130_fd_sc_hd__nor2_1 _23832_ (.A(_04081_),
    .B(_04077_),
    .Y(_04128_));
 sky130_fd_sc_hd__nor2_1 _23833_ (.A(_04076_),
    .B(_04128_),
    .Y(_04129_));
 sky130_fd_sc_hd__a211oi_1 _23834_ (.A1(_04074_),
    .A2(_04129_),
    .B1(_04089_),
    .C1(_03926_),
    .Y(_04130_));
 sky130_fd_sc_hd__and2_0 _23835_ (.A(_03926_),
    .B(_04089_),
    .X(_04131_));
 sky130_fd_sc_hd__o21a_1 _23836_ (.A1(_04077_),
    .A2(_04131_),
    .B1(_04129_),
    .X(_04132_));
 sky130_fd_sc_hd__nor2_1 _23837_ (.A(_04074_),
    .B(_04132_),
    .Y(_04133_));
 sky130_fd_sc_hd__a211oi_1 _23838_ (.A1(_04074_),
    .A2(_04090_),
    .B1(_04131_),
    .C1(_04081_),
    .Y(_04134_));
 sky130_fd_sc_hd__nor3_1 _23839_ (.A(_04130_),
    .B(_04133_),
    .C(_04134_),
    .Y(_04135_));
 sky130_fd_sc_hd__maj3_2 _23840_ (.A(_04015_),
    .B(_04019_),
    .C(_04040_),
    .X(_04136_));
 sky130_fd_sc_hd__nor2_1 _23841_ (.A(net1413),
    .B(_02932_),
    .Y(_04137_));
 sky130_fd_sc_hd__nor2_1 _23842_ (.A(_03142_),
    .B(net1243),
    .Y(_04138_));
 sky130_fd_sc_hd__nor2_1 _23843_ (.A(_02936_),
    .B(net1240),
    .Y(_04139_));
 sky130_fd_sc_hd__xnor3_1 _23844_ (.A(_04137_),
    .B(_04138_),
    .C(_04139_),
    .X(_04140_));
 sky130_fd_sc_hd__a221oi_4 _23845_ (.A1(net1165),
    .A2(net322),
    .B1(net1035),
    .B2(_02503_),
    .C1(_03160_),
    .Y(_04141_));
 sky130_fd_sc_hd__o211a_1 _23846_ (.A1(net979),
    .A2(net322),
    .B1(_02918_),
    .C1(_03309_),
    .X(_04142_));
 sky130_fd_sc_hd__xnor2_1 _23847_ (.A(_04141_),
    .B(_04142_),
    .Y(_04143_));
 sky130_fd_sc_hd__nand2_1 _23848_ (.A(net1069),
    .B(_03384_),
    .Y(_04144_));
 sky130_fd_sc_hd__xnor2_2 _23849_ (.A(_04143_),
    .B(_04144_),
    .Y(_04145_));
 sky130_fd_sc_hd__maj3_1 _23850_ (.A(_03994_),
    .B(_03995_),
    .C(_03993_),
    .X(_04146_));
 sky130_fd_sc_hd__xor3_1 _23851_ (.A(_04140_),
    .B(_04145_),
    .C(_04146_),
    .X(_04147_));
 sky130_fd_sc_hd__nand2b_1 _23852_ (.A_N(net1161),
    .B(_03265_),
    .Y(_04148_));
 sky130_fd_sc_hd__a211oi_4 _23853_ (.A1(_02895_),
    .A2(_02896_),
    .B1(_02723_),
    .C1(_02725_),
    .Y(_04149_));
 sky130_fd_sc_hd__a221oi_4 _23854_ (.A1(_02619_),
    .A2(_01712_),
    .B1(_03039_),
    .B2(_03040_),
    .C1(net855),
    .Y(_04150_));
 sky130_fd_sc_hd__xnor2_1 _23855_ (.A(_04149_),
    .B(_04150_),
    .Y(_04151_));
 sky130_fd_sc_hd__xnor2_1 _23856_ (.A(_04148_),
    .B(_04151_),
    .Y(_04152_));
 sky130_fd_sc_hd__maj3_1 _23857_ (.A(_03998_),
    .B(_03999_),
    .C(_04000_),
    .X(_04153_));
 sky130_fd_sc_hd__maj3_1 _23858_ (.A(_04006_),
    .B(_04005_),
    .C(_04007_),
    .X(_04154_));
 sky130_fd_sc_hd__xnor2_1 _23859_ (.A(_04153_),
    .B(_04154_),
    .Y(_04155_));
 sky130_fd_sc_hd__xnor2_1 _23860_ (.A(_04152_),
    .B(_04155_),
    .Y(_04156_));
 sky130_fd_sc_hd__maj3_1 _23861_ (.A(_04001_),
    .B(_03997_),
    .C(_04002_),
    .X(_04157_));
 sky130_fd_sc_hd__xnor3_2 _23862_ (.A(_04147_),
    .B(_04156_),
    .C(_04157_),
    .X(_04158_));
 sky130_fd_sc_hd__maj3_1 _23863_ (.A(_04004_),
    .B(_04013_),
    .C(_04014_),
    .X(_04159_));
 sky130_fd_sc_hd__o32ai_1 _23864_ (.A1(net898),
    .A2(_03119_),
    .A3(_03512_),
    .B1(_04020_),
    .B2(_02421_),
    .Y(_04160_));
 sky130_fd_sc_hd__nor2_1 _23865_ (.A(net1010),
    .B(_04020_),
    .Y(_04161_));
 sky130_fd_sc_hd__nor3_1 _23866_ (.A(_02289_),
    .B(_02421_),
    .C(_03512_),
    .Y(_04162_));
 sky130_fd_sc_hd__nor2_1 _23867_ (.A(_03119_),
    .B(_03689_),
    .Y(_04163_));
 sky130_fd_sc_hd__nor4_1 _23868_ (.A(net1167),
    .B(net1010),
    .C(_03265_),
    .D(_03670_),
    .Y(_04164_));
 sky130_fd_sc_hd__o21ai_0 _23869_ (.A1(_04163_),
    .A2(_04164_),
    .B1(net898),
    .Y(_04165_));
 sky130_fd_sc_hd__o21ai_1 _23870_ (.A1(_04161_),
    .A2(_04162_),
    .B1(_04165_),
    .Y(_04166_));
 sky130_fd_sc_hd__a21oi_2 _23871_ (.A1(net1167),
    .A2(_04160_),
    .B1(_04166_),
    .Y(_04167_));
 sky130_fd_sc_hd__maj3_1 _23872_ (.A(_04010_),
    .B(_04009_),
    .C(_04011_),
    .X(_04168_));
 sky130_fd_sc_hd__o41ai_1 _23873_ (.A1(_03883_),
    .A2(_03884_),
    .A3(_03885_),
    .A4(_03886_),
    .B1(_03428_),
    .Y(_04169_));
 sky130_fd_sc_hd__nand2_1 _23874_ (.A(_02421_),
    .B(_03265_),
    .Y(_04170_));
 sky130_fd_sc_hd__a211oi_1 _23875_ (.A1(_03271_),
    .A2(_03273_),
    .B1(_02299_),
    .C1(_02300_),
    .Y(_04171_));
 sky130_fd_sc_hd__o211ai_2 _23876_ (.A1(net915),
    .A2(net321),
    .B1(_02307_),
    .C1(_03428_),
    .Y(_04172_));
 sky130_fd_sc_hd__mux2i_4 _23877_ (.A0(_02289_),
    .A1(_04171_),
    .S(_04172_),
    .Y(_04173_));
 sky130_fd_sc_hd__xnor2_1 _23878_ (.A(_04170_),
    .B(_04173_),
    .Y(_04174_));
 sky130_fd_sc_hd__maj3_1 _23879_ (.A(_03890_),
    .B(_03891_),
    .C(_03893_),
    .X(_04175_));
 sky130_fd_sc_hd__maj3_2 _23880_ (.A(_04169_),
    .B(_04174_),
    .C(_04175_),
    .X(_04176_));
 sky130_fd_sc_hd__xnor2_1 _23881_ (.A(_04168_),
    .B(_04176_),
    .Y(_04177_));
 sky130_fd_sc_hd__xnor3_1 _23882_ (.A(_04035_),
    .B(_04167_),
    .C(_04177_),
    .X(_04178_));
 sky130_fd_sc_hd__xnor2_1 _23883_ (.A(_04159_),
    .B(_04178_),
    .Y(_04179_));
 sky130_fd_sc_hd__xnor2_2 _23884_ (.A(_04158_),
    .B(_04179_),
    .Y(_04180_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_281 ();
 sky130_fd_sc_hd__nand2_8 _23886_ (.A(_03689_),
    .B(_03936_),
    .Y(_04182_));
 sky130_fd_sc_hd__a21o_1 _23887_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[53] ),
    .A2(_08292_),
    .B1(_03778_),
    .X(_04183_));
 sky130_fd_sc_hd__a21oi_2 _23888_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[52] ),
    .A2(_08292_),
    .B1(_03778_),
    .Y(_04184_));
 sky130_fd_sc_hd__nand2_1 _23889_ (.A(_03516_),
    .B(_04184_),
    .Y(_04185_));
 sky130_fd_sc_hd__maj3_1 _23890_ (.A(_04182_),
    .B(_04183_),
    .C(_04185_),
    .X(_04186_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_279 ();
 sky130_fd_sc_hd__a21oi_1 _23893_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[53] ),
    .A2(_03509_),
    .B1(_03684_),
    .Y(_04189_));
 sky130_fd_sc_hd__nor2_2 _23894_ (.A(_03516_),
    .B(_04182_),
    .Y(_04190_));
 sky130_fd_sc_hd__a211oi_1 _23895_ (.A1(_04182_),
    .A2(_04189_),
    .B1(_04190_),
    .C1(_03695_),
    .Y(_04191_));
 sky130_fd_sc_hd__a21oi_2 _23896_ (.A1(_03695_),
    .A2(_04186_),
    .B1(_04191_),
    .Y(_04192_));
 sky130_fd_sc_hd__a21oi_4 _23897_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[54] ),
    .A2(_08292_),
    .B1(_03778_),
    .Y(_04193_));
 sky130_fd_sc_hd__xnor2_2 _23898_ (.A(_04192_),
    .B(_04193_),
    .Y(_04194_));
 sky130_fd_sc_hd__xnor2_1 _23899_ (.A(_04033_),
    .B(_04035_),
    .Y(_04195_));
 sky130_fd_sc_hd__nor2b_1 _23900_ (.A(_04038_),
    .B_N(_04036_),
    .Y(_04196_));
 sky130_fd_sc_hd__nand2b_1 _23901_ (.A_N(_04036_),
    .B(_04038_),
    .Y(_04197_));
 sky130_fd_sc_hd__o21ai_2 _23902_ (.A1(_04195_),
    .A2(_04196_),
    .B1(_04197_),
    .Y(_04198_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_278 ();
 sky130_fd_sc_hd__nand2_1 _23904_ (.A(_03690_),
    .B(_04184_),
    .Y(_04200_));
 sky130_fd_sc_hd__a21oi_1 _23905_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[51] ),
    .A2(_08292_),
    .B1(_03778_),
    .Y(_04201_));
 sky130_fd_sc_hd__a21o_1 _23906_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[52] ),
    .A2(_08292_),
    .B1(_03778_),
    .X(_04202_));
 sky130_fd_sc_hd__o21ai_0 _23907_ (.A1(_04201_),
    .A2(_04202_),
    .B1(_03695_),
    .Y(_04203_));
 sky130_fd_sc_hd__a21oi_1 _23908_ (.A1(_03516_),
    .A2(_04201_),
    .B1(_04184_),
    .Y(_04204_));
 sky130_fd_sc_hd__nor2_1 _23909_ (.A(_03698_),
    .B(_04182_),
    .Y(_04205_));
 sky130_fd_sc_hd__a32oi_1 _23910_ (.A1(_04182_),
    .A2(_04200_),
    .A3(_04203_),
    .B1(_04204_),
    .B2(_04205_),
    .Y(_04206_));
 sky130_fd_sc_hd__a21oi_1 _23911_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[53] ),
    .A2(_08292_),
    .B1(_03778_),
    .Y(_04207_));
 sky130_fd_sc_hd__a211o_1 _23912_ (.A1(_03695_),
    .A2(_04185_),
    .B1(_04207_),
    .C1(_04182_),
    .X(_04208_));
 sky130_fd_sc_hd__o21ai_2 _23913_ (.A1(_04183_),
    .A2(_04206_),
    .B1(_04208_),
    .Y(_04209_));
 sky130_fd_sc_hd__inv_1 _23914_ (.A(_04209_),
    .Y(_04210_));
 sky130_fd_sc_hd__xnor2_1 _23915_ (.A(_04198_),
    .B(_04210_),
    .Y(_04211_));
 sky130_fd_sc_hd__xnor2_1 _23916_ (.A(_04194_),
    .B(_04211_),
    .Y(_04212_));
 sky130_fd_sc_hd__xnor3_1 _23917_ (.A(_04136_),
    .B(_04180_),
    .C(_04212_),
    .X(_04213_));
 sky130_fd_sc_hd__inv_1 _23918_ (.A(_04213_),
    .Y(_04214_));
 sky130_fd_sc_hd__or2_0 _23919_ (.A(_04041_),
    .B(_04072_),
    .X(_04215_));
 sky130_fd_sc_hd__a21o_1 _23920_ (.A1(_03933_),
    .A2(_04060_),
    .B1(_04069_),
    .X(_04216_));
 sky130_fd_sc_hd__nor2_1 _23921_ (.A(_04054_),
    .B(_04216_),
    .Y(_04217_));
 sky130_fd_sc_hd__inv_1 _23922_ (.A(_04217_),
    .Y(_04218_));
 sky130_fd_sc_hd__nand2_1 _23923_ (.A(_04041_),
    .B(_04072_),
    .Y(_04219_));
 sky130_fd_sc_hd__nand2_1 _23924_ (.A(_04054_),
    .B(_04216_),
    .Y(_04220_));
 sky130_fd_sc_hd__nor2_1 _23925_ (.A(_04041_),
    .B(_04072_),
    .Y(_04221_));
 sky130_fd_sc_hd__o21ai_0 _23926_ (.A1(_04070_),
    .A2(_04221_),
    .B1(_04219_),
    .Y(_04222_));
 sky130_fd_sc_hd__o22ai_1 _23927_ (.A1(_04216_),
    .A2(_04215_),
    .B1(_04222_),
    .B2(_04054_),
    .Y(_04223_));
 sky130_fd_sc_hd__inv_1 _23928_ (.A(_04219_),
    .Y(_04224_));
 sky130_fd_sc_hd__inv_1 _23929_ (.A(_04043_),
    .Y(_04225_));
 sky130_fd_sc_hd__a221oi_1 _23930_ (.A1(_04216_),
    .A2(_04224_),
    .B1(_04222_),
    .B2(_04054_),
    .C1(_04225_),
    .Y(_04226_));
 sky130_fd_sc_hd__o21bai_1 _23931_ (.A1(_04043_),
    .A2(_04223_),
    .B1_N(_04226_),
    .Y(_04227_));
 sky130_fd_sc_hd__o221ai_1 _23932_ (.A1(_04215_),
    .A2(_04218_),
    .B1(_04219_),
    .B2(_04220_),
    .C1(_04227_),
    .Y(_04228_));
 sky130_fd_sc_hd__xnor2_1 _23933_ (.A(_04214_),
    .B(_04228_),
    .Y(_04229_));
 sky130_fd_sc_hd__or2_1 _23934_ (.A(_04135_),
    .B(_04229_),
    .X(_04230_));
 sky130_fd_sc_hd__nand2_1 _23935_ (.A(_04135_),
    .B(_04229_),
    .Y(_04231_));
 sky130_fd_sc_hd__nand2_1 _23936_ (.A(_04230_),
    .B(_04231_),
    .Y(_04232_));
 sky130_fd_sc_hd__xnor2_1 _23937_ (.A(_04232_),
    .B(_04127_),
    .Y(_04233_));
 sky130_fd_sc_hd__nor2_1 _23938_ (.A(_01698_),
    .B(_04233_),
    .Y(_04234_));
 sky130_fd_sc_hd__a21oi_2 _23939_ (.A1(_01698_),
    .A2(_02345_),
    .B1(_04234_),
    .Y(_04235_));
 sky130_fd_sc_hd__nand2_1 _23940_ (.A(net441),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[54] ),
    .Y(_04236_));
 sky130_fd_sc_hd__o21ai_4 _23941_ (.A1(_04235_),
    .A2(net441),
    .B1(_04236_),
    .Y(_04237_));
 sky130_fd_sc_hd__nor2_1 _23942_ (.A(_01762_),
    .B(_02561_),
    .Y(_04238_));
 sky130_fd_sc_hd__a21oi_1 _23943_ (.A1(_01762_),
    .A2(_02567_),
    .B1(_04238_),
    .Y(_04239_));
 sky130_fd_sc_hd__nor2_1 _23944_ (.A(_10205_),
    .B(_01898_),
    .Y(_04240_));
 sky130_fd_sc_hd__a22oi_1 _23945_ (.A1(_10205_),
    .A2(_01896_),
    .B1(_04240_),
    .B2(_10172_),
    .Y(_04241_));
 sky130_fd_sc_hd__nor2_1 _23946_ (.A(_10205_),
    .B(_01903_),
    .Y(_04242_));
 sky130_fd_sc_hd__o22ai_1 _23947_ (.A1(_01893_),
    .A2(_04241_),
    .B1(_04242_),
    .B2(_10172_),
    .Y(_04243_));
 sky130_fd_sc_hd__o21ai_0 _23948_ (.A1(_01761_),
    .A2(_04239_),
    .B1(_04243_),
    .Y(_04244_));
 sky130_fd_sc_hd__a21oi_1 _23949_ (.A1(net1547),
    .A2(_01929_),
    .B1(_04244_),
    .Y(_04245_));
 sky130_fd_sc_hd__nor2_1 _23950_ (.A(net314),
    .B(_04245_),
    .Y(_04246_));
 sky130_fd_sc_hd__a21oi_4 _23951_ (.A1(_04237_),
    .A2(net314),
    .B1(_04246_),
    .Y(_04247_));
 sky130_fd_sc_hd__nor2_8 _23952_ (.A(_04247_),
    .B(_08632_),
    .Y(_04248_));
 sky130_fd_sc_hd__mux4_1 _23953_ (.A0(net41),
    .A1(net55),
    .A2(\load_store_unit_i.rdata_q[30] ),
    .A3(net32),
    .S0(\load_store_unit_i.rdata_offset_q[1] ),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .X(_04249_));
 sky130_fd_sc_hd__nand2_1 _23954_ (.A(_01674_),
    .B(_04249_),
    .Y(_04250_));
 sky130_fd_sc_hd__nand3_1 _23955_ (.A(_02646_),
    .B(_03478_),
    .C(_04250_),
    .Y(_04251_));
 sky130_fd_sc_hd__o31a_4 _23956_ (.A1(_04248_),
    .A2(_02646_),
    .A3(_11641_),
    .B1(_04251_),
    .X(_04252_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_277 ();
 sky130_fd_sc_hd__mux2_4 _23958_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[150] ),
    .A1(_04252_),
    .S(_02119_),
    .X(_00534_));
 sky130_fd_sc_hd__mux2i_1 _23959_ (.A0(\load_store_unit_i.rdata_q[31] ),
    .A1(net33),
    .S(\load_store_unit_i.rdata_offset_q[1] ),
    .Y(_04254_));
 sky130_fd_sc_hd__nand2_1 _23960_ (.A(\load_store_unit_i.rdata_offset_q[0] ),
    .B(_04254_),
    .Y(_04255_));
 sky130_fd_sc_hd__o211ai_2 _23961_ (.A1(\load_store_unit_i.rdata_offset_q[0] ),
    .A2(_03475_),
    .B1(_04255_),
    .C1(_01674_),
    .Y(_04256_));
 sky130_fd_sc_hd__o21a_1 _23962_ (.A1(_04213_),
    .A2(_04217_),
    .B1(_04225_),
    .X(_04257_));
 sky130_fd_sc_hd__a21oi_1 _23963_ (.A1(_04213_),
    .A2(_04220_),
    .B1(_04257_),
    .Y(_04258_));
 sky130_fd_sc_hd__a21oi_1 _23964_ (.A1(_04225_),
    .A2(_04220_),
    .B1(_04217_),
    .Y(_04259_));
 sky130_fd_sc_hd__maj3_1 _23965_ (.A(_04214_),
    .B(_04215_),
    .C(_04259_),
    .X(_04260_));
 sky130_fd_sc_hd__o21ai_1 _23966_ (.A1(_04224_),
    .A2(_04258_),
    .B1(_04260_),
    .Y(_04261_));
 sky130_fd_sc_hd__o211ai_1 _23967_ (.A1(_03265_),
    .A2(_03428_),
    .B1(_04027_),
    .C1(_03274_),
    .Y(_04262_));
 sky130_fd_sc_hd__o21ai_0 _23968_ (.A1(_03889_),
    .A2(_04167_),
    .B1(_04262_),
    .Y(_04263_));
 sky130_fd_sc_hd__o32ai_1 _23969_ (.A1(net1168),
    .A2(_03889_),
    .A3(_04166_),
    .B1(_04262_),
    .B2(_03689_),
    .Y(_04264_));
 sky130_fd_sc_hd__a21oi_2 _23970_ (.A1(net1169),
    .A2(_04263_),
    .B1(_04264_),
    .Y(_04265_));
 sky130_fd_sc_hd__nand2_1 _23971_ (.A(_04153_),
    .B(_04154_),
    .Y(_04266_));
 sky130_fd_sc_hd__nor2_1 _23972_ (.A(_04153_),
    .B(_04154_),
    .Y(_04267_));
 sky130_fd_sc_hd__a21oi_2 _23973_ (.A1(_04152_),
    .A2(_04266_),
    .B1(_04267_),
    .Y(_04268_));
 sky130_fd_sc_hd__a211oi_1 _23974_ (.A1(_02289_),
    .A2(_03274_),
    .B1(net1010),
    .C1(net910),
    .Y(_04269_));
 sky130_fd_sc_hd__a31oi_2 _23975_ (.A1(net910),
    .A2(_02289_),
    .A3(net1010),
    .B1(_04269_),
    .Y(_04270_));
 sky130_fd_sc_hd__xnor2_2 _23976_ (.A(_03887_),
    .B(_04270_),
    .Y(_04271_));
 sky130_fd_sc_hd__nor2_8 _23977_ (.A(_03670_),
    .B(_04271_),
    .Y(_04272_));
 sky130_fd_sc_hd__xor2_1 _23978_ (.A(_04268_),
    .B(_04272_),
    .X(_04273_));
 sky130_fd_sc_hd__xnor2_2 _23979_ (.A(_04265_),
    .B(_04273_),
    .Y(_04274_));
 sky130_fd_sc_hd__maj3_1 _23980_ (.A(_04147_),
    .B(_04156_),
    .C(_04157_),
    .X(_04275_));
 sky130_fd_sc_hd__nor2_1 _23981_ (.A(net1239),
    .B(net899),
    .Y(_04276_));
 sky130_fd_sc_hd__nor2_1 _23982_ (.A(net1413),
    .B(net1263),
    .Y(_04277_));
 sky130_fd_sc_hd__nor2_1 _23983_ (.A(_02936_),
    .B(_03097_),
    .Y(_04278_));
 sky130_fd_sc_hd__xnor2_1 _23984_ (.A(_04277_),
    .B(_04278_),
    .Y(_04279_));
 sky130_fd_sc_hd__xnor2_1 _23985_ (.A(_04276_),
    .B(_04279_),
    .Y(_04280_));
 sky130_fd_sc_hd__nor2_1 _23986_ (.A(_04141_),
    .B(_04142_),
    .Y(_04281_));
 sky130_fd_sc_hd__nand2_1 _23987_ (.A(_04141_),
    .B(_04142_),
    .Y(_04282_));
 sky130_fd_sc_hd__o21ai_0 _23988_ (.A1(_04144_),
    .A2(_04281_),
    .B1(_04282_),
    .Y(_04283_));
 sky130_fd_sc_hd__inv_1 _23989_ (.A(_04283_),
    .Y(_04284_));
 sky130_fd_sc_hd__nand2_1 _23990_ (.A(_02589_),
    .B(_03161_),
    .Y(_04285_));
 sky130_fd_sc_hd__nand2_1 _23991_ (.A(_03004_),
    .B(_03310_),
    .Y(_04286_));
 sky130_fd_sc_hd__xor2_1 _23992_ (.A(_04285_),
    .B(_04286_),
    .X(_04287_));
 sky130_fd_sc_hd__nand2_1 _23993_ (.A(net1228),
    .B(_03376_),
    .Y(_04288_));
 sky130_fd_sc_hd__xor2_1 _23994_ (.A(_04287_),
    .B(_04288_),
    .X(_04289_));
 sky130_fd_sc_hd__xnor2_1 _23995_ (.A(_04284_),
    .B(_04289_),
    .Y(_04290_));
 sky130_fd_sc_hd__maj3_1 _23996_ (.A(_04140_),
    .B(_04145_),
    .C(_04146_),
    .X(_04291_));
 sky130_fd_sc_hd__maj3_1 _23997_ (.A(_04137_),
    .B(_04138_),
    .C(_04139_),
    .X(_04292_));
 sky130_fd_sc_hd__nor2_1 _23998_ (.A(net1161),
    .B(_04020_),
    .Y(_04293_));
 sky130_fd_sc_hd__nor2_1 _23999_ (.A(net1158),
    .B(_03100_),
    .Y(_04294_));
 sky130_fd_sc_hd__nor2_1 _24000_ (.A(net1173),
    .B(_03119_),
    .Y(_04295_));
 sky130_fd_sc_hd__xnor3_1 _24001_ (.A(_04293_),
    .B(_04294_),
    .C(_04295_),
    .X(_04296_));
 sky130_fd_sc_hd__nor2_1 _24002_ (.A(_04149_),
    .B(_04150_),
    .Y(_04297_));
 sky130_fd_sc_hd__nand2_1 _24003_ (.A(_04149_),
    .B(_04150_),
    .Y(_04298_));
 sky130_fd_sc_hd__o21ai_2 _24004_ (.A1(_04148_),
    .A2(_04297_),
    .B1(_04298_),
    .Y(_04299_));
 sky130_fd_sc_hd__xnor3_1 _24005_ (.A(_04292_),
    .B(_04296_),
    .C(_04299_),
    .X(_04300_));
 sky130_fd_sc_hd__xor2_1 _24006_ (.A(_04291_),
    .B(_04300_),
    .X(_04301_));
 sky130_fd_sc_hd__xnor3_1 _24007_ (.A(_04280_),
    .B(_04290_),
    .C(_04301_),
    .X(_04302_));
 sky130_fd_sc_hd__nor2_2 _24008_ (.A(_04275_),
    .B(_04302_),
    .Y(_04303_));
 sky130_fd_sc_hd__and2_1 _24009_ (.A(_04275_),
    .B(_04302_),
    .X(_04304_));
 sky130_fd_sc_hd__nor2_1 _24010_ (.A(_04303_),
    .B(_04304_),
    .Y(_04305_));
 sky130_fd_sc_hd__xor2_2 _24011_ (.A(_04274_),
    .B(_04305_),
    .X(_04306_));
 sky130_fd_sc_hd__nor2_1 _24012_ (.A(_04159_),
    .B(_04178_),
    .Y(_04307_));
 sky130_fd_sc_hd__nand2_1 _24013_ (.A(_04159_),
    .B(_04178_),
    .Y(_04308_));
 sky130_fd_sc_hd__o21a_1 _24014_ (.A1(_04158_),
    .A2(_04307_),
    .B1(_04308_),
    .X(_04309_));
 sky130_fd_sc_hd__o21a_1 _24015_ (.A1(_04010_),
    .A2(_04011_),
    .B1(_04009_),
    .X(_04310_));
 sky130_fd_sc_hd__a21oi_1 _24016_ (.A1(_04010_),
    .A2(_04011_),
    .B1(_04310_),
    .Y(_04311_));
 sky130_fd_sc_hd__xnor2_1 _24017_ (.A(_04035_),
    .B(_04167_),
    .Y(_04312_));
 sky130_fd_sc_hd__maj3_4 _24018_ (.A(_04311_),
    .B(_04312_),
    .C(_04176_),
    .X(_04313_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_276 ();
 sky130_fd_sc_hd__nand2_1 _24020_ (.A(_03695_),
    .B(_04061_),
    .Y(_04315_));
 sky130_fd_sc_hd__nand2_1 _24021_ (.A(_04183_),
    .B(_04193_),
    .Y(_04316_));
 sky130_fd_sc_hd__nor2_1 _24022_ (.A(_04182_),
    .B(_04193_),
    .Y(_04317_));
 sky130_fd_sc_hd__nor2_1 _24023_ (.A(_04061_),
    .B(_04316_),
    .Y(_04318_));
 sky130_fd_sc_hd__o21ai_0 _24024_ (.A1(_04317_),
    .A2(_04318_),
    .B1(_03698_),
    .Y(_04319_));
 sky130_fd_sc_hd__o21ai_0 _24025_ (.A1(_04315_),
    .A2(_04316_),
    .B1(_04319_),
    .Y(_04320_));
 sky130_fd_sc_hd__nand3_1 _24026_ (.A(_04182_),
    .B(_04202_),
    .C(_04193_),
    .Y(_04321_));
 sky130_fd_sc_hd__o21ai_0 _24027_ (.A1(_04182_),
    .A2(_04193_),
    .B1(_04321_),
    .Y(_04322_));
 sky130_fd_sc_hd__nand2_1 _24028_ (.A(_04061_),
    .B(_04193_),
    .Y(_04323_));
 sky130_fd_sc_hd__or3_1 _24029_ (.A(_04061_),
    .B(_04183_),
    .C(_04193_),
    .X(_04324_));
 sky130_fd_sc_hd__a21oi_1 _24030_ (.A1(_04323_),
    .A2(_04324_),
    .B1(_03695_),
    .Y(_04325_));
 sky130_fd_sc_hd__a31oi_1 _24031_ (.A1(_03695_),
    .A2(_04207_),
    .A3(_04322_),
    .B1(_04325_),
    .Y(_04326_));
 sky130_fd_sc_hd__o311ai_1 _24032_ (.A1(_04182_),
    .A2(_04184_),
    .A3(_04316_),
    .B1(_04326_),
    .C1(_03516_),
    .Y(_04327_));
 sky130_fd_sc_hd__o21ai_2 _24033_ (.A1(_03516_),
    .A2(_04320_),
    .B1(_04327_),
    .Y(_04328_));
 sky130_fd_sc_hd__o211ai_1 _24034_ (.A1(_04061_),
    .A2(_04193_),
    .B1(_04207_),
    .C1(_03516_),
    .Y(_04329_));
 sky130_fd_sc_hd__a21oi_2 _24035_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[54] ),
    .A2(_03509_),
    .B1(_03684_),
    .Y(_04330_));
 sky130_fd_sc_hd__a211oi_1 _24036_ (.A1(_04182_),
    .A2(_04330_),
    .B1(_04190_),
    .C1(_03695_),
    .Y(_04331_));
 sky130_fd_sc_hd__a31oi_2 _24037_ (.A1(_03695_),
    .A2(_04323_),
    .A3(_04329_),
    .B1(_04331_),
    .Y(_04332_));
 sky130_fd_sc_hd__a21oi_1 _24038_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[55] ),
    .A2(_08292_),
    .B1(_03778_),
    .Y(_04333_));
 sky130_fd_sc_hd__xnor2_2 _24039_ (.A(_04332_),
    .B(_04333_),
    .Y(_04334_));
 sky130_fd_sc_hd__inv_1 _24040_ (.A(_04334_),
    .Y(_04335_));
 sky130_fd_sc_hd__xnor2_1 _24041_ (.A(_04328_),
    .B(_04335_),
    .Y(_04336_));
 sky130_fd_sc_hd__xnor2_1 _24042_ (.A(_04313_),
    .B(_04336_),
    .Y(_04337_));
 sky130_fd_sc_hd__xnor2_1 _24043_ (.A(_04309_),
    .B(_04337_),
    .Y(_04338_));
 sky130_fd_sc_hd__xnor2_2 _24044_ (.A(_04306_),
    .B(_04338_),
    .Y(_04339_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_272 ();
 sky130_fd_sc_hd__a21oi_1 _24049_ (.A1(_03927_),
    .A2(_03939_),
    .B1(_03941_),
    .Y(_04344_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_269 ();
 sky130_fd_sc_hd__a21oi_1 _24053_ (.A1(_03942_),
    .A2(_03939_),
    .B1(_03941_),
    .Y(_04348_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_268 ();
 sky130_fd_sc_hd__o32a_1 _24055_ (.A1(_03670_),
    .A2(_03515_),
    .A3(_04348_),
    .B1(_03939_),
    .B2(_03933_),
    .X(_04350_));
 sky130_fd_sc_hd__nor2_1 _24056_ (.A(_03937_),
    .B(_04350_),
    .Y(_04351_));
 sky130_fd_sc_hd__nand2_4 _24057_ (.A(_03933_),
    .B(_03937_),
    .Y(_04352_));
 sky130_fd_sc_hd__a211oi_1 _24058_ (.A1(_03927_),
    .A2(_03773_),
    .B1(_03939_),
    .C1(_04352_),
    .Y(_04353_));
 sky130_fd_sc_hd__o21ai_0 _24059_ (.A1(_04351_),
    .A2(_04353_),
    .B1(_04046_),
    .Y(_04354_));
 sky130_fd_sc_hd__o31ai_2 _24060_ (.A1(_04049_),
    .A2(_04046_),
    .A3(_04344_),
    .B1(_04354_),
    .Y(_04355_));
 sky130_fd_sc_hd__nor2_1 _24061_ (.A(_04180_),
    .B(_04198_),
    .Y(_04356_));
 sky130_fd_sc_hd__and2_1 _24062_ (.A(_04180_),
    .B(_04198_),
    .X(_04357_));
 sky130_fd_sc_hd__xnor2_1 _24063_ (.A(_04192_),
    .B(_04330_),
    .Y(_04358_));
 sky130_fd_sc_hd__nor2_1 _24064_ (.A(_04357_),
    .B(_04358_),
    .Y(_04359_));
 sky130_fd_sc_hd__nand2_1 _24065_ (.A(_04357_),
    .B(_04358_),
    .Y(_04360_));
 sky130_fd_sc_hd__o31ai_1 _24066_ (.A1(_04136_),
    .A2(_04356_),
    .A3(_04359_),
    .B1(_04360_),
    .Y(_04361_));
 sky130_fd_sc_hd__nor4_1 _24067_ (.A(_04180_),
    .B(_04198_),
    .C(_04194_),
    .D(_04209_),
    .Y(_04362_));
 sky130_fd_sc_hd__nor2_1 _24068_ (.A(_04194_),
    .B(_04209_),
    .Y(_04363_));
 sky130_fd_sc_hd__nand2_1 _24069_ (.A(_04136_),
    .B(_04363_),
    .Y(_04364_));
 sky130_fd_sc_hd__xor2_1 _24070_ (.A(_04192_),
    .B(_04193_),
    .X(_04365_));
 sky130_fd_sc_hd__nor2_1 _24071_ (.A(_04136_),
    .B(_04365_),
    .Y(_04366_));
 sky130_fd_sc_hd__nand2_1 _24072_ (.A(_04357_),
    .B(_04366_),
    .Y(_04367_));
 sky130_fd_sc_hd__o211ai_1 _24073_ (.A1(_04365_),
    .A2(_04210_),
    .B1(_04136_),
    .C1(_04356_),
    .Y(_04368_));
 sky130_fd_sc_hd__o211ai_1 _24074_ (.A1(_04357_),
    .A2(_04364_),
    .B1(_04367_),
    .C1(_04368_),
    .Y(_04369_));
 sky130_fd_sc_hd__a211oi_1 _24075_ (.A1(_04355_),
    .A2(_04361_),
    .B1(_04362_),
    .C1(_04369_),
    .Y(_04370_));
 sky130_fd_sc_hd__xor2_1 _24076_ (.A(_04339_),
    .B(_04370_),
    .X(_04371_));
 sky130_fd_sc_hd__xnor2_1 _24077_ (.A(_04261_),
    .B(_04371_),
    .Y(_04372_));
 sky130_fd_sc_hd__nor2_4 _24078_ (.A(_03992_),
    .B(_04101_),
    .Y(_04373_));
 sky130_fd_sc_hd__o21ai_1 _24079_ (.A1(_04100_),
    .A2(_04373_),
    .B1(_04231_),
    .Y(_04374_));
 sky130_fd_sc_hd__nand2_1 _24080_ (.A(_04230_),
    .B(_04374_),
    .Y(_04375_));
 sky130_fd_sc_hd__xor2_2 _24081_ (.A(_04372_),
    .B(_04375_),
    .X(_04376_));
 sky130_fd_sc_hd__nand2_2 _24082_ (.A(_02169_),
    .B(_04376_),
    .Y(_04377_));
 sky130_fd_sc_hd__o21ai_4 _24083_ (.A1(_02169_),
    .A2(_02451_),
    .B1(_04377_),
    .Y(_04378_));
 sky130_fd_sc_hd__mux2i_4 _24084_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[55] ),
    .A1(_04378_),
    .S(_08100_),
    .Y(_04379_));
 sky130_fd_sc_hd__nor2_1 _24085_ (.A(_01762_),
    .B(_02476_),
    .Y(_04380_));
 sky130_fd_sc_hd__a21oi_1 _24086_ (.A1(_01762_),
    .A2(_02472_),
    .B1(_04380_),
    .Y(_04381_));
 sky130_fd_sc_hd__nor3_1 _24087_ (.A(_10266_),
    .B(_10272_),
    .C(_01898_),
    .Y(_04382_));
 sky130_fd_sc_hd__a21oi_1 _24088_ (.A1(_10266_),
    .A2(_01896_),
    .B1(_04382_),
    .Y(_04383_));
 sky130_fd_sc_hd__o21ai_0 _24089_ (.A1(_10266_),
    .A2(_01903_),
    .B1(_10272_),
    .Y(_04384_));
 sky130_fd_sc_hd__o21ai_0 _24090_ (.A1(_01893_),
    .A2(_04383_),
    .B1(_04384_),
    .Y(_04385_));
 sky130_fd_sc_hd__o21ai_0 _24091_ (.A1(_01761_),
    .A2(_04381_),
    .B1(_04385_),
    .Y(_04386_));
 sky130_fd_sc_hd__a211oi_1 _24092_ (.A1(net164),
    .A2(_01929_),
    .B1(_04386_),
    .C1(net1103),
    .Y(_04387_));
 sky130_fd_sc_hd__a21oi_4 _24093_ (.A1(_04379_),
    .A2(net1103),
    .B1(_04387_),
    .Y(_04388_));
 sky130_fd_sc_hd__nor3_4 _24094_ (.A(_11661_),
    .B(_02646_),
    .C(_04388_),
    .Y(_04389_));
 sky130_fd_sc_hd__a31oi_4 _24095_ (.A1(_02646_),
    .A2(_03478_),
    .A3(_04256_),
    .B1(_04389_),
    .Y(_04390_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_267 ();
 sky130_fd_sc_hd__nand2_1 _24097_ (.A(_04390_),
    .B(_02119_),
    .Y(_04392_));
 sky130_fd_sc_hd__nand2_1 _24098_ (.A(\gen_regfile_ff.register_file_i.rf_reg[151] ),
    .B(_02123_),
    .Y(_04393_));
 sky130_fd_sc_hd__nand2_1 _24099_ (.A(_04392_),
    .B(_04393_),
    .Y(_00535_));
 sky130_fd_sc_hd__nand2_1 _24100_ (.A(_01916_),
    .B(_02849_),
    .Y(_04394_));
 sky130_fd_sc_hd__nand2_1 _24101_ (.A(\gen_regfile_ff.register_file_i.rf_reg[43] ),
    .B(_01921_),
    .Y(_04395_));
 sky130_fd_sc_hd__nand2_1 _24102_ (.A(_04394_),
    .B(_04395_),
    .Y(_00536_));
 sky130_fd_sc_hd__mux4_1 _24103_ (.A0(net43),
    .A1(net57),
    .A2(net27),
    .A3(net34),
    .S0(\load_store_unit_i.rdata_offset_q[1] ),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .X(_04396_));
 sky130_fd_sc_hd__a21oi_1 _24104_ (.A1(_01674_),
    .A2(_04396_),
    .B1(_03479_),
    .Y(_04397_));
 sky130_fd_sc_hd__nand3_1 _24105_ (.A(_10368_),
    .B(_10396_),
    .C(_02228_),
    .Y(_04398_));
 sky130_fd_sc_hd__o21ai_0 _24106_ (.A1(_10368_),
    .A2(_01902_),
    .B1(_04398_),
    .Y(_04399_));
 sky130_fd_sc_hd__a21oi_1 _24107_ (.A1(_10368_),
    .A2(_02233_),
    .B1(_10396_),
    .Y(_04400_));
 sky130_fd_sc_hd__a21oi_1 _24108_ (.A1(_02225_),
    .A2(_04399_),
    .B1(_04400_),
    .Y(_04401_));
 sky130_fd_sc_hd__nor2_1 _24109_ (.A(_01762_),
    .B(_02378_),
    .Y(_04402_));
 sky130_fd_sc_hd__a21oi_1 _24110_ (.A1(_01762_),
    .A2(_02377_),
    .B1(_04402_),
    .Y(_04403_));
 sky130_fd_sc_hd__nor2_1 _24111_ (.A(_01761_),
    .B(_04403_),
    .Y(_04404_));
 sky130_fd_sc_hd__nand3_1 _24112_ (.A(_08290_),
    .B(_11682_),
    .C(net1483),
    .Y(_04405_));
 sky130_fd_sc_hd__a2111oi_4 _24113_ (.A1(net774),
    .A2(_01929_),
    .B1(_04401_),
    .C1(_04404_),
    .D1(_04405_),
    .Y(_04406_));
 sky130_fd_sc_hd__o21a_1 _24114_ (.A1(_04261_),
    .A2(_04371_),
    .B1(_04231_),
    .X(_04407_));
 sky130_fd_sc_hd__nand2_1 _24115_ (.A(_03959_),
    .B(_04099_),
    .Y(_04408_));
 sky130_fd_sc_hd__a21oi_2 _24116_ (.A1(_03958_),
    .A2(_04125_),
    .B1(_04408_),
    .Y(_04409_));
 sky130_fd_sc_hd__o21ai_2 _24117_ (.A1(_04409_),
    .A2(_04101_),
    .B1(_04230_),
    .Y(_04410_));
 sky130_fd_sc_hd__nand2_1 _24118_ (.A(_04261_),
    .B(_04371_),
    .Y(_04411_));
 sky130_fd_sc_hd__inv_1 _24119_ (.A(_04411_),
    .Y(_04412_));
 sky130_fd_sc_hd__a21oi_2 _24120_ (.A1(_04407_),
    .A2(_04410_),
    .B1(_04412_),
    .Y(_04413_));
 sky130_fd_sc_hd__o21ai_0 _24121_ (.A1(_04356_),
    .A2(_04339_),
    .B1(_04136_),
    .Y(_04414_));
 sky130_fd_sc_hd__inv_1 _24122_ (.A(_04357_),
    .Y(_04415_));
 sky130_fd_sc_hd__nand2_1 _24123_ (.A(_04415_),
    .B(_04339_),
    .Y(_04416_));
 sky130_fd_sc_hd__a22oi_1 _24124_ (.A1(_04194_),
    .A2(_04209_),
    .B1(_04414_),
    .B2(_04416_),
    .Y(_04417_));
 sky130_fd_sc_hd__a21oi_1 _24125_ (.A1(_04136_),
    .A2(_04415_),
    .B1(_04356_),
    .Y(_04418_));
 sky130_fd_sc_hd__nor2_1 _24126_ (.A(_04339_),
    .B(_04363_),
    .Y(_04419_));
 sky130_fd_sc_hd__nor2_1 _24127_ (.A(_04418_),
    .B(_04419_),
    .Y(_04420_));
 sky130_fd_sc_hd__a211oi_1 _24128_ (.A1(_04339_),
    .A2(_04363_),
    .B1(_04417_),
    .C1(_04420_),
    .Y(_04421_));
 sky130_fd_sc_hd__inv_1 _24129_ (.A(_04304_),
    .Y(_04422_));
 sky130_fd_sc_hd__a21oi_2 _24130_ (.A1(_04274_),
    .A2(_04422_),
    .B1(_04303_),
    .Y(_04423_));
 sky130_fd_sc_hd__a21o_1 _24131_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[54] ),
    .A2(_03509_),
    .B1(_03684_),
    .X(_04424_));
 sky130_fd_sc_hd__nand2_1 _24132_ (.A(_04182_),
    .B(_04424_),
    .Y(_04425_));
 sky130_fd_sc_hd__a21oi_2 _24133_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[55] ),
    .A2(_03509_),
    .B1(_03684_),
    .Y(_04426_));
 sky130_fd_sc_hd__o21ai_0 _24134_ (.A1(_04330_),
    .A2(_04426_),
    .B1(_04061_),
    .Y(_04427_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_266 ();
 sky130_fd_sc_hd__a21oi_1 _24136_ (.A1(_04425_),
    .A2(_04427_),
    .B1(_03698_),
    .Y(_04429_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_265 ();
 sky130_fd_sc_hd__nor2_1 _24138_ (.A(_04061_),
    .B(_04426_),
    .Y(_04431_));
 sky130_fd_sc_hd__a21o_1 _24139_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[55] ),
    .A2(_03509_),
    .B1(_03684_),
    .X(_04432_));
 sky130_fd_sc_hd__nand2_1 _24140_ (.A(_04061_),
    .B(_04432_),
    .Y(_04433_));
 sky130_fd_sc_hd__nand3_1 _24141_ (.A(_03698_),
    .B(_04182_),
    .C(_04426_),
    .Y(_04434_));
 sky130_fd_sc_hd__o211ai_1 _24142_ (.A1(_03698_),
    .A2(_04433_),
    .B1(_04434_),
    .C1(_03690_),
    .Y(_04435_));
 sky130_fd_sc_hd__o31ai_2 _24143_ (.A1(_03690_),
    .A2(_04429_),
    .A3(_04431_),
    .B1(_04435_),
    .Y(_04436_));
 sky130_fd_sc_hd__a21oi_4 _24144_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[56] ),
    .A2(net311),
    .B1(_03772_),
    .Y(_04437_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_264 ();
 sky130_fd_sc_hd__a21oi_1 _24146_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[56] ),
    .A2(_03509_),
    .B1(_03684_),
    .Y(_04439_));
 sky130_fd_sc_hd__nand2_1 _24147_ (.A(_04436_),
    .B(_04439_),
    .Y(_04440_));
 sky130_fd_sc_hd__o21ai_2 _24148_ (.A1(_04436_),
    .A2(_04437_),
    .B1(_04440_),
    .Y(_04441_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_263 ();
 sky130_fd_sc_hd__nor2_1 _24150_ (.A(_04268_),
    .B(_04272_),
    .Y(_04443_));
 sky130_fd_sc_hd__nand2_1 _24151_ (.A(_04268_),
    .B(_04272_),
    .Y(_04444_));
 sky130_fd_sc_hd__o21ai_1 _24152_ (.A1(_04265_),
    .A2(_04443_),
    .B1(_04444_),
    .Y(_04445_));
 sky130_fd_sc_hd__o21ai_0 _24153_ (.A1(_04189_),
    .A2(_04330_),
    .B1(_03695_),
    .Y(_04446_));
 sky130_fd_sc_hd__a21o_1 _24154_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[53] ),
    .A2(_03509_),
    .B1(_03684_),
    .X(_04447_));
 sky130_fd_sc_hd__nor2_1 _24155_ (.A(_03698_),
    .B(_04432_),
    .Y(_04448_));
 sky130_fd_sc_hd__nor2_1 _24156_ (.A(_03695_),
    .B(_04426_),
    .Y(_04449_));
 sky130_fd_sc_hd__a21oi_1 _24157_ (.A1(_04447_),
    .A2(_04448_),
    .B1(_04449_),
    .Y(_04450_));
 sky130_fd_sc_hd__o22ai_1 _24158_ (.A1(_03698_),
    .A2(_04433_),
    .B1(_04450_),
    .B2(_04061_),
    .Y(_04451_));
 sky130_fd_sc_hd__a32oi_1 _24159_ (.A1(_04061_),
    .A2(_04426_),
    .A3(_04446_),
    .B1(_04451_),
    .B2(_04330_),
    .Y(_04452_));
 sky130_fd_sc_hd__nor2_1 _24160_ (.A(_04182_),
    .B(_04330_),
    .Y(_04453_));
 sky130_fd_sc_hd__nand3_1 _24161_ (.A(_04182_),
    .B(_04424_),
    .C(_04426_),
    .Y(_04454_));
 sky130_fd_sc_hd__a21oi_1 _24162_ (.A1(_04433_),
    .A2(_04454_),
    .B1(_03695_),
    .Y(_04455_));
 sky130_fd_sc_hd__a211oi_1 _24163_ (.A1(_04453_),
    .A2(_04448_),
    .B1(_04455_),
    .C1(_03516_),
    .Y(_04456_));
 sky130_fd_sc_hd__a21o_1 _24164_ (.A1(_03516_),
    .A2(_04452_),
    .B1(_04456_),
    .X(_04457_));
 sky130_fd_sc_hd__xor2_1 _24165_ (.A(_04445_),
    .B(_04457_),
    .X(_04458_));
 sky130_fd_sc_hd__xnor2_2 _24166_ (.A(_04441_),
    .B(_04458_),
    .Y(_04459_));
 sky130_fd_sc_hd__xnor2_2 _24167_ (.A(_04423_),
    .B(_04459_),
    .Y(_04460_));
 sky130_fd_sc_hd__nor2_1 _24168_ (.A(_03097_),
    .B(net899),
    .Y(_04461_));
 sky130_fd_sc_hd__nor2_1 _24169_ (.A(_02936_),
    .B(_03100_),
    .Y(_04462_));
 sky130_fd_sc_hd__nand2_1 _24170_ (.A(_02889_),
    .B(_03017_),
    .Y(_04463_));
 sky130_fd_sc_hd__xnor2_1 _24171_ (.A(_04462_),
    .B(_04463_),
    .Y(_04464_));
 sky130_fd_sc_hd__xnor2_2 _24172_ (.A(_04461_),
    .B(_04464_),
    .Y(_04465_));
 sky130_fd_sc_hd__o21a_1 _24173_ (.A1(_04285_),
    .A2(_04286_),
    .B1(_04288_),
    .X(_04466_));
 sky130_fd_sc_hd__a21oi_1 _24174_ (.A1(_04285_),
    .A2(_04286_),
    .B1(_04466_),
    .Y(_04467_));
 sky130_fd_sc_hd__nor2_1 _24175_ (.A(net1413),
    .B(_03313_),
    .Y(_04468_));
 sky130_fd_sc_hd__nor2_1 _24176_ (.A(_03142_),
    .B(_03373_),
    .Y(_04469_));
 sky130_fd_sc_hd__nand2_1 _24177_ (.A(net1004),
    .B(_03384_),
    .Y(_04470_));
 sky130_fd_sc_hd__xnor2_1 _24178_ (.A(_04469_),
    .B(_04470_),
    .Y(_04471_));
 sky130_fd_sc_hd__xnor2_1 _24179_ (.A(_04468_),
    .B(_04471_),
    .Y(_04472_));
 sky130_fd_sc_hd__xor2_1 _24180_ (.A(_04467_),
    .B(_04472_),
    .X(_04473_));
 sky130_fd_sc_hd__xnor2_2 _24181_ (.A(_04465_),
    .B(_04473_),
    .Y(_04474_));
 sky130_fd_sc_hd__xor2_1 _24182_ (.A(_04276_),
    .B(_04279_),
    .X(_04475_));
 sky130_fd_sc_hd__maj3_1 _24183_ (.A(_04475_),
    .B(_04284_),
    .C(_04289_),
    .X(_04476_));
 sky130_fd_sc_hd__nand2_1 _24184_ (.A(_02727_),
    .B(_03265_),
    .Y(_04477_));
 sky130_fd_sc_hd__nor2_1 _24185_ (.A(net1173),
    .B(_04020_),
    .Y(_04478_));
 sky130_fd_sc_hd__nor2_1 _24186_ (.A(net1161),
    .B(_03512_),
    .Y(_04479_));
 sky130_fd_sc_hd__xor2_1 _24187_ (.A(_04478_),
    .B(_04479_),
    .X(_04480_));
 sky130_fd_sc_hd__xnor2_1 _24188_ (.A(_04477_),
    .B(_04480_),
    .Y(_04481_));
 sky130_fd_sc_hd__maj3_1 _24189_ (.A(_04276_),
    .B(_04277_),
    .C(_04278_),
    .X(_04482_));
 sky130_fd_sc_hd__maj3_1 _24190_ (.A(_04293_),
    .B(_04294_),
    .C(_04295_),
    .X(_04483_));
 sky130_fd_sc_hd__xor2_1 _24191_ (.A(_04482_),
    .B(_04483_),
    .X(_04484_));
 sky130_fd_sc_hd__xnor2_1 _24192_ (.A(_04481_),
    .B(_04484_),
    .Y(_04485_));
 sky130_fd_sc_hd__nor2_1 _24193_ (.A(_04476_),
    .B(_04485_),
    .Y(_04486_));
 sky130_fd_sc_hd__and2_0 _24194_ (.A(_04476_),
    .B(_04485_),
    .X(_04487_));
 sky130_fd_sc_hd__nor2_1 _24195_ (.A(_04486_),
    .B(_04487_),
    .Y(_04488_));
 sky130_fd_sc_hd__xor2_2 _24196_ (.A(_04474_),
    .B(_04488_),
    .X(_04489_));
 sky130_fd_sc_hd__nand2b_1 _24197_ (.A_N(_04291_),
    .B(_04300_),
    .Y(_04490_));
 sky130_fd_sc_hd__xnor2_1 _24198_ (.A(_04280_),
    .B(_04290_),
    .Y(_04491_));
 sky130_fd_sc_hd__nand2b_1 _24199_ (.A_N(_04300_),
    .B(_04291_),
    .Y(_04492_));
 sky130_fd_sc_hd__nand2_1 _24200_ (.A(_04491_),
    .B(_04492_),
    .Y(_04493_));
 sky130_fd_sc_hd__nand2_1 _24201_ (.A(_04490_),
    .B(_04493_),
    .Y(_04494_));
 sky130_fd_sc_hd__nand2_1 _24202_ (.A(_04292_),
    .B(_04299_),
    .Y(_04495_));
 sky130_fd_sc_hd__nand2_1 _24203_ (.A(_04296_),
    .B(_04495_),
    .Y(_04496_));
 sky130_fd_sc_hd__o21ai_4 _24204_ (.A1(_04292_),
    .A2(_04299_),
    .B1(_04496_),
    .Y(_04497_));
 sky130_fd_sc_hd__xnor2_1 _24205_ (.A(_04494_),
    .B(_04497_),
    .Y(_04498_));
 sky130_fd_sc_hd__xnor2_2 _24206_ (.A(_04489_),
    .B(_04498_),
    .Y(_04499_));
 sky130_fd_sc_hd__nor2_2 _24207_ (.A(_03690_),
    .B(_04061_),
    .Y(_04500_));
 sky130_fd_sc_hd__nor2_8 _24208_ (.A(_04190_),
    .B(_04500_),
    .Y(_04501_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_262 ();
 sky130_fd_sc_hd__nand2_1 _24210_ (.A(_02289_),
    .B(net1010),
    .Y(_04503_));
 sky130_fd_sc_hd__nor2_1 _24211_ (.A(_03887_),
    .B(_04027_),
    .Y(_04504_));
 sky130_fd_sc_hd__nor2_1 _24212_ (.A(net911),
    .B(_04504_),
    .Y(_04505_));
 sky130_fd_sc_hd__a21oi_2 _24213_ (.A1(_03887_),
    .A2(_04503_),
    .B1(_04505_),
    .Y(_04506_));
 sky130_fd_sc_hd__nor2_4 _24214_ (.A(_03512_),
    .B(_04506_),
    .Y(_04507_));
 sky130_fd_sc_hd__xnor2_4 _24215_ (.A(_04272_),
    .B(_04507_),
    .Y(_04508_));
 sky130_fd_sc_hd__xor2_4 _24216_ (.A(_04501_),
    .B(_04508_),
    .X(_04509_));
 sky130_fd_sc_hd__xnor2_2 _24217_ (.A(_04499_),
    .B(_04509_),
    .Y(_04510_));
 sky130_fd_sc_hd__xnor2_4 _24218_ (.A(_04460_),
    .B(_04510_),
    .Y(_04511_));
 sky130_fd_sc_hd__nor2_2 _24219_ (.A(_04309_),
    .B(_04306_),
    .Y(_04512_));
 sky130_fd_sc_hd__nand3_1 _24220_ (.A(_04313_),
    .B(_04335_),
    .C(_04512_),
    .Y(_04513_));
 sky130_fd_sc_hd__inv_1 _24221_ (.A(_04313_),
    .Y(_04514_));
 sky130_fd_sc_hd__and2_0 _24222_ (.A(_04309_),
    .B(_04306_),
    .X(_04515_));
 sky130_fd_sc_hd__nand3_1 _24223_ (.A(_04514_),
    .B(_04334_),
    .C(_04515_),
    .Y(_04516_));
 sky130_fd_sc_hd__nand2_1 _24224_ (.A(_04309_),
    .B(_04306_),
    .Y(_04517_));
 sky130_fd_sc_hd__a21oi_1 _24225_ (.A1(_04313_),
    .A2(_04517_),
    .B1(_04512_),
    .Y(_04518_));
 sky130_fd_sc_hd__a22o_1 _24226_ (.A1(_04514_),
    .A2(_04515_),
    .B1(_04518_),
    .B2(_04334_),
    .X(_04519_));
 sky130_fd_sc_hd__nand2_1 _24227_ (.A(_04313_),
    .B(_04512_),
    .Y(_04520_));
 sky130_fd_sc_hd__o21ai_0 _24228_ (.A1(_04334_),
    .A2(_04518_),
    .B1(_04520_),
    .Y(_04521_));
 sky130_fd_sc_hd__mux2i_1 _24229_ (.A0(_04519_),
    .A1(_04521_),
    .S(_04328_),
    .Y(_04522_));
 sky130_fd_sc_hd__and3_1 _24230_ (.A(_04513_),
    .B(_04516_),
    .C(_04522_),
    .X(_04523_));
 sky130_fd_sc_hd__xor2_4 _24231_ (.A(_04511_),
    .B(_04523_),
    .X(_04524_));
 sky130_fd_sc_hd__nand2b_1 _24232_ (.A_N(_04421_),
    .B(_04524_),
    .Y(_04525_));
 sky130_fd_sc_hd__nor2b_1 _24233_ (.A(_04524_),
    .B_N(_04421_),
    .Y(_04526_));
 sky130_fd_sc_hd__inv_1 _24234_ (.A(_04526_),
    .Y(_04527_));
 sky130_fd_sc_hd__nand2_1 _24235_ (.A(_04525_),
    .B(_04527_),
    .Y(_04528_));
 sky130_fd_sc_hd__xor2_1 _24236_ (.A(_04413_),
    .B(_04528_),
    .X(_04529_));
 sky130_fd_sc_hd__nand2_2 _24237_ (.A(_02169_),
    .B(_04529_),
    .Y(_04530_));
 sky130_fd_sc_hd__or2_0 _24238_ (.A(_02169_),
    .B(_02539_),
    .X(_04531_));
 sky130_fd_sc_hd__a21oi_4 _24239_ (.A1(_04530_),
    .A2(_04531_),
    .B1(net443),
    .Y(_04532_));
 sky130_fd_sc_hd__a21oi_4 _24240_ (.A1(net443),
    .A2(_10343_),
    .B1(_04532_),
    .Y(_04533_));
 sky130_fd_sc_hd__nor3_4 _24241_ (.A(net739),
    .B(_04533_),
    .C(_02646_),
    .Y(_04534_));
 sky130_fd_sc_hd__nor3_4 _24242_ (.A(_04397_),
    .B(_04406_),
    .C(net1262),
    .Y(_04535_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_261 ();
 sky130_fd_sc_hd__nand2_1 _24244_ (.A(_02119_),
    .B(net1270),
    .Y(_04537_));
 sky130_fd_sc_hd__nand2_1 _24245_ (.A(\gen_regfile_ff.register_file_i.rf_reg[152] ),
    .B(_02123_),
    .Y(_04538_));
 sky130_fd_sc_hd__nand2_1 _24246_ (.A(_04537_),
    .B(_04538_),
    .Y(_00537_));
 sky130_fd_sc_hd__nand2_1 _24247_ (.A(_04099_),
    .B(_04230_),
    .Y(_04539_));
 sky130_fd_sc_hd__nor2_1 _24248_ (.A(_04372_),
    .B(_04539_),
    .Y(_04540_));
 sky130_fd_sc_hd__nand2_1 _24249_ (.A(_04101_),
    .B(_04230_),
    .Y(_04541_));
 sky130_fd_sc_hd__a21oi_1 _24250_ (.A1(_04407_),
    .A2(_04541_),
    .B1(_04412_),
    .Y(_04542_));
 sky130_fd_sc_hd__a21o_1 _24251_ (.A1(_03992_),
    .A2(_04540_),
    .B1(_04542_),
    .X(_04543_));
 sky130_fd_sc_hd__a21oi_2 _24252_ (.A1(_04525_),
    .A2(_04543_),
    .B1(_04526_),
    .Y(_04544_));
 sky130_fd_sc_hd__nor2_1 _24253_ (.A(_04511_),
    .B(_04512_),
    .Y(_04545_));
 sky130_fd_sc_hd__a21oi_1 _24254_ (.A1(_04511_),
    .A2(_04517_),
    .B1(_04328_),
    .Y(_04546_));
 sky130_fd_sc_hd__o22ai_2 _24255_ (.A1(_04514_),
    .A2(_04334_),
    .B1(_04545_),
    .B2(_04546_),
    .Y(_04547_));
 sky130_fd_sc_hd__nor2_1 _24256_ (.A(_04328_),
    .B(_04512_),
    .Y(_04548_));
 sky130_fd_sc_hd__o21ai_0 _24257_ (.A1(_04313_),
    .A2(_04335_),
    .B1(_04511_),
    .Y(_04549_));
 sky130_fd_sc_hd__o21ai_1 _24258_ (.A1(_04515_),
    .A2(_04548_),
    .B1(_04549_),
    .Y(_04550_));
 sky130_fd_sc_hd__o311ai_4 _24259_ (.A1(_04313_),
    .A2(_04335_),
    .A3(_04511_),
    .B1(_04547_),
    .C1(_04550_),
    .Y(_04551_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_260 ();
 sky130_fd_sc_hd__xor2_1 _24261_ (.A(_04499_),
    .B(_04508_),
    .X(_04553_));
 sky130_fd_sc_hd__xnor2_1 _24262_ (.A(_04459_),
    .B(_04501_),
    .Y(_04554_));
 sky130_fd_sc_hd__maj3_1 _24263_ (.A(_04423_),
    .B(_04553_),
    .C(_04554_),
    .X(_04555_));
 sky130_fd_sc_hd__inv_1 _24264_ (.A(_04494_),
    .Y(_04556_));
 sky130_fd_sc_hd__xnor2_1 _24265_ (.A(_04497_),
    .B(_04508_),
    .Y(_04557_));
 sky130_fd_sc_hd__maj3_1 _24266_ (.A(_04556_),
    .B(_04489_),
    .C(_04557_),
    .X(_04558_));
 sky130_fd_sc_hd__inv_1 _24267_ (.A(_04497_),
    .Y(_04559_));
 sky130_fd_sc_hd__nor2_1 _24268_ (.A(_03670_),
    .B(_04506_),
    .Y(_04560_));
 sky130_fd_sc_hd__maj3_1 _24269_ (.A(_04272_),
    .B(_04559_),
    .C(_04560_),
    .X(_04561_));
 sky130_fd_sc_hd__a21oi_2 _24270_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[57] ),
    .A2(net311),
    .B1(_03772_),
    .Y(_04562_));
 sky130_fd_sc_hd__a21oi_2 _24271_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[55] ),
    .A2(net311),
    .B1(_03772_),
    .Y(_04563_));
 sky130_fd_sc_hd__o21ai_0 _24272_ (.A1(_04563_),
    .A2(_04437_),
    .B1(_03937_),
    .Y(_04564_));
 sky130_fd_sc_hd__o21ai_0 _24273_ (.A1(_03937_),
    .A2(_04563_),
    .B1(_04564_),
    .Y(_04565_));
 sky130_fd_sc_hd__nand2_1 _24274_ (.A(_03933_),
    .B(_04565_),
    .Y(_04566_));
 sky130_fd_sc_hd__o21ai_0 _24275_ (.A1(_03937_),
    .A2(_04437_),
    .B1(_04566_),
    .Y(_04567_));
 sky130_fd_sc_hd__nand3_1 _24276_ (.A(_03941_),
    .B(_04049_),
    .C(_04437_),
    .Y(_04568_));
 sky130_fd_sc_hd__nor2_1 _24277_ (.A(_04049_),
    .B(_04437_),
    .Y(_04569_));
 sky130_fd_sc_hd__nand2_1 _24278_ (.A(_03933_),
    .B(_04569_),
    .Y(_04570_));
 sky130_fd_sc_hd__a21oi_1 _24279_ (.A1(_04568_),
    .A2(_04570_),
    .B1(_03927_),
    .Y(_04571_));
 sky130_fd_sc_hd__a21oi_1 _24280_ (.A1(_03927_),
    .A2(_04567_),
    .B1(_04571_),
    .Y(_04572_));
 sky130_fd_sc_hd__xnor2_2 _24281_ (.A(_04562_),
    .B(_04572_),
    .Y(_04573_));
 sky130_fd_sc_hd__nand2_1 _24282_ (.A(_03933_),
    .B(_04563_),
    .Y(_04574_));
 sky130_fd_sc_hd__a21oi_1 _24283_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[54] ),
    .A2(net311),
    .B1(_03772_),
    .Y(_04575_));
 sky130_fd_sc_hd__nor2_1 _24284_ (.A(_03937_),
    .B(_04575_),
    .Y(_04576_));
 sky130_fd_sc_hd__a21oi_1 _24285_ (.A1(_04576_),
    .A2(_04437_),
    .B1(_04569_),
    .Y(_04577_));
 sky130_fd_sc_hd__nor3_1 _24286_ (.A(_04061_),
    .B(_04432_),
    .C(_04439_),
    .Y(_04578_));
 sky130_fd_sc_hd__a21oi_1 _24287_ (.A1(_04061_),
    .A2(_04439_),
    .B1(_04578_),
    .Y(_04579_));
 sky130_fd_sc_hd__nor2_1 _24288_ (.A(_03695_),
    .B(_04579_),
    .Y(_04580_));
 sky130_fd_sc_hd__a31oi_1 _24289_ (.A1(_04453_),
    .A2(_04432_),
    .A3(_04439_),
    .B1(_04580_),
    .Y(_04581_));
 sky130_fd_sc_hd__o21ai_0 _24290_ (.A1(_04574_),
    .A2(_04577_),
    .B1(_04581_),
    .Y(_04582_));
 sky130_fd_sc_hd__nand2_1 _24291_ (.A(_03941_),
    .B(_04049_),
    .Y(_04583_));
 sky130_fd_sc_hd__a21oi_1 _24292_ (.A1(_04352_),
    .A2(_04583_),
    .B1(_04563_),
    .Y(_04584_));
 sky130_fd_sc_hd__nor3_1 _24293_ (.A(_03933_),
    .B(_04049_),
    .C(_04437_),
    .Y(_04585_));
 sky130_fd_sc_hd__a21oi_1 _24294_ (.A1(_04437_),
    .A2(_04584_),
    .B1(_04585_),
    .Y(_04586_));
 sky130_fd_sc_hd__nor2_1 _24295_ (.A(_03927_),
    .B(_04586_),
    .Y(_04587_));
 sky130_fd_sc_hd__a21oi_2 _24296_ (.A1(_03927_),
    .A2(_04582_),
    .B1(_04587_),
    .Y(_04588_));
 sky130_fd_sc_hd__xnor3_1 _24297_ (.A(_04561_),
    .B(_04573_),
    .C(_04588_),
    .X(_04589_));
 sky130_fd_sc_hd__xnor2_1 _24298_ (.A(_04558_),
    .B(_04589_),
    .Y(_04590_));
 sky130_fd_sc_hd__nand2_1 _24299_ (.A(_02889_),
    .B(_03161_),
    .Y(_04591_));
 sky130_fd_sc_hd__nand2_1 _24300_ (.A(_03142_),
    .B(_03376_),
    .Y(_04592_));
 sky130_fd_sc_hd__nand2_1 _24301_ (.A(_03407_),
    .B(_03310_),
    .Y(_04593_));
 sky130_fd_sc_hd__xor2_1 _24302_ (.A(_04592_),
    .B(_04593_),
    .X(_04594_));
 sky130_fd_sc_hd__xor2_2 _24303_ (.A(_04591_),
    .B(_04594_),
    .X(_04595_));
 sky130_fd_sc_hd__nor2_1 _24304_ (.A(net899),
    .B(_03100_),
    .Y(_04596_));
 sky130_fd_sc_hd__nor2_1 _24305_ (.A(_02936_),
    .B(_03119_),
    .Y(_04597_));
 sky130_fd_sc_hd__nor2_1 _24306_ (.A(_03097_),
    .B(net1263),
    .Y(_04598_));
 sky130_fd_sc_hd__xnor2_1 _24307_ (.A(_04597_),
    .B(_04598_),
    .Y(_04599_));
 sky130_fd_sc_hd__xor2_1 _24308_ (.A(_04596_),
    .B(_04599_),
    .X(_04600_));
 sky130_fd_sc_hd__a22o_1 _24309_ (.A1(net1004),
    .A2(_03376_),
    .B1(_04468_),
    .B2(_04469_),
    .X(_04601_));
 sky130_fd_sc_hd__o21ai_2 _24310_ (.A1(_04468_),
    .A2(_04469_),
    .B1(_04601_),
    .Y(_04602_));
 sky130_fd_sc_hd__xnor2_1 _24311_ (.A(_04600_),
    .B(_04602_),
    .Y(_04603_));
 sky130_fd_sc_hd__xnor2_2 _24312_ (.A(_04595_),
    .B(_04603_),
    .Y(_04604_));
 sky130_fd_sc_hd__nand3_1 _24313_ (.A(net1173),
    .B(_02727_),
    .C(_03274_),
    .Y(_04605_));
 sky130_fd_sc_hd__o31ai_1 _24314_ (.A1(net1173),
    .A2(_02727_),
    .A3(_03512_),
    .B1(_04605_),
    .Y(_04606_));
 sky130_fd_sc_hd__nand2b_2 _24315_ (.A_N(net1173),
    .B(_02727_),
    .Y(_04607_));
 sky130_fd_sc_hd__o21ai_0 _24316_ (.A1(net1158),
    .A2(_04020_),
    .B1(net1173),
    .Y(_04608_));
 sky130_fd_sc_hd__nand2_1 _24317_ (.A(_04607_),
    .B(_04608_),
    .Y(_04609_));
 sky130_fd_sc_hd__a32o_1 _24318_ (.A1(_02727_),
    .A2(_03274_),
    .A3(_03512_),
    .B1(_04479_),
    .B2(_04609_),
    .X(_04610_));
 sky130_fd_sc_hd__a21oi_1 _24319_ (.A1(net1161),
    .A2(_04606_),
    .B1(_04610_),
    .Y(_04611_));
 sky130_fd_sc_hd__nand2_1 _24320_ (.A(_04461_),
    .B(_04462_),
    .Y(_04612_));
 sky130_fd_sc_hd__nor2_1 _24321_ (.A(_04461_),
    .B(_04462_),
    .Y(_04613_));
 sky130_fd_sc_hd__a21oi_1 _24322_ (.A1(_04463_),
    .A2(_04612_),
    .B1(_04613_),
    .Y(_04614_));
 sky130_fd_sc_hd__o21ai_0 _24323_ (.A1(net1173),
    .A2(_04020_),
    .B1(_04477_),
    .Y(_04615_));
 sky130_fd_sc_hd__nor3_1 _24324_ (.A(net1173),
    .B(_04020_),
    .C(_04477_),
    .Y(_04616_));
 sky130_fd_sc_hd__a21oi_1 _24325_ (.A1(_04479_),
    .A2(_04615_),
    .B1(_04616_),
    .Y(_04617_));
 sky130_fd_sc_hd__xnor2_1 _24326_ (.A(_04614_),
    .B(_04617_),
    .Y(_04618_));
 sky130_fd_sc_hd__xnor2_1 _24327_ (.A(_04611_),
    .B(_04618_),
    .Y(_04619_));
 sky130_fd_sc_hd__nand2_1 _24328_ (.A(_04465_),
    .B(_04472_),
    .Y(_04620_));
 sky130_fd_sc_hd__nor2_1 _24329_ (.A(_04465_),
    .B(_04472_),
    .Y(_04621_));
 sky130_fd_sc_hd__a21o_1 _24330_ (.A1(_04467_),
    .A2(_04620_),
    .B1(_04621_),
    .X(_04622_));
 sky130_fd_sc_hd__nor2_1 _24331_ (.A(_04619_),
    .B(_04622_),
    .Y(_04623_));
 sky130_fd_sc_hd__nand2_1 _24332_ (.A(_04619_),
    .B(_04622_),
    .Y(_04624_));
 sky130_fd_sc_hd__nor2b_1 _24333_ (.A(_04623_),
    .B_N(_04624_),
    .Y(_04625_));
 sky130_fd_sc_hd__xnor2_2 _24334_ (.A(_04604_),
    .B(_04625_),
    .Y(_04626_));
 sky130_fd_sc_hd__inv_1 _24335_ (.A(_04486_),
    .Y(_04627_));
 sky130_fd_sc_hd__a21oi_2 _24336_ (.A1(_04474_),
    .A2(_04627_),
    .B1(_04487_),
    .Y(_04628_));
 sky130_fd_sc_hd__maj3_2 _24337_ (.A(_04482_),
    .B(_04481_),
    .C(_04483_),
    .X(_04629_));
 sky130_fd_sc_hd__xor2_1 _24338_ (.A(_04628_),
    .B(_04629_),
    .X(_04630_));
 sky130_fd_sc_hd__xnor2_1 _24339_ (.A(_04626_),
    .B(_04630_),
    .Y(_04631_));
 sky130_fd_sc_hd__xor2_1 _24340_ (.A(_04509_),
    .B(_04631_),
    .X(_04632_));
 sky130_fd_sc_hd__xnor2_1 _24341_ (.A(_04590_),
    .B(_04632_),
    .Y(_04633_));
 sky130_fd_sc_hd__xnor2_1 _24342_ (.A(_04441_),
    .B(_04501_),
    .Y(_04634_));
 sky130_fd_sc_hd__nand2_1 _24343_ (.A(_04457_),
    .B(_04634_),
    .Y(_04635_));
 sky130_fd_sc_hd__nand2_1 _24344_ (.A(_04445_),
    .B(_04635_),
    .Y(_04636_));
 sky130_fd_sc_hd__o21ai_1 _24345_ (.A1(_04457_),
    .A2(_04634_),
    .B1(_04636_),
    .Y(_04637_));
 sky130_fd_sc_hd__xnor2_1 _24346_ (.A(_04633_),
    .B(_04637_),
    .Y(_04638_));
 sky130_fd_sc_hd__xnor2_1 _24347_ (.A(_04555_),
    .B(_04638_),
    .Y(_04639_));
 sky130_fd_sc_hd__or2_0 _24348_ (.A(_04551_),
    .B(_04639_),
    .X(_04640_));
 sky130_fd_sc_hd__nand2_1 _24349_ (.A(_04551_),
    .B(_04639_),
    .Y(_04641_));
 sky130_fd_sc_hd__nand2_1 _24350_ (.A(_04640_),
    .B(_04641_),
    .Y(_04642_));
 sky130_fd_sc_hd__xor2_1 _24351_ (.A(_04642_),
    .B(_04544_),
    .X(_04643_));
 sky130_fd_sc_hd__nand2_1 _24352_ (.A(_02169_),
    .B(_04643_),
    .Y(_04644_));
 sky130_fd_sc_hd__o21ai_2 _24353_ (.A1(_02169_),
    .A2(_02641_),
    .B1(_04644_),
    .Y(_04645_));
 sky130_fd_sc_hd__mux2i_4 _24354_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[57] ),
    .A1(_04645_),
    .S(_08100_),
    .Y(_04646_));
 sky130_fd_sc_hd__and2_0 _24355_ (.A(_02646_),
    .B(_03478_),
    .X(_04647_));
 sky130_fd_sc_hd__mux4_1 _24356_ (.A0(net44),
    .A1(net58),
    .A2(net38),
    .A3(net35),
    .S0(\load_store_unit_i.rdata_offset_q[1] ),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .X(_04648_));
 sky130_fd_sc_hd__nand2_1 _24357_ (.A(_01674_),
    .B(_04648_),
    .Y(_04649_));
 sky130_fd_sc_hd__nand2_1 _24358_ (.A(_04647_),
    .B(_04649_),
    .Y(_04650_));
 sky130_fd_sc_hd__nor2_1 _24359_ (.A(_01773_),
    .B(_02272_),
    .Y(_04651_));
 sky130_fd_sc_hd__a21oi_1 _24360_ (.A1(_01773_),
    .A2(_02276_),
    .B1(_04651_),
    .Y(_04652_));
 sky130_fd_sc_hd__nor3_1 _24361_ (.A(_10303_),
    .B(_10335_),
    .C(_01898_),
    .Y(_04653_));
 sky130_fd_sc_hd__a21oi_1 _24362_ (.A1(_10335_),
    .A2(_01896_),
    .B1(_04653_),
    .Y(_04654_));
 sky130_fd_sc_hd__o21ai_0 _24363_ (.A1(_10335_),
    .A2(_01903_),
    .B1(_10303_),
    .Y(_04655_));
 sky130_fd_sc_hd__o21ai_0 _24364_ (.A1(_01893_),
    .A2(_04654_),
    .B1(_04655_),
    .Y(_04656_));
 sky130_fd_sc_hd__nand2_1 _24365_ (.A(_08290_),
    .B(_04656_),
    .Y(_04657_));
 sky130_fd_sc_hd__a21oi_1 _24366_ (.A1(_01734_),
    .A2(_04652_),
    .B1(_04657_),
    .Y(_04658_));
 sky130_fd_sc_hd__o2111ai_4 _24367_ (.A1(net684),
    .A2(_01889_),
    .B1(_04658_),
    .C1(_11704_),
    .D1(net1484),
    .Y(_04659_));
 sky130_fd_sc_hd__nand2_1 _24368_ (.A(_04650_),
    .B(_04659_),
    .Y(_04660_));
 sky130_fd_sc_hd__a31oi_4 _24369_ (.A1(_04646_),
    .A2(net265),
    .A3(net1101),
    .B1(_04660_),
    .Y(_04661_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_259 ();
 sky130_fd_sc_hd__nand2_2 _24371_ (.A(net1564),
    .B(_02119_),
    .Y(_04663_));
 sky130_fd_sc_hd__nand2_1 _24372_ (.A(\gen_regfile_ff.register_file_i.rf_reg[153] ),
    .B(_02123_),
    .Y(_04664_));
 sky130_fd_sc_hd__nand2_1 _24373_ (.A(_04663_),
    .B(_04664_),
    .Y(_00538_));
 sky130_fd_sc_hd__o21a_1 _24374_ (.A1(_04526_),
    .A2(_04413_),
    .B1(_04525_),
    .X(_04665_));
 sky130_fd_sc_hd__maj3_2 _24375_ (.A(_04665_),
    .B(_04639_),
    .C(_04551_),
    .X(_04666_));
 sky130_fd_sc_hd__inv_1 _24376_ (.A(_04633_),
    .Y(_04667_));
 sky130_fd_sc_hd__nand2_1 _24377_ (.A(_04667_),
    .B(_04637_),
    .Y(_04668_));
 sky130_fd_sc_hd__nor2_1 _24378_ (.A(_04667_),
    .B(_04637_),
    .Y(_04669_));
 sky130_fd_sc_hd__a21oi_2 _24379_ (.A1(_04555_),
    .A2(_04668_),
    .B1(_04669_),
    .Y(_04670_));
 sky130_fd_sc_hd__xnor2_1 _24380_ (.A(_04508_),
    .B(_04631_),
    .Y(_04671_));
 sky130_fd_sc_hd__nand3_4 _24381_ (.A(_03428_),
    .B(_03515_),
    .C(_03936_),
    .Y(_04672_));
 sky130_fd_sc_hd__nand2_2 _24382_ (.A(_03927_),
    .B(_04049_),
    .Y(_04673_));
 sky130_fd_sc_hd__nand2_8 _24383_ (.A(_04672_),
    .B(_04673_),
    .Y(_04674_));
 sky130_fd_sc_hd__xor2_1 _24384_ (.A(_04674_),
    .B(_04589_),
    .X(_04675_));
 sky130_fd_sc_hd__maj3_1 _24385_ (.A(_04558_),
    .B(_04671_),
    .C(_04675_),
    .X(_04676_));
 sky130_fd_sc_hd__nor2_1 _24386_ (.A(_03941_),
    .B(_04049_),
    .Y(_04677_));
 sky130_fd_sc_hd__a21o_1 _24387_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[57] ),
    .A2(net311),
    .B1(_03772_),
    .X(_04678_));
 sky130_fd_sc_hd__nor2_1 _24388_ (.A(_04437_),
    .B(_04678_),
    .Y(_04679_));
 sky130_fd_sc_hd__nor2_1 _24389_ (.A(_04049_),
    .B(_04562_),
    .Y(_04680_));
 sky130_fd_sc_hd__a21oi_1 _24390_ (.A1(_04049_),
    .A2(_04679_),
    .B1(_04680_),
    .Y(_04681_));
 sky130_fd_sc_hd__nor2_1 _24391_ (.A(_03933_),
    .B(_04681_),
    .Y(_04682_));
 sky130_fd_sc_hd__a21oi_1 _24392_ (.A1(_04677_),
    .A2(_04679_),
    .B1(_04682_),
    .Y(_04683_));
 sky130_fd_sc_hd__nor4_1 _24393_ (.A(_04049_),
    .B(_04563_),
    .C(_04437_),
    .D(_04678_),
    .Y(_04684_));
 sky130_fd_sc_hd__nor3_1 _24394_ (.A(_03937_),
    .B(_04563_),
    .C(_04678_),
    .Y(_04685_));
 sky130_fd_sc_hd__o21ai_0 _24395_ (.A1(_04680_),
    .A2(_04685_),
    .B1(_04437_),
    .Y(_04686_));
 sky130_fd_sc_hd__nand3_1 _24396_ (.A(_04049_),
    .B(_04437_),
    .C(_04678_),
    .Y(_04687_));
 sky130_fd_sc_hd__o21ai_0 _24397_ (.A1(_04049_),
    .A2(_04678_),
    .B1(_04687_),
    .Y(_04688_));
 sky130_fd_sc_hd__nor2_1 _24398_ (.A(_03933_),
    .B(_04688_),
    .Y(_04689_));
 sky130_fd_sc_hd__a21oi_1 _24399_ (.A1(_03933_),
    .A2(_04686_),
    .B1(_04689_),
    .Y(_04690_));
 sky130_fd_sc_hd__o21ai_0 _24400_ (.A1(_04684_),
    .A2(_04690_),
    .B1(_03927_),
    .Y(_04691_));
 sky130_fd_sc_hd__o21ai_2 _24401_ (.A1(_03927_),
    .A2(_04683_),
    .B1(_04691_),
    .Y(_04692_));
 sky130_fd_sc_hd__a21o_1 _24402_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[58] ),
    .A2(net311),
    .B1(_03772_),
    .X(_04693_));
 sky130_fd_sc_hd__o21ai_0 _24403_ (.A1(_04437_),
    .A2(_04562_),
    .B1(_03937_),
    .Y(_04694_));
 sky130_fd_sc_hd__o21ai_0 _24404_ (.A1(_03937_),
    .A2(_04437_),
    .B1(_04694_),
    .Y(_04695_));
 sky130_fd_sc_hd__nand2_1 _24405_ (.A(_03933_),
    .B(_04695_),
    .Y(_04696_));
 sky130_fd_sc_hd__o21ai_0 _24406_ (.A1(_03937_),
    .A2(_04562_),
    .B1(_04696_),
    .Y(_04697_));
 sky130_fd_sc_hd__nand3_1 _24407_ (.A(_03941_),
    .B(_04049_),
    .C(_04562_),
    .Y(_04698_));
 sky130_fd_sc_hd__nand2_1 _24408_ (.A(_03933_),
    .B(_04680_),
    .Y(_04699_));
 sky130_fd_sc_hd__a21oi_1 _24409_ (.A1(_04698_),
    .A2(_04699_),
    .B1(_03927_),
    .Y(_04700_));
 sky130_fd_sc_hd__a21oi_1 _24410_ (.A1(_03927_),
    .A2(_04697_),
    .B1(_04700_),
    .Y(_04701_));
 sky130_fd_sc_hd__xor2_2 _24411_ (.A(_04693_),
    .B(_04701_),
    .X(_04702_));
 sky130_fd_sc_hd__maj3_1 _24412_ (.A(_04272_),
    .B(_04560_),
    .C(_04629_),
    .X(_04703_));
 sky130_fd_sc_hd__xnor2_1 _24413_ (.A(_04702_),
    .B(_04703_),
    .Y(_04704_));
 sky130_fd_sc_hd__xnor2_1 _24414_ (.A(_04692_),
    .B(_04704_),
    .Y(_04705_));
 sky130_fd_sc_hd__xnor2_1 _24415_ (.A(_04508_),
    .B(_04629_),
    .Y(_04706_));
 sky130_fd_sc_hd__maj3_1 _24416_ (.A(_04628_),
    .B(_04626_),
    .C(_04706_),
    .X(_04707_));
 sky130_fd_sc_hd__a21oi_2 _24417_ (.A1(_04604_),
    .A2(_04624_),
    .B1(_04623_),
    .Y(_04708_));
 sky130_fd_sc_hd__nand2_1 _24418_ (.A(net1414),
    .B(_03376_),
    .Y(_04709_));
 sky130_fd_sc_hd__nand2_1 _24419_ (.A(_02889_),
    .B(_03310_),
    .Y(_04710_));
 sky130_fd_sc_hd__nand2_1 _24420_ (.A(_02897_),
    .B(_03161_),
    .Y(_04711_));
 sky130_fd_sc_hd__xor2_1 _24421_ (.A(_04710_),
    .B(_04711_),
    .X(_04712_));
 sky130_fd_sc_hd__xnor2_1 _24422_ (.A(_04709_),
    .B(_04712_),
    .Y(_04713_));
 sky130_fd_sc_hd__inv_1 _24423_ (.A(_04713_),
    .Y(_04714_));
 sky130_fd_sc_hd__maj3_1 _24424_ (.A(_04591_),
    .B(_04592_),
    .C(_04593_),
    .X(_04715_));
 sky130_fd_sc_hd__nor2_1 _24425_ (.A(net899),
    .B(_03119_),
    .Y(_04716_));
 sky130_fd_sc_hd__nor2_1 _24426_ (.A(net1264),
    .B(_03100_),
    .Y(_04717_));
 sky130_fd_sc_hd__nor2_1 _24427_ (.A(_02936_),
    .B(_04020_),
    .Y(_04718_));
 sky130_fd_sc_hd__xnor2_1 _24428_ (.A(_04717_),
    .B(_04718_),
    .Y(_04719_));
 sky130_fd_sc_hd__xor2_1 _24429_ (.A(_04716_),
    .B(_04719_),
    .X(_04720_));
 sky130_fd_sc_hd__xnor2_1 _24430_ (.A(_04715_),
    .B(_04720_),
    .Y(_04721_));
 sky130_fd_sc_hd__xnor2_1 _24431_ (.A(_04714_),
    .B(_04721_),
    .Y(_04722_));
 sky130_fd_sc_hd__maj3_1 _24432_ (.A(_04600_),
    .B(_04595_),
    .C(_04602_),
    .X(_04723_));
 sky130_fd_sc_hd__maj3_1 _24433_ (.A(_04596_),
    .B(_04597_),
    .C(_04598_),
    .X(_04724_));
 sky130_fd_sc_hd__nand3_1 _24434_ (.A(net1161),
    .B(net1173),
    .C(net1158),
    .Y(_04725_));
 sky130_fd_sc_hd__o21ai_1 _24435_ (.A1(net1161),
    .A2(_04607_),
    .B1(_04725_),
    .Y(_04726_));
 sky130_fd_sc_hd__nor2_2 _24436_ (.A(_03512_),
    .B(_04726_),
    .Y(_04727_));
 sky130_fd_sc_hd__xnor2_1 _24437_ (.A(_04724_),
    .B(_04727_),
    .Y(_04728_));
 sky130_fd_sc_hd__xor2_1 _24438_ (.A(_04723_),
    .B(_04728_),
    .X(_04729_));
 sky130_fd_sc_hd__xnor2_2 _24439_ (.A(_04722_),
    .B(_04729_),
    .Y(_04730_));
 sky130_fd_sc_hd__inv_1 _24440_ (.A(_04611_),
    .Y(_04731_));
 sky130_fd_sc_hd__inv_1 _24441_ (.A(_04617_),
    .Y(_04732_));
 sky130_fd_sc_hd__maj3_2 _24442_ (.A(_04614_),
    .B(_04731_),
    .C(_04732_),
    .X(_04733_));
 sky130_fd_sc_hd__xnor2_1 _24443_ (.A(_04730_),
    .B(_04733_),
    .Y(_04734_));
 sky130_fd_sc_hd__xnor2_1 _24444_ (.A(_04708_),
    .B(_04734_),
    .Y(_04735_));
 sky130_fd_sc_hd__xor2_1 _24445_ (.A(_04509_),
    .B(_04735_),
    .X(_04736_));
 sky130_fd_sc_hd__xnor2_1 _24446_ (.A(_04707_),
    .B(_04736_),
    .Y(_04737_));
 sky130_fd_sc_hd__xnor2_1 _24447_ (.A(_04705_),
    .B(_04737_),
    .Y(_04738_));
 sky130_fd_sc_hd__xnor2_1 _24448_ (.A(_04674_),
    .B(_04573_),
    .Y(_04739_));
 sky130_fd_sc_hd__nand2_1 _24449_ (.A(_04561_),
    .B(_04739_),
    .Y(_04740_));
 sky130_fd_sc_hd__nor2_1 _24450_ (.A(_04561_),
    .B(_04739_),
    .Y(_04741_));
 sky130_fd_sc_hd__a21oi_1 _24451_ (.A1(_04588_),
    .A2(_04740_),
    .B1(_04741_),
    .Y(_04742_));
 sky130_fd_sc_hd__xnor2_1 _24452_ (.A(_04738_),
    .B(_04742_),
    .Y(_04743_));
 sky130_fd_sc_hd__xnor2_2 _24453_ (.A(_04676_),
    .B(_04743_),
    .Y(_04744_));
 sky130_fd_sc_hd__xnor2_1 _24454_ (.A(_04670_),
    .B(_04744_),
    .Y(_04745_));
 sky130_fd_sc_hd__xnor2_2 _24455_ (.A(_04666_),
    .B(_04745_),
    .Y(_04746_));
 sky130_fd_sc_hd__mux2_4 _24456_ (.A0(_02751_),
    .A1(_04746_),
    .S(_02169_),
    .X(_04747_));
 sky130_fd_sc_hd__mux2i_4 _24457_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[58] ),
    .A1(_04747_),
    .S(_08100_),
    .Y(_04748_));
 sky130_fd_sc_hd__mux4_1 _24458_ (.A0(net45),
    .A1(net28),
    .A2(net49),
    .A3(net36),
    .S0(\load_store_unit_i.rdata_offset_q[1] ),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .X(_04749_));
 sky130_fd_sc_hd__nand2_1 _24459_ (.A(_01674_),
    .B(_04749_),
    .Y(_04750_));
 sky130_fd_sc_hd__nand2_1 _24460_ (.A(_04647_),
    .B(_04750_),
    .Y(_04751_));
 sky130_fd_sc_hd__nand2_1 _24461_ (.A(net295),
    .B(_02214_),
    .Y(_04752_));
 sky130_fd_sc_hd__o21ai_0 _24462_ (.A1(net295),
    .A2(_02222_),
    .B1(_04752_),
    .Y(_04753_));
 sky130_fd_sc_hd__nand2_1 _24463_ (.A(_10468_),
    .B(_02233_),
    .Y(_04754_));
 sky130_fd_sc_hd__nor2_1 _24464_ (.A(_10440_),
    .B(_01898_),
    .Y(_04755_));
 sky130_fd_sc_hd__nor2_1 _24465_ (.A(_10468_),
    .B(_01902_),
    .Y(_04756_));
 sky130_fd_sc_hd__a21oi_1 _24466_ (.A1(_10468_),
    .A2(_04755_),
    .B1(_04756_),
    .Y(_04757_));
 sky130_fd_sc_hd__nor2_1 _24467_ (.A(_01893_),
    .B(_04757_),
    .Y(_04758_));
 sky130_fd_sc_hd__a21oi_1 _24468_ (.A1(_10440_),
    .A2(_04754_),
    .B1(_04758_),
    .Y(_04759_));
 sky130_fd_sc_hd__a221oi_2 _24469_ (.A1(net167),
    .A2(_01929_),
    .B1(_04753_),
    .B2(_01734_),
    .C1(_04759_),
    .Y(_04760_));
 sky130_fd_sc_hd__nand4_4 _24470_ (.A(_08290_),
    .B(_11724_),
    .C(net1485),
    .D(_04760_),
    .Y(_04761_));
 sky130_fd_sc_hd__nand2_1 _24471_ (.A(_04751_),
    .B(_04761_),
    .Y(_04762_));
 sky130_fd_sc_hd__a31oi_4 _24472_ (.A1(net1102),
    .A2(net265),
    .A3(_04748_),
    .B1(_04762_),
    .Y(_04763_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_258 ();
 sky130_fd_sc_hd__nand2_1 _24474_ (.A(_02119_),
    .B(net1515),
    .Y(_04765_));
 sky130_fd_sc_hd__nand2_1 _24475_ (.A(\gen_regfile_ff.register_file_i.rf_reg[154] ),
    .B(_02123_),
    .Y(_04766_));
 sky130_fd_sc_hd__nand2_1 _24476_ (.A(_04765_),
    .B(_04766_),
    .Y(_00539_));
 sky130_fd_sc_hd__o211a_1 _24477_ (.A1(_04539_),
    .A2(_04373_),
    .B1(_04524_),
    .C1(_04407_),
    .X(_04767_));
 sky130_fd_sc_hd__nor3_1 _24478_ (.A(_04372_),
    .B(_04524_),
    .C(_04539_),
    .Y(_04768_));
 sky130_fd_sc_hd__a211oi_1 _24479_ (.A1(_04407_),
    .A2(_04541_),
    .B1(_04524_),
    .C1(_04412_),
    .Y(_04769_));
 sky130_fd_sc_hd__a21boi_0 _24480_ (.A1(_04412_),
    .A2(_04524_),
    .B1_N(_04421_),
    .Y(_04770_));
 sky130_fd_sc_hd__a211oi_2 _24481_ (.A1(_03992_),
    .A2(_04768_),
    .B1(_04769_),
    .C1(_04770_),
    .Y(_04771_));
 sky130_fd_sc_hd__or2_0 _24482_ (.A(_04670_),
    .B(_04744_),
    .X(_04772_));
 sky130_fd_sc_hd__nand2_1 _24483_ (.A(_04640_),
    .B(_04772_),
    .Y(_04773_));
 sky130_fd_sc_hd__a22o_1 _24484_ (.A1(_04551_),
    .A2(_04639_),
    .B1(_04670_),
    .B2(_04744_),
    .X(_04774_));
 sky130_fd_sc_hd__nand2_2 _24485_ (.A(_04772_),
    .B(_04774_),
    .Y(_04775_));
 sky130_fd_sc_hd__o31ai_4 _24486_ (.A1(_04767_),
    .A2(_04771_),
    .A3(_04773_),
    .B1(_04775_),
    .Y(_04776_));
 sky130_fd_sc_hd__xnor2_1 _24487_ (.A(_04508_),
    .B(_04735_),
    .Y(_04777_));
 sky130_fd_sc_hd__xnor2_1 _24488_ (.A(_04674_),
    .B(_04705_),
    .Y(_04778_));
 sky130_fd_sc_hd__maj3_1 _24489_ (.A(_04707_),
    .B(_04777_),
    .C(_04778_),
    .X(_04779_));
 sky130_fd_sc_hd__xnor2_1 _24490_ (.A(_04508_),
    .B(_04733_),
    .Y(_04780_));
 sky130_fd_sc_hd__maj3_1 _24491_ (.A(_04708_),
    .B(_04730_),
    .C(_04780_),
    .X(_04781_));
 sky130_fd_sc_hd__xor2_1 _24492_ (.A(_04509_),
    .B(_04781_),
    .X(_04782_));
 sky130_fd_sc_hd__maj3_1 _24493_ (.A(_04722_),
    .B(_04723_),
    .C(_04728_),
    .X(_04783_));
 sky130_fd_sc_hd__nor2_1 _24494_ (.A(net1265),
    .B(_03119_),
    .Y(_04784_));
 sky130_fd_sc_hd__nor2_1 _24495_ (.A(net899),
    .B(_04020_),
    .Y(_04785_));
 sky130_fd_sc_hd__nor2_1 _24496_ (.A(_02936_),
    .B(_03512_),
    .Y(_04786_));
 sky130_fd_sc_hd__xnor2_1 _24497_ (.A(_04785_),
    .B(_04786_),
    .Y(_04787_));
 sky130_fd_sc_hd__xor2_1 _24498_ (.A(_04784_),
    .B(_04787_),
    .X(_04788_));
 sky130_fd_sc_hd__nor2_1 _24499_ (.A(_03097_),
    .B(_03373_),
    .Y(_04789_));
 sky130_fd_sc_hd__nor2_1 _24500_ (.A(_03100_),
    .B(_03313_),
    .Y(_04790_));
 sky130_fd_sc_hd__nor2_1 _24501_ (.A(_02889_),
    .B(_03370_),
    .Y(_04791_));
 sky130_fd_sc_hd__xor2_1 _24502_ (.A(_04790_),
    .B(_04791_),
    .X(_04792_));
 sky130_fd_sc_hd__xnor2_2 _24503_ (.A(_04789_),
    .B(_04792_),
    .Y(_04793_));
 sky130_fd_sc_hd__maj3_1 _24504_ (.A(_04710_),
    .B(_04711_),
    .C(_04709_),
    .X(_04794_));
 sky130_fd_sc_hd__xnor2_1 _24505_ (.A(_04793_),
    .B(_04794_),
    .Y(_04795_));
 sky130_fd_sc_hd__xnor2_1 _24506_ (.A(_04788_),
    .B(_04795_),
    .Y(_04796_));
 sky130_fd_sc_hd__maj3_1 _24507_ (.A(_04714_),
    .B(_04715_),
    .C(_04720_),
    .X(_04797_));
 sky130_fd_sc_hd__maj3_1 _24508_ (.A(_04716_),
    .B(_04717_),
    .C(_04718_),
    .X(_04798_));
 sky130_fd_sc_hd__xnor2_1 _24509_ (.A(_04727_),
    .B(_04798_),
    .Y(_04799_));
 sky130_fd_sc_hd__xnor2_1 _24510_ (.A(_04797_),
    .B(_04799_),
    .Y(_04800_));
 sky130_fd_sc_hd__xnor2_2 _24511_ (.A(_04796_),
    .B(_04800_),
    .Y(_04801_));
 sky130_fd_sc_hd__nand2_1 _24512_ (.A(net1173),
    .B(net1158),
    .Y(_04802_));
 sky130_fd_sc_hd__inv_1 _24513_ (.A(_04724_),
    .Y(_04803_));
 sky130_fd_sc_hd__a21oi_1 _24514_ (.A1(_04607_),
    .A2(_04803_),
    .B1(net1161),
    .Y(_04804_));
 sky130_fd_sc_hd__a21oi_1 _24515_ (.A1(_04724_),
    .A2(_04802_),
    .B1(_04804_),
    .Y(_04805_));
 sky130_fd_sc_hd__nor2_1 _24516_ (.A(_03512_),
    .B(_04805_),
    .Y(_04806_));
 sky130_fd_sc_hd__xnor2_1 _24517_ (.A(_04801_),
    .B(_04806_),
    .Y(_04807_));
 sky130_fd_sc_hd__xor2_1 _24518_ (.A(_04783_),
    .B(_04807_),
    .X(_04808_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_257 ();
 sky130_fd_sc_hd__a21oi_4 _24520_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[58] ),
    .A2(_03509_),
    .B1(_03684_),
    .Y(_04810_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_256 ();
 sky130_fd_sc_hd__nand3_1 _24522_ (.A(_03698_),
    .B(_04182_),
    .C(_04810_),
    .Y(_04812_));
 sky130_fd_sc_hd__nor2_1 _24523_ (.A(_04182_),
    .B(_04810_),
    .Y(_04813_));
 sky130_fd_sc_hd__nand2_1 _24524_ (.A(_03695_),
    .B(_04813_),
    .Y(_04814_));
 sky130_fd_sc_hd__a21o_1 _24525_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[57] ),
    .A2(_03509_),
    .B1(_03684_),
    .X(_04815_));
 sky130_fd_sc_hd__nand2_1 _24526_ (.A(_04182_),
    .B(_04815_),
    .Y(_04816_));
 sky130_fd_sc_hd__a21oi_1 _24527_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[57] ),
    .A2(_03509_),
    .B1(_03684_),
    .Y(_04817_));
 sky130_fd_sc_hd__o21ai_0 _24528_ (.A1(_04817_),
    .A2(_04810_),
    .B1(_04061_),
    .Y(_04818_));
 sky130_fd_sc_hd__a21oi_1 _24529_ (.A1(_04816_),
    .A2(_04818_),
    .B1(_03698_),
    .Y(_04819_));
 sky130_fd_sc_hd__nor2_1 _24530_ (.A(_04061_),
    .B(_04810_),
    .Y(_04820_));
 sky130_fd_sc_hd__nor3_1 _24531_ (.A(_03690_),
    .B(_04819_),
    .C(_04820_),
    .Y(_04821_));
 sky130_fd_sc_hd__a31oi_2 _24532_ (.A1(_03690_),
    .A2(_04812_),
    .A3(_04814_),
    .B1(_04821_),
    .Y(_04822_));
 sky130_fd_sc_hd__a21o_1 _24533_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[59] ),
    .A2(_03509_),
    .B1(_03684_),
    .X(_04823_));
 sky130_fd_sc_hd__xnor2_2 _24534_ (.A(_04822_),
    .B(_04823_),
    .Y(_04824_));
 sky130_fd_sc_hd__nand2_1 _24535_ (.A(_04815_),
    .B(_04810_),
    .Y(_04825_));
 sky130_fd_sc_hd__nor2_1 _24536_ (.A(_04061_),
    .B(_04825_),
    .Y(_04826_));
 sky130_fd_sc_hd__o21ai_0 _24537_ (.A1(_04813_),
    .A2(_04826_),
    .B1(_03698_),
    .Y(_04827_));
 sky130_fd_sc_hd__o21ai_1 _24538_ (.A1(_04315_),
    .A2(_04825_),
    .B1(_04827_),
    .Y(_04828_));
 sky130_fd_sc_hd__a21o_1 _24539_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[56] ),
    .A2(_03509_),
    .B1(_03684_),
    .X(_04829_));
 sky130_fd_sc_hd__nand2_1 _24540_ (.A(_04061_),
    .B(_04829_),
    .Y(_04830_));
 sky130_fd_sc_hd__nor3_1 _24541_ (.A(_04061_),
    .B(_04815_),
    .C(_04810_),
    .Y(_04831_));
 sky130_fd_sc_hd__a21oi_1 _24542_ (.A1(_04061_),
    .A2(_04810_),
    .B1(_04831_),
    .Y(_04832_));
 sky130_fd_sc_hd__and3_1 _24543_ (.A(_04182_),
    .B(_04829_),
    .C(_04810_),
    .X(_04833_));
 sky130_fd_sc_hd__o211ai_1 _24544_ (.A1(_04813_),
    .A2(_04833_),
    .B1(_03695_),
    .C1(_04817_),
    .Y(_04834_));
 sky130_fd_sc_hd__o221ai_2 _24545_ (.A1(_04830_),
    .A2(_04825_),
    .B1(_04832_),
    .B2(_03695_),
    .C1(_04834_),
    .Y(_04835_));
 sky130_fd_sc_hd__mux2i_1 _24546_ (.A0(_04828_),
    .A1(_04835_),
    .S(_03516_),
    .Y(_04836_));
 sky130_fd_sc_hd__maj3_2 _24547_ (.A(_04272_),
    .B(_04560_),
    .C(_04733_),
    .X(_04837_));
 sky130_fd_sc_hd__xor2_1 _24548_ (.A(_04836_),
    .B(_04837_),
    .X(_04838_));
 sky130_fd_sc_hd__xnor2_2 _24549_ (.A(_04824_),
    .B(_04838_),
    .Y(_04839_));
 sky130_fd_sc_hd__xnor2_1 _24550_ (.A(_04808_),
    .B(_04839_),
    .Y(_04840_));
 sky130_fd_sc_hd__xnor2_1 _24551_ (.A(_04782_),
    .B(_04840_),
    .Y(_04841_));
 sky130_fd_sc_hd__xnor2_1 _24552_ (.A(_04674_),
    .B(_04702_),
    .Y(_04842_));
 sky130_fd_sc_hd__maj3_1 _24553_ (.A(_04692_),
    .B(_04703_),
    .C(_04842_),
    .X(_04843_));
 sky130_fd_sc_hd__xnor2_1 _24554_ (.A(_04841_),
    .B(_04843_),
    .Y(_04844_));
 sky130_fd_sc_hd__xnor2_2 _24555_ (.A(_04779_),
    .B(_04844_),
    .Y(_04845_));
 sky130_fd_sc_hd__a211o_1 _24556_ (.A1(_04676_),
    .A2(_04738_),
    .B1(_04741_),
    .C1(_04588_),
    .X(_04846_));
 sky130_fd_sc_hd__maj3_1 _24557_ (.A(_04676_),
    .B(_04738_),
    .C(_04740_),
    .X(_04847_));
 sky130_fd_sc_hd__nand2_1 _24558_ (.A(_04846_),
    .B(_04847_),
    .Y(_04848_));
 sky130_fd_sc_hd__xnor2_1 _24559_ (.A(_04845_),
    .B(_04848_),
    .Y(_04849_));
 sky130_fd_sc_hd__xnor2_2 _24560_ (.A(_04776_),
    .B(_04849_),
    .Y(_04850_));
 sky130_fd_sc_hd__nand2_1 _24561_ (.A(_02169_),
    .B(_04850_),
    .Y(_04851_));
 sky130_fd_sc_hd__o21ai_2 _24562_ (.A1(_02169_),
    .A2(_02827_),
    .B1(_04851_),
    .Y(_04852_));
 sky130_fd_sc_hd__mux2i_4 _24563_ (.A0(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[59] ),
    .A1(_04852_),
    .S(_08100_),
    .Y(_04853_));
 sky130_fd_sc_hd__nand3_1 _24564_ (.A(_10497_),
    .B(_10524_),
    .C(_02228_),
    .Y(_04854_));
 sky130_fd_sc_hd__o21ai_0 _24565_ (.A1(_10497_),
    .A2(_01902_),
    .B1(_04854_),
    .Y(_04855_));
 sky130_fd_sc_hd__a21oi_1 _24566_ (.A1(_10497_),
    .A2(_02233_),
    .B1(_10524_),
    .Y(_04856_));
 sky130_fd_sc_hd__a21oi_1 _24567_ (.A1(_02225_),
    .A2(_04855_),
    .B1(_04856_),
    .Y(_04857_));
 sky130_fd_sc_hd__nor2_1 _24568_ (.A(_01773_),
    .B(_01955_),
    .Y(_04858_));
 sky130_fd_sc_hd__a211oi_2 _24569_ (.A1(_01773_),
    .A2(_01944_),
    .B1(_04858_),
    .C1(_01761_),
    .Y(_04859_));
 sky130_fd_sc_hd__a2111oi_0 _24570_ (.A1(net168),
    .A2(_01929_),
    .B1(_04857_),
    .C1(_04859_),
    .D1(net314),
    .Y(_04860_));
 sky130_fd_sc_hd__mux4_1 _24571_ (.A0(net46),
    .A1(net29),
    .A2(net52),
    .A3(net37),
    .S0(\load_store_unit_i.rdata_offset_q[1] ),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .X(_04861_));
 sky130_fd_sc_hd__a21oi_2 _24572_ (.A1(_01674_),
    .A2(_04861_),
    .B1(_03479_),
    .Y(_04862_));
 sky130_fd_sc_hd__a211oi_4 _24573_ (.A1(_04853_),
    .A2(net314),
    .B1(_04860_),
    .C1(_04862_),
    .Y(_04863_));
 sky130_fd_sc_hd__a21oi_2 _24574_ (.A1(_11744_),
    .A2(net265),
    .B1(_04862_),
    .Y(_04864_));
 sky130_fd_sc_hd__or2_4 _24575_ (.A(_04864_),
    .B(_04863_),
    .X(_04865_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_255 ();
 sky130_fd_sc_hd__nand2_2 _24577_ (.A(net1529),
    .B(_02119_),
    .Y(_04867_));
 sky130_fd_sc_hd__nand2_1 _24578_ (.A(\gen_regfile_ff.register_file_i.rf_reg[155] ),
    .B(_02123_),
    .Y(_04868_));
 sky130_fd_sc_hd__nand2_1 _24579_ (.A(_04868_),
    .B(_04867_),
    .Y(_00540_));
 sky130_fd_sc_hd__nor2_1 _24580_ (.A(_10655_),
    .B(_01902_),
    .Y(_04869_));
 sky130_fd_sc_hd__a31oi_1 _24581_ (.A1(_10622_),
    .A2(_10655_),
    .A3(_02228_),
    .B1(_04869_),
    .Y(_04870_));
 sky130_fd_sc_hd__nor2_1 _24582_ (.A(_01893_),
    .B(_04870_),
    .Y(_04871_));
 sky130_fd_sc_hd__a21oi_1 _24583_ (.A1(_10655_),
    .A2(_02233_),
    .B1(_10622_),
    .Y(_04872_));
 sky130_fd_sc_hd__o21ai_0 _24584_ (.A1(_04871_),
    .A2(_04872_),
    .B1(net739),
    .Y(_04873_));
 sky130_fd_sc_hd__nor2_1 _24585_ (.A(_01738_),
    .B(_02835_),
    .Y(_04874_));
 sky130_fd_sc_hd__nor2_1 _24586_ (.A(_01758_),
    .B(_02374_),
    .Y(_04875_));
 sky130_fd_sc_hd__nor2_1 _24587_ (.A(net300),
    .B(_01856_),
    .Y(_04876_));
 sky130_fd_sc_hd__a21oi_1 _24588_ (.A1(net300),
    .A2(_01832_),
    .B1(_04876_),
    .Y(_04877_));
 sky130_fd_sc_hd__nor2_1 _24589_ (.A(_01771_),
    .B(_02190_),
    .Y(_04878_));
 sky130_fd_sc_hd__a211oi_1 _24590_ (.A1(_01771_),
    .A2(_04877_),
    .B1(_04878_),
    .C1(_01748_),
    .Y(_04879_));
 sky130_fd_sc_hd__nor3_1 _24591_ (.A(_01826_),
    .B(_04875_),
    .C(_04879_),
    .Y(_04880_));
 sky130_fd_sc_hd__nand2_1 _24592_ (.A(_02558_),
    .B(_02863_),
    .Y(_04881_));
 sky130_fd_sc_hd__o31ai_2 _24593_ (.A1(_02558_),
    .A2(_04874_),
    .A3(_04880_),
    .B1(_04881_),
    .Y(_04882_));
 sky130_fd_sc_hd__nand2_1 _24594_ (.A(_01762_),
    .B(_04882_),
    .Y(_04883_));
 sky130_fd_sc_hd__nor2_1 _24595_ (.A(_01735_),
    .B(_01743_),
    .Y(_04884_));
 sky130_fd_sc_hd__a21oi_1 _24596_ (.A1(_01743_),
    .A2(_02866_),
    .B1(_04884_),
    .Y(_04885_));
 sky130_fd_sc_hd__nand2_1 _24597_ (.A(_01773_),
    .B(_04885_),
    .Y(_04886_));
 sky130_fd_sc_hd__a21oi_2 _24598_ (.A1(_04883_),
    .A2(_04886_),
    .B1(_01761_),
    .Y(_04887_));
 sky130_fd_sc_hd__a211oi_2 _24599_ (.A1(net169),
    .A2(_01929_),
    .B1(_04873_),
    .C1(_04887_),
    .Y(_04888_));
 sky130_fd_sc_hd__mux2_1 _24600_ (.A0(net47),
    .A1(net30),
    .S(\load_store_unit_i.rdata_offset_q[1] ),
    .X(_04889_));
 sky130_fd_sc_hd__nor2_1 _24601_ (.A(\load_store_unit_i.rdata_offset_q[0] ),
    .B(_04889_),
    .Y(_04890_));
 sky130_fd_sc_hd__a311o_1 _24602_ (.A1(\load_store_unit_i.rdata_offset_q[0] ),
    .A2(_02103_),
    .A3(_02109_),
    .B1(_04890_),
    .C1(_01684_),
    .X(_04891_));
 sky130_fd_sc_hd__nand2_2 _24603_ (.A(_04647_),
    .B(_04891_),
    .Y(_04892_));
 sky130_fd_sc_hd__o21ai_1 _24604_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[60] ),
    .A2(_03724_),
    .B1(_04892_),
    .Y(_04893_));
 sky130_fd_sc_hd__maj3_1 _24605_ (.A(_04779_),
    .B(_04841_),
    .C(_04843_),
    .X(_04894_));
 sky130_fd_sc_hd__xor2_1 _24606_ (.A(_04508_),
    .B(_04808_),
    .X(_04895_));
 sky130_fd_sc_hd__xor2_1 _24607_ (.A(_04501_),
    .B(_04839_),
    .X(_04896_));
 sky130_fd_sc_hd__maj3_1 _24608_ (.A(_04781_),
    .B(_04895_),
    .C(_04896_),
    .X(_04897_));
 sky130_fd_sc_hd__xor2_1 _24609_ (.A(_04508_),
    .B(_04806_),
    .X(_04898_));
 sky130_fd_sc_hd__maj3_1 _24610_ (.A(_04801_),
    .B(_04783_),
    .C(_04898_),
    .X(_04899_));
 sky130_fd_sc_hd__xnor2_1 _24611_ (.A(_04509_),
    .B(_04899_),
    .Y(_04900_));
 sky130_fd_sc_hd__maj3_1 _24612_ (.A(_04796_),
    .B(_04797_),
    .C(_04799_),
    .X(_04901_));
 sky130_fd_sc_hd__nand2_1 _24613_ (.A(_03017_),
    .B(_03274_),
    .Y(_04902_));
 sky130_fd_sc_hd__xnor2_1 _24614_ (.A(_02936_),
    .B(net899),
    .Y(_04903_));
 sky130_fd_sc_hd__nor2_1 _24615_ (.A(_03512_),
    .B(_04903_),
    .Y(_04904_));
 sky130_fd_sc_hd__xnor2_1 _24616_ (.A(_04902_),
    .B(_04904_),
    .Y(_04905_));
 sky130_fd_sc_hd__maj3_1 _24617_ (.A(_04789_),
    .B(_04790_),
    .C(_04791_),
    .X(_04906_));
 sky130_fd_sc_hd__nand2_1 _24618_ (.A(_03041_),
    .B(_03310_),
    .Y(_04907_));
 sky130_fd_sc_hd__nand2_1 _24619_ (.A(_03097_),
    .B(_03376_),
    .Y(_04908_));
 sky130_fd_sc_hd__nand2_1 _24620_ (.A(_03161_),
    .B(_03265_),
    .Y(_04909_));
 sky130_fd_sc_hd__xor2_1 _24621_ (.A(_04908_),
    .B(_04909_),
    .X(_04910_));
 sky130_fd_sc_hd__xnor2_1 _24622_ (.A(_04907_),
    .B(_04910_),
    .Y(_04911_));
 sky130_fd_sc_hd__xor2_1 _24623_ (.A(_04906_),
    .B(_04911_),
    .X(_04912_));
 sky130_fd_sc_hd__xnor2_1 _24624_ (.A(_04905_),
    .B(_04912_),
    .Y(_04913_));
 sky130_fd_sc_hd__maj3_1 _24625_ (.A(_04793_),
    .B(_04788_),
    .C(_04794_),
    .X(_04914_));
 sky130_fd_sc_hd__maj3_1 _24626_ (.A(_04785_),
    .B(_04784_),
    .C(_04786_),
    .X(_04915_));
 sky130_fd_sc_hd__xnor2_1 _24627_ (.A(_04727_),
    .B(_04915_),
    .Y(_04916_));
 sky130_fd_sc_hd__xnor2_1 _24628_ (.A(_04914_),
    .B(_04916_),
    .Y(_04917_));
 sky130_fd_sc_hd__xnor2_1 _24629_ (.A(_04913_),
    .B(_04917_),
    .Y(_04918_));
 sky130_fd_sc_hd__inv_1 _24630_ (.A(_04798_),
    .Y(_04919_));
 sky130_fd_sc_hd__a21oi_1 _24631_ (.A1(_04607_),
    .A2(_04919_),
    .B1(net1161),
    .Y(_04920_));
 sky130_fd_sc_hd__a21oi_1 _24632_ (.A1(_04802_),
    .A2(_04798_),
    .B1(_04920_),
    .Y(_04921_));
 sky130_fd_sc_hd__nor2_2 _24633_ (.A(_03512_),
    .B(_04921_),
    .Y(_04922_));
 sky130_fd_sc_hd__xnor2_1 _24634_ (.A(_04918_),
    .B(_04922_),
    .Y(_04923_));
 sky130_fd_sc_hd__xnor2_2 _24635_ (.A(_04901_),
    .B(_04923_),
    .Y(_04924_));
 sky130_fd_sc_hd__maj3_1 _24636_ (.A(_04272_),
    .B(_04507_),
    .C(_04806_),
    .X(_04925_));
 sky130_fd_sc_hd__nand2_1 _24637_ (.A(_04061_),
    .B(_04823_),
    .Y(_04926_));
 sky130_fd_sc_hd__o21ai_0 _24638_ (.A1(_04816_),
    .A2(_04823_),
    .B1(_04926_),
    .Y(_04927_));
 sky130_fd_sc_hd__nand3_1 _24639_ (.A(_03695_),
    .B(_04810_),
    .C(_04927_),
    .Y(_04928_));
 sky130_fd_sc_hd__nand3_1 _24640_ (.A(_04182_),
    .B(_04810_),
    .C(_04823_),
    .Y(_04929_));
 sky130_fd_sc_hd__o21ai_0 _24641_ (.A1(_04182_),
    .A2(_04823_),
    .B1(_04929_),
    .Y(_04930_));
 sky130_fd_sc_hd__nor2_1 _24642_ (.A(_04810_),
    .B(_04823_),
    .Y(_04931_));
 sky130_fd_sc_hd__nor2_1 _24643_ (.A(_04182_),
    .B(_04817_),
    .Y(_04932_));
 sky130_fd_sc_hd__a22oi_1 _24644_ (.A1(_03698_),
    .A2(_04930_),
    .B1(_04931_),
    .B2(_04932_),
    .Y(_04933_));
 sky130_fd_sc_hd__nand2_1 _24645_ (.A(_04182_),
    .B(_04931_),
    .Y(_04934_));
 sky130_fd_sc_hd__a21oi_1 _24646_ (.A1(_04926_),
    .A2(_04934_),
    .B1(_03695_),
    .Y(_04935_));
 sky130_fd_sc_hd__a211oi_1 _24647_ (.A1(_04205_),
    .A2(_04931_),
    .B1(_04935_),
    .C1(_03516_),
    .Y(_04936_));
 sky130_fd_sc_hd__a31o_1 _24648_ (.A1(_03516_),
    .A2(_04928_),
    .A3(_04933_),
    .B1(_04936_),
    .X(_04937_));
 sky130_fd_sc_hd__xnor2_1 _24649_ (.A(_04925_),
    .B(_04937_),
    .Y(_04938_));
 sky130_fd_sc_hd__a21oi_1 _24650_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[59] ),
    .A2(_03509_),
    .B1(_03684_),
    .Y(_04939_));
 sky130_fd_sc_hd__nand3_1 _24651_ (.A(_03698_),
    .B(_04182_),
    .C(_04939_),
    .Y(_04940_));
 sky130_fd_sc_hd__o21ai_0 _24652_ (.A1(_03698_),
    .A2(_04926_),
    .B1(_04940_),
    .Y(_04941_));
 sky130_fd_sc_hd__nor2_1 _24653_ (.A(_04810_),
    .B(_04939_),
    .Y(_04942_));
 sky130_fd_sc_hd__nor2_1 _24654_ (.A(_04182_),
    .B(_04942_),
    .Y(_04943_));
 sky130_fd_sc_hd__o21ai_0 _24655_ (.A1(_04820_),
    .A2(_04943_),
    .B1(_03695_),
    .Y(_04944_));
 sky130_fd_sc_hd__o211ai_1 _24656_ (.A1(_04061_),
    .A2(_04939_),
    .B1(_04944_),
    .C1(_03516_),
    .Y(_04945_));
 sky130_fd_sc_hd__o21ai_1 _24657_ (.A1(_03516_),
    .A2(_04941_),
    .B1(_04945_),
    .Y(_04946_));
 sky130_fd_sc_hd__a21oi_2 _24658_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[60] ),
    .A2(_03509_),
    .B1(_03684_),
    .Y(_04947_));
 sky130_fd_sc_hd__xnor2_2 _24659_ (.A(_04946_),
    .B(_04947_),
    .Y(_04948_));
 sky130_fd_sc_hd__xnor2_1 _24660_ (.A(_04938_),
    .B(_04948_),
    .Y(_04949_));
 sky130_fd_sc_hd__xnor2_1 _24661_ (.A(_04924_),
    .B(_04949_),
    .Y(_04950_));
 sky130_fd_sc_hd__xnor2_1 _24662_ (.A(_04900_),
    .B(_04950_),
    .Y(_04951_));
 sky130_fd_sc_hd__nor2_1 _24663_ (.A(_04828_),
    .B(_04837_),
    .Y(_04952_));
 sky130_fd_sc_hd__xnor2_1 _24664_ (.A(_04182_),
    .B(_04824_),
    .Y(_04953_));
 sky130_fd_sc_hd__nor2_1 _24665_ (.A(_04952_),
    .B(_04953_),
    .Y(_04954_));
 sky130_fd_sc_hd__a211oi_1 _24666_ (.A1(_04828_),
    .A2(_04837_),
    .B1(_04954_),
    .C1(_03516_),
    .Y(_04955_));
 sky130_fd_sc_hd__maj3_1 _24667_ (.A(_04835_),
    .B(_04837_),
    .C(_04953_),
    .X(_04956_));
 sky130_fd_sc_hd__nor2_1 _24668_ (.A(_03690_),
    .B(_04956_),
    .Y(_04957_));
 sky130_fd_sc_hd__nor2_1 _24669_ (.A(_04955_),
    .B(_04957_),
    .Y(_04958_));
 sky130_fd_sc_hd__xnor2_1 _24670_ (.A(_04951_),
    .B(_04958_),
    .Y(_04959_));
 sky130_fd_sc_hd__xnor2_1 _24671_ (.A(_04897_),
    .B(_04959_),
    .Y(_04960_));
 sky130_fd_sc_hd__nor2_1 _24672_ (.A(_04894_),
    .B(_04960_),
    .Y(_04961_));
 sky130_fd_sc_hd__and2_0 _24673_ (.A(_04894_),
    .B(_04960_),
    .X(_04962_));
 sky130_fd_sc_hd__nor2_1 _24674_ (.A(_04961_),
    .B(_04962_),
    .Y(_04963_));
 sky130_fd_sc_hd__nand2_1 _24675_ (.A(_04411_),
    .B(_04525_),
    .Y(_04964_));
 sky130_fd_sc_hd__a21oi_2 _24676_ (.A1(_04410_),
    .A2(_04407_),
    .B1(_04964_),
    .Y(_04965_));
 sky130_fd_sc_hd__o21bai_2 _24677_ (.A1(_04965_),
    .A2(_04526_),
    .B1_N(_04773_),
    .Y(_04966_));
 sky130_fd_sc_hd__nand2_1 _24678_ (.A(_04966_),
    .B(_04775_),
    .Y(_04967_));
 sky130_fd_sc_hd__maj3_2 _24679_ (.A(_04845_),
    .B(_04967_),
    .C(_04848_),
    .X(_04968_));
 sky130_fd_sc_hd__xnor2_4 _24680_ (.A(_04963_),
    .B(_04968_),
    .Y(_04969_));
 sky130_fd_sc_hd__nand2_4 _24681_ (.A(_02169_),
    .B(_04969_),
    .Y(_04970_));
 sky130_fd_sc_hd__or2_1 _24682_ (.A(_02169_),
    .B(_02968_),
    .X(_04971_));
 sky130_fd_sc_hd__a211oi_4 _24683_ (.A1(_04970_),
    .A2(_04971_),
    .B1(net441),
    .C1(net739),
    .Y(_04972_));
 sky130_fd_sc_hd__nand2_1 _24684_ (.A(_11763_),
    .B(net265),
    .Y(_04973_));
 sky130_fd_sc_hd__nand2_1 _24685_ (.A(_04892_),
    .B(_04973_),
    .Y(_04974_));
 sky130_fd_sc_hd__o31ai_4 _24686_ (.A1(_04888_),
    .A2(_04893_),
    .A3(_04972_),
    .B1(_04974_),
    .Y(_04975_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_254 ();
 sky130_fd_sc_hd__mux2_4 _24688_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[156] ),
    .A1(_04975_),
    .S(_02119_),
    .X(_00541_));
 sky130_fd_sc_hd__nor2_1 _24689_ (.A(_04845_),
    .B(_04848_),
    .Y(_04977_));
 sky130_fd_sc_hd__a21oi_2 _24690_ (.A1(_04845_),
    .A2(_04848_),
    .B1(_04776_),
    .Y(_04978_));
 sky130_fd_sc_hd__nor2_1 _24691_ (.A(_04977_),
    .B(_04978_),
    .Y(_04979_));
 sky130_fd_sc_hd__a21oi_1 _24692_ (.A1(_04894_),
    .A2(_04960_),
    .B1(_04979_),
    .Y(_04980_));
 sky130_fd_sc_hd__nor2_1 _24693_ (.A(_04980_),
    .B(_04961_),
    .Y(_04981_));
 sky130_fd_sc_hd__maj3_1 _24694_ (.A(_04897_),
    .B(_04951_),
    .C(_04958_),
    .X(_04982_));
 sky130_fd_sc_hd__xor2_1 _24695_ (.A(_04508_),
    .B(_04924_),
    .X(_04983_));
 sky130_fd_sc_hd__xor2_1 _24696_ (.A(_04501_),
    .B(_04949_),
    .X(_04984_));
 sky130_fd_sc_hd__maj3_1 _24697_ (.A(_04899_),
    .B(_04983_),
    .C(_04984_),
    .X(_04985_));
 sky130_fd_sc_hd__maj3_1 _24698_ (.A(_04272_),
    .B(_04507_),
    .C(_04922_),
    .X(_04986_));
 sky130_fd_sc_hd__a21o_1 _24699_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[59] ),
    .A2(net311),
    .B1(_03772_),
    .X(_04987_));
 sky130_fd_sc_hd__a21oi_4 _24700_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[60] ),
    .A2(net311),
    .B1(_03772_),
    .Y(_04988_));
 sky130_fd_sc_hd__nand2_1 _24701_ (.A(_04987_),
    .B(_04988_),
    .Y(_04989_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_252 ();
 sky130_fd_sc_hd__a21o_1 _24704_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[60] ),
    .A2(net311),
    .B1(_03772_),
    .X(_04992_));
 sky130_fd_sc_hd__nand2_1 _24705_ (.A(_03937_),
    .B(_04992_),
    .Y(_04993_));
 sky130_fd_sc_hd__o21ai_0 _24706_ (.A1(_03937_),
    .A2(_04989_),
    .B1(_04993_),
    .Y(_04994_));
 sky130_fd_sc_hd__nor2_1 _24707_ (.A(_04352_),
    .B(_04989_),
    .Y(_04995_));
 sky130_fd_sc_hd__a21oi_1 _24708_ (.A1(_03941_),
    .A2(_04994_),
    .B1(_04995_),
    .Y(_04996_));
 sky130_fd_sc_hd__nand2_1 _24709_ (.A(_03937_),
    .B(_04693_),
    .Y(_04997_));
 sky130_fd_sc_hd__nor3_1 _24710_ (.A(_03937_),
    .B(_04987_),
    .C(_04988_),
    .Y(_04998_));
 sky130_fd_sc_hd__a211oi_1 _24711_ (.A1(_03937_),
    .A2(_04988_),
    .B1(_04998_),
    .C1(_03933_),
    .Y(_04999_));
 sky130_fd_sc_hd__nand3_1 _24712_ (.A(_04049_),
    .B(_04693_),
    .C(_04988_),
    .Y(_05000_));
 sky130_fd_sc_hd__a21oi_1 _24713_ (.A1(_04993_),
    .A2(_05000_),
    .B1(_04987_),
    .Y(_05001_));
 sky130_fd_sc_hd__nor2_1 _24714_ (.A(_03941_),
    .B(_05001_),
    .Y(_05002_));
 sky130_fd_sc_hd__o22ai_1 _24715_ (.A1(_04997_),
    .A2(_04989_),
    .B1(_04999_),
    .B2(_05002_),
    .Y(_05003_));
 sky130_fd_sc_hd__nand2_1 _24716_ (.A(_03927_),
    .B(_05003_),
    .Y(_05004_));
 sky130_fd_sc_hd__o21ai_1 _24717_ (.A1(_03927_),
    .A2(_04996_),
    .B1(_05004_),
    .Y(_05005_));
 sky130_fd_sc_hd__xnor2_1 _24718_ (.A(_04986_),
    .B(_05005_),
    .Y(_05006_));
 sky130_fd_sc_hd__nand3_1 _24719_ (.A(_03698_),
    .B(_04182_),
    .C(_04947_),
    .Y(_05007_));
 sky130_fd_sc_hd__o21ai_0 _24720_ (.A1(_03941_),
    .A2(_04993_),
    .B1(_05007_),
    .Y(_05008_));
 sky130_fd_sc_hd__a21oi_1 _24721_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[59] ),
    .A2(net311),
    .B1(_03772_),
    .Y(_05009_));
 sky130_fd_sc_hd__nand3_1 _24722_ (.A(_03933_),
    .B(_03937_),
    .C(_05009_),
    .Y(_05010_));
 sky130_fd_sc_hd__o221ai_1 _24723_ (.A1(_03937_),
    .A2(_04988_),
    .B1(_04989_),
    .B2(_03941_),
    .C1(_05010_),
    .Y(_05011_));
 sky130_fd_sc_hd__mux2i_2 _24724_ (.A0(_05008_),
    .A1(_05011_),
    .S(_03927_),
    .Y(_05012_));
 sky130_fd_sc_hd__a21oi_4 _24725_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[61] ),
    .A2(net311),
    .B1(_03772_),
    .Y(_05013_));
 sky130_fd_sc_hd__xnor2_2 _24726_ (.A(_05012_),
    .B(_05013_),
    .Y(_05014_));
 sky130_fd_sc_hd__xnor2_1 _24727_ (.A(_05006_),
    .B(_05014_),
    .Y(_05015_));
 sky130_fd_sc_hd__maj3_1 _24728_ (.A(_04908_),
    .B(_04909_),
    .C(_04907_),
    .X(_05016_));
 sky130_fd_sc_hd__nand2_1 _24729_ (.A(_03100_),
    .B(_03376_),
    .Y(_05017_));
 sky130_fd_sc_hd__nand2_1 _24730_ (.A(_03161_),
    .B(_03274_),
    .Y(_05018_));
 sky130_fd_sc_hd__nand2_1 _24731_ (.A(_03265_),
    .B(_03310_),
    .Y(_05019_));
 sky130_fd_sc_hd__xor2_1 _24732_ (.A(_05018_),
    .B(_05019_),
    .X(_05020_));
 sky130_fd_sc_hd__xor2_1 _24733_ (.A(_05017_),
    .B(_05020_),
    .X(_05021_));
 sky130_fd_sc_hd__or2_0 _24734_ (.A(_05016_),
    .B(_05021_),
    .X(_05022_));
 sky130_fd_sc_hd__nand2_1 _24735_ (.A(_05016_),
    .B(_05021_),
    .Y(_05023_));
 sky130_fd_sc_hd__nand2_1 _24736_ (.A(_05022_),
    .B(_05023_),
    .Y(_05024_));
 sky130_fd_sc_hd__maj3_1 _24737_ (.A(_04905_),
    .B(_04906_),
    .C(_04911_),
    .X(_05025_));
 sky130_fd_sc_hd__xnor2_2 _24738_ (.A(net1266),
    .B(_04903_),
    .Y(_05026_));
 sky130_fd_sc_hd__nor2_1 _24739_ (.A(_03512_),
    .B(_05026_),
    .Y(_05027_));
 sky130_fd_sc_hd__maj3_1 _24740_ (.A(_02936_),
    .B(net899),
    .C(_04902_),
    .X(_05028_));
 sky130_fd_sc_hd__nand2b_1 _24741_ (.A_N(_05028_),
    .B(_03689_),
    .Y(_05029_));
 sky130_fd_sc_hd__xor2_2 _24742_ (.A(_04727_),
    .B(_05029_),
    .X(_05030_));
 sky130_fd_sc_hd__xnor2_2 _24743_ (.A(_05027_),
    .B(_05030_),
    .Y(_05031_));
 sky130_fd_sc_hd__xor2_1 _24744_ (.A(_05025_),
    .B(_05031_),
    .X(_05032_));
 sky130_fd_sc_hd__xnor2_2 _24745_ (.A(_05024_),
    .B(_05032_),
    .Y(_05033_));
 sky130_fd_sc_hd__maj3_1 _24746_ (.A(_04913_),
    .B(_04914_),
    .C(_04916_),
    .X(_05034_));
 sky130_fd_sc_hd__inv_1 _24747_ (.A(_04915_),
    .Y(_05035_));
 sky130_fd_sc_hd__a21oi_1 _24748_ (.A1(_04607_),
    .A2(_05035_),
    .B1(net1161),
    .Y(_05036_));
 sky130_fd_sc_hd__a21oi_1 _24749_ (.A1(_04802_),
    .A2(_04915_),
    .B1(_05036_),
    .Y(_05037_));
 sky130_fd_sc_hd__nor2_2 _24750_ (.A(_03512_),
    .B(_05037_),
    .Y(_05038_));
 sky130_fd_sc_hd__xnor2_1 _24751_ (.A(_05034_),
    .B(_05038_),
    .Y(_05039_));
 sky130_fd_sc_hd__xnor2_2 _24752_ (.A(_05033_),
    .B(_05039_),
    .Y(_05040_));
 sky130_fd_sc_hd__xnor2_1 _24753_ (.A(_04509_),
    .B(_05040_),
    .Y(_05041_));
 sky130_fd_sc_hd__xor2_1 _24754_ (.A(_04508_),
    .B(_04922_),
    .X(_05042_));
 sky130_fd_sc_hd__maj3_2 _24755_ (.A(_04918_),
    .B(_04901_),
    .C(_05042_),
    .X(_05043_));
 sky130_fd_sc_hd__xnor2_1 _24756_ (.A(_05041_),
    .B(_05043_),
    .Y(_05044_));
 sky130_fd_sc_hd__xnor2_1 _24757_ (.A(_05015_),
    .B(_05044_),
    .Y(_05045_));
 sky130_fd_sc_hd__inv_1 _24758_ (.A(_04937_),
    .Y(_05046_));
 sky130_fd_sc_hd__xor2_1 _24759_ (.A(_04501_),
    .B(_04948_),
    .X(_05047_));
 sky130_fd_sc_hd__maj3_1 _24760_ (.A(_04925_),
    .B(_05046_),
    .C(_05047_),
    .X(_05048_));
 sky130_fd_sc_hd__nand2_1 _24761_ (.A(_05045_),
    .B(_05048_),
    .Y(_05049_));
 sky130_fd_sc_hd__or2_0 _24762_ (.A(_05045_),
    .B(_05048_),
    .X(_05050_));
 sky130_fd_sc_hd__nand2_1 _24763_ (.A(_05049_),
    .B(_05050_),
    .Y(_05051_));
 sky130_fd_sc_hd__xor2_1 _24764_ (.A(_04985_),
    .B(_05051_),
    .X(_05052_));
 sky130_fd_sc_hd__and2_1 _24765_ (.A(_04982_),
    .B(_05052_),
    .X(_05053_));
 sky130_fd_sc_hd__nor2_1 _24766_ (.A(_04982_),
    .B(_05052_),
    .Y(_05054_));
 sky130_fd_sc_hd__nor2_1 _24767_ (.A(_05053_),
    .B(_05054_),
    .Y(_05055_));
 sky130_fd_sc_hd__xnor2_2 _24768_ (.A(_05055_),
    .B(_04981_),
    .Y(_05056_));
 sky130_fd_sc_hd__nand2_1 _24769_ (.A(_01698_),
    .B(_03073_),
    .Y(_05057_));
 sky130_fd_sc_hd__o21ai_4 _24770_ (.A1(_01698_),
    .A2(_05056_),
    .B1(_05057_),
    .Y(_05058_));
 sky130_fd_sc_hd__nor2_8 _24771_ (.A(net441),
    .B(_05058_),
    .Y(_05059_));
 sky130_fd_sc_hd__o21ai_1 _24772_ (.A1(_08100_),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[61] ),
    .B1(net314),
    .Y(_05060_));
 sky130_fd_sc_hd__nor4_4 _24773_ (.A(_08581_),
    .B(_11774_),
    .C(_11777_),
    .D(_11781_),
    .Y(_05061_));
 sky130_fd_sc_hd__nand3_1 _24774_ (.A(_10561_),
    .B(_10592_),
    .C(_02228_),
    .Y(_05062_));
 sky130_fd_sc_hd__o21ai_0 _24775_ (.A1(_10561_),
    .A2(_01902_),
    .B1(_05062_),
    .Y(_05063_));
 sky130_fd_sc_hd__a21oi_1 _24776_ (.A1(_10561_),
    .A2(_02233_),
    .B1(_10592_),
    .Y(_05064_));
 sky130_fd_sc_hd__a21oi_1 _24777_ (.A1(_02225_),
    .A2(_05063_),
    .B1(_05064_),
    .Y(_05065_));
 sky130_fd_sc_hd__nor2_1 _24778_ (.A(_01771_),
    .B(_01834_),
    .Y(_05066_));
 sky130_fd_sc_hd__nor2_1 _24779_ (.A(_01751_),
    .B(_01857_),
    .Y(_05067_));
 sky130_fd_sc_hd__nand2_1 _24780_ (.A(_01748_),
    .B(_02268_),
    .Y(_05068_));
 sky130_fd_sc_hd__o311ai_2 _24781_ (.A1(_01748_),
    .A2(_05066_),
    .A3(_05067_),
    .B1(_01738_),
    .C1(_05068_),
    .Y(_05069_));
 sky130_fd_sc_hd__o211ai_1 _24782_ (.A1(_01738_),
    .A2(_02661_),
    .B1(_05069_),
    .C1(_01743_),
    .Y(_05070_));
 sky130_fd_sc_hd__o21ai_1 _24783_ (.A1(_01743_),
    .A2(_02986_),
    .B1(_05070_),
    .Y(_05071_));
 sky130_fd_sc_hd__nand2_1 _24784_ (.A(net295),
    .B(_05071_),
    .Y(_05072_));
 sky130_fd_sc_hd__a21oi_1 _24785_ (.A1(_01743_),
    .A2(_02983_),
    .B1(_04884_),
    .Y(_05073_));
 sky130_fd_sc_hd__nand2_1 _24786_ (.A(_01773_),
    .B(_05073_),
    .Y(_05074_));
 sky130_fd_sc_hd__a21oi_2 _24787_ (.A1(_05072_),
    .A2(_05074_),
    .B1(_01761_),
    .Y(_05075_));
 sky130_fd_sc_hd__nor2_1 _24788_ (.A(_05065_),
    .B(_05075_),
    .Y(_05076_));
 sky130_fd_sc_hd__o21ai_1 _24789_ (.A1(_10665_),
    .A2(_01889_),
    .B1(_05076_),
    .Y(_05077_));
 sky130_fd_sc_hd__a21oi_2 _24790_ (.A1(net739),
    .A2(_05077_),
    .B1(_08632_),
    .Y(_05078_));
 sky130_fd_sc_hd__o221ai_4 _24791_ (.A1(_05059_),
    .A2(_05060_),
    .B1(_05061_),
    .B2(_05078_),
    .C1(net265),
    .Y(_05079_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_251 ();
 sky130_fd_sc_hd__mux2_1 _24793_ (.A0(net48),
    .A1(net31),
    .S(\load_store_unit_i.rdata_offset_q[1] ),
    .X(_05081_));
 sky130_fd_sc_hd__nor2_1 _24794_ (.A(\load_store_unit_i.rdata_offset_q[0] ),
    .B(_05081_),
    .Y(_05082_));
 sky130_fd_sc_hd__a31oi_4 _24795_ (.A1(\load_store_unit_i.rdata_offset_q[0] ),
    .A2(_02241_),
    .A3(_02247_),
    .B1(_05082_),
    .Y(_05083_));
 sky130_fd_sc_hd__a21oi_4 _24796_ (.A1(_01674_),
    .A2(_05083_),
    .B1(_03479_),
    .Y(_05084_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_250 ();
 sky130_fd_sc_hd__nor2_1 _24798_ (.A(_02123_),
    .B(_05084_),
    .Y(_05086_));
 sky130_fd_sc_hd__a22o_1 _24799_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[157] ),
    .A2(_02123_),
    .B1(_05086_),
    .B2(_05079_),
    .X(_00542_));
 sky130_fd_sc_hd__inv_1 _24800_ (.A(_05050_),
    .Y(_05087_));
 sky130_fd_sc_hd__o21ai_1 _24801_ (.A1(_04985_),
    .A2(_05087_),
    .B1(_05049_),
    .Y(_05088_));
 sky130_fd_sc_hd__xnor2_1 _24802_ (.A(_04508_),
    .B(_05040_),
    .Y(_05089_));
 sky130_fd_sc_hd__xor2_1 _24803_ (.A(_04674_),
    .B(_05015_),
    .X(_05090_));
 sky130_fd_sc_hd__maj3_1 _24804_ (.A(_05043_),
    .B(_05089_),
    .C(_05090_),
    .X(_05091_));
 sky130_fd_sc_hd__a21o_2 _24805_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[62] ),
    .A2(net311),
    .B1(_03772_),
    .X(_05092_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_249 ();
 sky130_fd_sc_hd__nand2_1 _24807_ (.A(_04049_),
    .B(_05013_),
    .Y(_05094_));
 sky130_fd_sc_hd__a21o_1 _24808_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[61] ),
    .A2(net311),
    .B1(_03772_),
    .X(_05095_));
 sky130_fd_sc_hd__nand2_1 _24809_ (.A(_04049_),
    .B(_05095_),
    .Y(_05096_));
 sky130_fd_sc_hd__nor2_1 _24810_ (.A(_04049_),
    .B(_05095_),
    .Y(_05097_));
 sky130_fd_sc_hd__a311oi_1 _24811_ (.A1(_03927_),
    .A2(_04988_),
    .A3(_05096_),
    .B1(_05097_),
    .C1(_03941_),
    .Y(_05098_));
 sky130_fd_sc_hd__a31oi_1 _24812_ (.A1(_03941_),
    .A2(_04672_),
    .A3(_05094_),
    .B1(_05098_),
    .Y(_05099_));
 sky130_fd_sc_hd__xnor2_1 _24813_ (.A(_05092_),
    .B(_05099_),
    .Y(_05100_));
 sky130_fd_sc_hd__nand2_1 _24814_ (.A(_04992_),
    .B(_05013_),
    .Y(_05101_));
 sky130_fd_sc_hd__nor2_1 _24815_ (.A(_03937_),
    .B(_05013_),
    .Y(_05102_));
 sky130_fd_sc_hd__a211oi_1 _24816_ (.A1(_04988_),
    .A2(_05102_),
    .B1(_05097_),
    .C1(_03933_),
    .Y(_05103_));
 sky130_fd_sc_hd__nand2_1 _24817_ (.A(_03937_),
    .B(_05095_),
    .Y(_05104_));
 sky130_fd_sc_hd__o21ai_0 _24818_ (.A1(_05009_),
    .A2(_05094_),
    .B1(_05104_),
    .Y(_05105_));
 sky130_fd_sc_hd__a21oi_1 _24819_ (.A1(_04988_),
    .A2(_05105_),
    .B1(_03941_),
    .Y(_05106_));
 sky130_fd_sc_hd__o32ai_1 _24820_ (.A1(_04049_),
    .A2(_05009_),
    .A3(_05101_),
    .B1(_05103_),
    .B2(_05106_),
    .Y(_05107_));
 sky130_fd_sc_hd__o21ai_0 _24821_ (.A1(_03937_),
    .A2(_05101_),
    .B1(_05104_),
    .Y(_05108_));
 sky130_fd_sc_hd__nor2_1 _24822_ (.A(_04352_),
    .B(_05101_),
    .Y(_05109_));
 sky130_fd_sc_hd__a21oi_1 _24823_ (.A1(_03941_),
    .A2(_05108_),
    .B1(_05109_),
    .Y(_05110_));
 sky130_fd_sc_hd__nor2_1 _24824_ (.A(_03927_),
    .B(_05110_),
    .Y(_05111_));
 sky130_fd_sc_hd__a21oi_1 _24825_ (.A1(_03927_),
    .A2(_05107_),
    .B1(_05111_),
    .Y(_05112_));
 sky130_fd_sc_hd__a21o_1 _24826_ (.A1(_04507_),
    .A2(_05038_),
    .B1(_04272_),
    .X(_05113_));
 sky130_fd_sc_hd__o21ai_2 _24827_ (.A1(_04507_),
    .A2(_05038_),
    .B1(_05113_),
    .Y(_05114_));
 sky130_fd_sc_hd__xor2_1 _24828_ (.A(_05112_),
    .B(_05114_),
    .X(_05115_));
 sky130_fd_sc_hd__xnor2_1 _24829_ (.A(_05100_),
    .B(_05115_),
    .Y(_05116_));
 sky130_fd_sc_hd__nor2_1 _24830_ (.A(_03670_),
    .B(_05028_),
    .Y(_05117_));
 sky130_fd_sc_hd__a21oi_1 _24831_ (.A1(_04607_),
    .A2(_05029_),
    .B1(net1161),
    .Y(_05118_));
 sky130_fd_sc_hd__a21oi_1 _24832_ (.A1(_04802_),
    .A2(_05117_),
    .B1(_05118_),
    .Y(_05119_));
 sky130_fd_sc_hd__nor2_2 _24833_ (.A(_03512_),
    .B(_05119_),
    .Y(_05120_));
 sky130_fd_sc_hd__xnor2_2 _24834_ (.A(_04508_),
    .B(_05120_),
    .Y(_05121_));
 sky130_fd_sc_hd__a21boi_2 _24835_ (.A1(_05023_),
    .A2(_05027_),
    .B1_N(_05022_),
    .Y(_05122_));
 sky130_fd_sc_hd__maj3_1 _24836_ (.A(_05018_),
    .B(_05019_),
    .C(_05017_),
    .X(_05123_));
 sky130_fd_sc_hd__nor2_1 _24837_ (.A(_03313_),
    .B(_03512_),
    .Y(_05124_));
 sky130_fd_sc_hd__nor2_1 _24838_ (.A(_04020_),
    .B(_03373_),
    .Y(_05125_));
 sky130_fd_sc_hd__xnor2_1 _24839_ (.A(_05124_),
    .B(_05125_),
    .Y(_05126_));
 sky130_fd_sc_hd__nand2_1 _24840_ (.A(_03119_),
    .B(_03376_),
    .Y(_05127_));
 sky130_fd_sc_hd__xnor2_1 _24841_ (.A(_05126_),
    .B(_05127_),
    .Y(_05128_));
 sky130_fd_sc_hd__xnor2_1 _24842_ (.A(_05123_),
    .B(_05128_),
    .Y(_05129_));
 sky130_fd_sc_hd__xnor2_1 _24843_ (.A(_05122_),
    .B(_05129_),
    .Y(_05130_));
 sky130_fd_sc_hd__xnor2_1 _24844_ (.A(_05031_),
    .B(_05130_),
    .Y(_05131_));
 sky130_fd_sc_hd__nor2_1 _24845_ (.A(_03670_),
    .B(_04726_),
    .Y(_05132_));
 sky130_fd_sc_hd__xnor2_2 _24846_ (.A(_05132_),
    .B(_05117_),
    .Y(_05133_));
 sky130_fd_sc_hd__nand2b_1 _24847_ (.A_N(_05026_),
    .B(_03689_),
    .Y(_05134_));
 sky130_fd_sc_hd__xnor2_1 _24848_ (.A(_05024_),
    .B(_05134_),
    .Y(_05135_));
 sky130_fd_sc_hd__nor2_1 _24849_ (.A(_05030_),
    .B(_05135_),
    .Y(_05136_));
 sky130_fd_sc_hd__nor2_1 _24850_ (.A(_05025_),
    .B(_05136_),
    .Y(_05137_));
 sky130_fd_sc_hd__a21oi_2 _24851_ (.A1(_05133_),
    .A2(_05135_),
    .B1(_05137_),
    .Y(_05138_));
 sky130_fd_sc_hd__xnor2_1 _24852_ (.A(_05131_),
    .B(_05138_),
    .Y(_05139_));
 sky130_fd_sc_hd__xnor2_2 _24853_ (.A(_05121_),
    .B(_05139_),
    .Y(_05140_));
 sky130_fd_sc_hd__inv_1 _24854_ (.A(_05034_),
    .Y(_05141_));
 sky130_fd_sc_hd__xnor2_1 _24855_ (.A(_04508_),
    .B(_05038_),
    .Y(_05142_));
 sky130_fd_sc_hd__maj3_2 _24856_ (.A(_05033_),
    .B(_05141_),
    .C(_05142_),
    .X(_05143_));
 sky130_fd_sc_hd__xnor2_1 _24857_ (.A(_05140_),
    .B(_05143_),
    .Y(_05144_));
 sky130_fd_sc_hd__xnor2_1 _24858_ (.A(_05116_),
    .B(_05144_),
    .Y(_05145_));
 sky130_fd_sc_hd__xnor2_1 _24859_ (.A(_04674_),
    .B(_05014_),
    .Y(_05146_));
 sky130_fd_sc_hd__maj3_1 _24860_ (.A(_04986_),
    .B(_05005_),
    .C(_05146_),
    .X(_05147_));
 sky130_fd_sc_hd__xor2_1 _24861_ (.A(_05145_),
    .B(_05147_),
    .X(_05148_));
 sky130_fd_sc_hd__xnor2_1 _24862_ (.A(_05091_),
    .B(_05148_),
    .Y(_05149_));
 sky130_fd_sc_hd__and2_0 _24863_ (.A(_05088_),
    .B(_05149_),
    .X(_05150_));
 sky130_fd_sc_hd__nor2_1 _24864_ (.A(_05088_),
    .B(_05149_),
    .Y(_05151_));
 sky130_fd_sc_hd__nor2_1 _24865_ (.A(_05150_),
    .B(_05151_),
    .Y(_05152_));
 sky130_fd_sc_hd__nor2_1 _24866_ (.A(_05053_),
    .B(_05152_),
    .Y(_05153_));
 sky130_fd_sc_hd__a221oi_2 _24867_ (.A1(_04846_),
    .A2(_04847_),
    .B1(_04966_),
    .B2(_04775_),
    .C1(_04961_),
    .Y(_05154_));
 sky130_fd_sc_hd__o22ai_2 _24868_ (.A1(_04982_),
    .A2(_05052_),
    .B1(_04962_),
    .B2(_05154_),
    .Y(_05155_));
 sky130_fd_sc_hd__o21ai_0 _24869_ (.A1(_04640_),
    .A2(_04744_),
    .B1(_04670_),
    .Y(_05156_));
 sky130_fd_sc_hd__nand2_1 _24870_ (.A(_04640_),
    .B(_04744_),
    .Y(_05157_));
 sky130_fd_sc_hd__a2bb2oi_2 _24871_ (.A1_N(_04774_),
    .A2_N(_04665_),
    .B1(_05156_),
    .B2(_05157_),
    .Y(_05158_));
 sky130_fd_sc_hd__nor2_1 _24872_ (.A(_04961_),
    .B(_05054_),
    .Y(_05159_));
 sky130_fd_sc_hd__o211ai_2 _24873_ (.A1(_05158_),
    .A2(_04848_),
    .B1(_05159_),
    .C1(_04845_),
    .Y(_05160_));
 sky130_fd_sc_hd__nand2_2 _24874_ (.A(_05155_),
    .B(_05160_),
    .Y(_05161_));
 sky130_fd_sc_hd__mux2i_4 _24875_ (.A0(_05153_),
    .A1(_05152_),
    .S(_05161_),
    .Y(_05162_));
 sky130_fd_sc_hd__nand3_1 _24876_ (.A(_02169_),
    .B(_05053_),
    .C(_05152_),
    .Y(_05163_));
 sky130_fd_sc_hd__o21ai_1 _24877_ (.A1(_02169_),
    .A2(_03192_),
    .B1(_05163_),
    .Y(_05164_));
 sky130_fd_sc_hd__nand2_1 _24878_ (.A(net441),
    .B(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[62] ),
    .Y(_05165_));
 sky130_fd_sc_hd__o21ai_1 _24879_ (.A1(net441),
    .A2(_05164_),
    .B1(_05165_),
    .Y(_05166_));
 sky130_fd_sc_hd__o311ai_4 _24880_ (.A1(net441),
    .A2(_01698_),
    .A3(_05162_),
    .B1(_05166_),
    .C1(net312),
    .Y(_05167_));
 sky130_fd_sc_hd__nand3_1 _24881_ (.A(_10764_),
    .B(_10799_),
    .C(_02228_),
    .Y(_05168_));
 sky130_fd_sc_hd__o21ai_0 _24882_ (.A1(_10799_),
    .A2(_01902_),
    .B1(_05168_),
    .Y(_05169_));
 sky130_fd_sc_hd__a21oi_1 _24883_ (.A1(_10799_),
    .A2(_02233_),
    .B1(_10764_),
    .Y(_05170_));
 sky130_fd_sc_hd__a21oi_1 _24884_ (.A1(_02225_),
    .A2(_05169_),
    .B1(_05170_),
    .Y(_05171_));
 sky130_fd_sc_hd__nor2_1 _24885_ (.A(net300),
    .B(_01848_),
    .Y(_05172_));
 sky130_fd_sc_hd__a21oi_1 _24886_ (.A1(net300),
    .A2(_01854_),
    .B1(_05172_),
    .Y(_05173_));
 sky130_fd_sc_hd__nand2_1 _24887_ (.A(_01751_),
    .B(_04877_),
    .Y(_05174_));
 sky130_fd_sc_hd__o211ai_2 _24888_ (.A1(_01751_),
    .A2(_05173_),
    .B1(_05174_),
    .C1(_01758_),
    .Y(_05175_));
 sky130_fd_sc_hd__o211ai_1 _24889_ (.A1(_01758_),
    .A2(_02193_),
    .B1(_05175_),
    .C1(_01738_),
    .Y(_05176_));
 sky130_fd_sc_hd__o21ai_1 _24890_ (.A1(_01738_),
    .A2(_02564_),
    .B1(_05176_),
    .Y(_05177_));
 sky130_fd_sc_hd__nor2_1 _24891_ (.A(_02558_),
    .B(_05177_),
    .Y(_05178_));
 sky130_fd_sc_hd__a21o_1 _24892_ (.A1(_02558_),
    .A2(_03206_),
    .B1(_05178_),
    .X(_05179_));
 sky130_fd_sc_hd__nand2_1 _24893_ (.A(net295),
    .B(_05179_),
    .Y(_05180_));
 sky130_fd_sc_hd__a21oi_1 _24894_ (.A1(_01743_),
    .A2(_03201_),
    .B1(_04884_),
    .Y(_05181_));
 sky130_fd_sc_hd__nand2_1 _24895_ (.A(_01773_),
    .B(_05181_),
    .Y(_05182_));
 sky130_fd_sc_hd__a21oi_1 _24896_ (.A1(_05180_),
    .A2(_05182_),
    .B1(_01761_),
    .Y(_05183_));
 sky130_fd_sc_hd__a211oi_1 _24897_ (.A1(net172),
    .A2(_01929_),
    .B1(_05171_),
    .C1(_05183_),
    .Y(_05184_));
 sky130_fd_sc_hd__o21ai_1 _24898_ (.A1(net313),
    .A2(_05184_),
    .B1(_08581_),
    .Y(_05185_));
 sky130_fd_sc_hd__o21ai_4 _24899_ (.A1(_08581_),
    .A2(_11806_),
    .B1(_05185_),
    .Y(_05186_));
 sky130_fd_sc_hd__mux2_1 _24900_ (.A0(net50),
    .A1(net32),
    .S(\load_store_unit_i.rdata_offset_q[1] ),
    .X(_05187_));
 sky130_fd_sc_hd__nor2_1 _24901_ (.A(\load_store_unit_i.rdata_offset_q[0] ),
    .B(_05187_),
    .Y(_05188_));
 sky130_fd_sc_hd__a31oi_2 _24902_ (.A1(\load_store_unit_i.rdata_offset_q[0] ),
    .A2(_02351_),
    .A3(_02357_),
    .B1(_05188_),
    .Y(_05189_));
 sky130_fd_sc_hd__a21oi_4 _24903_ (.A1(_01674_),
    .A2(_05189_),
    .B1(_03479_),
    .Y(_05190_));
 sky130_fd_sc_hd__a31oi_4 _24904_ (.A1(net266),
    .A2(net860),
    .A3(_05186_),
    .B1(_05190_),
    .Y(_05191_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_248 ();
 sky130_fd_sc_hd__mux2_4 _24906_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[158] ),
    .A1(_05191_),
    .S(_02119_),
    .X(_00543_));
 sky130_fd_sc_hd__nor2_1 _24907_ (.A(net314),
    .B(_02646_),
    .Y(_05193_));
 sky130_fd_sc_hd__nor2_1 _24908_ (.A(_04962_),
    .B(_05053_),
    .Y(_05194_));
 sky130_fd_sc_hd__nor2_1 _24909_ (.A(_05054_),
    .B(_05194_),
    .Y(_05195_));
 sky130_fd_sc_hd__nor4_4 _24910_ (.A(_05054_),
    .B(_04961_),
    .C(_04977_),
    .D(_04978_),
    .Y(_05196_));
 sky130_fd_sc_hd__o21ai_1 _24911_ (.A1(_05196_),
    .A2(_05195_),
    .B1(_05088_),
    .Y(_05197_));
 sky130_fd_sc_hd__o31ai_1 _24912_ (.A1(_05088_),
    .A2(_05195_),
    .A3(_05196_),
    .B1(_05149_),
    .Y(_05198_));
 sky130_fd_sc_hd__nand2_2 _24913_ (.A(_05198_),
    .B(_05197_),
    .Y(_05199_));
 sky130_fd_sc_hd__maj3_1 _24914_ (.A(_05116_),
    .B(_05140_),
    .C(_05143_),
    .X(_05200_));
 sky130_fd_sc_hd__maj3_1 _24915_ (.A(_05134_),
    .B(_05123_),
    .C(_05128_),
    .X(_05201_));
 sky130_fd_sc_hd__nor2_1 _24916_ (.A(_04020_),
    .B(_05127_),
    .Y(_05202_));
 sky130_fd_sc_hd__a21oi_1 _24917_ (.A1(_03689_),
    .A2(_05202_),
    .B1(_03373_),
    .Y(_05203_));
 sky130_fd_sc_hd__nor2_1 _24918_ (.A(_03370_),
    .B(_04023_),
    .Y(_05204_));
 sky130_fd_sc_hd__o22a_1 _24919_ (.A1(_03161_),
    .A2(_05203_),
    .B1(_05204_),
    .B2(_03428_),
    .X(_05205_));
 sky130_fd_sc_hd__xnor2_1 _24920_ (.A(_05201_),
    .B(_05205_),
    .Y(_05206_));
 sky130_fd_sc_hd__xor2_1 _24921_ (.A(_05031_),
    .B(_05206_),
    .X(_05207_));
 sky130_fd_sc_hd__xnor2_1 _24922_ (.A(_05134_),
    .B(_05129_),
    .Y(_05208_));
 sky130_fd_sc_hd__maj3_1 _24923_ (.A(_05030_),
    .B(_05122_),
    .C(_05208_),
    .X(_05209_));
 sky130_fd_sc_hd__xnor2_1 _24924_ (.A(_05207_),
    .B(_05209_),
    .Y(_05210_));
 sky130_fd_sc_hd__xor2_2 _24925_ (.A(_05121_),
    .B(_05210_),
    .X(_05211_));
 sky130_fd_sc_hd__maj3_2 _24926_ (.A(_05131_),
    .B(_05138_),
    .C(_05121_),
    .X(_05212_));
 sky130_fd_sc_hd__xor2_1 _24927_ (.A(_05211_),
    .B(_05212_),
    .X(_05213_));
 sky130_fd_sc_hd__a21oi_4 _24928_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[63] ),
    .A2(net311),
    .B1(_03772_),
    .Y(_05214_));
 sky130_fd_sc_hd__a21oi_2 _24929_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[62] ),
    .A2(net311),
    .B1(_03772_),
    .Y(_05215_));
 sky130_fd_sc_hd__nand2_1 _24930_ (.A(_04049_),
    .B(_05215_),
    .Y(_05216_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_247 ();
 sky130_fd_sc_hd__nand2_1 _24932_ (.A(_04049_),
    .B(_05092_),
    .Y(_05218_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_246 ();
 sky130_fd_sc_hd__nor2_1 _24934_ (.A(_04049_),
    .B(_05092_),
    .Y(_05220_));
 sky130_fd_sc_hd__a311oi_1 _24935_ (.A1(_03927_),
    .A2(_05013_),
    .A3(_05218_),
    .B1(_05220_),
    .C1(_03941_),
    .Y(_05221_));
 sky130_fd_sc_hd__a31oi_1 _24936_ (.A1(_03941_),
    .A2(_04672_),
    .A3(_05216_),
    .B1(_05221_),
    .Y(_05222_));
 sky130_fd_sc_hd__xnor2_1 _24937_ (.A(_05214_),
    .B(_05222_),
    .Y(_05223_));
 sky130_fd_sc_hd__a21o_1 _24938_ (.A1(_04507_),
    .A2(_05120_),
    .B1(_04272_),
    .X(_05224_));
 sky130_fd_sc_hd__o21ai_4 _24939_ (.A1(_04507_),
    .A2(_05120_),
    .B1(_05224_),
    .Y(_05225_));
 sky130_fd_sc_hd__nand2_1 _24940_ (.A(_05095_),
    .B(_05215_),
    .Y(_05226_));
 sky130_fd_sc_hd__nand2_1 _24941_ (.A(_03937_),
    .B(_05092_),
    .Y(_05227_));
 sky130_fd_sc_hd__o21ai_0 _24942_ (.A1(_03937_),
    .A2(_05226_),
    .B1(_05227_),
    .Y(_05228_));
 sky130_fd_sc_hd__nor2_1 _24943_ (.A(_04352_),
    .B(_05226_),
    .Y(_05229_));
 sky130_fd_sc_hd__a21oi_1 _24944_ (.A1(_03941_),
    .A2(_05228_),
    .B1(_05229_),
    .Y(_05230_));
 sky130_fd_sc_hd__nor2_1 _24945_ (.A(_05095_),
    .B(_05218_),
    .Y(_05231_));
 sky130_fd_sc_hd__nor3_1 _24946_ (.A(_03933_),
    .B(_05220_),
    .C(_05231_),
    .Y(_05232_));
 sky130_fd_sc_hd__o21ai_0 _24947_ (.A1(_04988_),
    .A2(_05216_),
    .B1(_05227_),
    .Y(_05233_));
 sky130_fd_sc_hd__a21oi_1 _24948_ (.A1(_05013_),
    .A2(_05233_),
    .B1(_03941_),
    .Y(_05234_));
 sky130_fd_sc_hd__o22ai_1 _24949_ (.A1(_04993_),
    .A2(_05226_),
    .B1(_05232_),
    .B2(_05234_),
    .Y(_05235_));
 sky130_fd_sc_hd__nand2_1 _24950_ (.A(_03927_),
    .B(_05235_),
    .Y(_05236_));
 sky130_fd_sc_hd__o21ai_1 _24951_ (.A1(_03927_),
    .A2(_05230_),
    .B1(_05236_),
    .Y(_05237_));
 sky130_fd_sc_hd__xor2_1 _24952_ (.A(_05225_),
    .B(_05237_),
    .X(_05238_));
 sky130_fd_sc_hd__xnor2_1 _24953_ (.A(_05223_),
    .B(_05238_),
    .Y(_05239_));
 sky130_fd_sc_hd__xnor2_1 _24954_ (.A(_05213_),
    .B(_05239_),
    .Y(_05240_));
 sky130_fd_sc_hd__maj3_1 _24955_ (.A(_05100_),
    .B(_05112_),
    .C(_05114_),
    .X(_05241_));
 sky130_fd_sc_hd__xnor2_1 _24956_ (.A(_05240_),
    .B(_05241_),
    .Y(_05242_));
 sky130_fd_sc_hd__xnor2_2 _24957_ (.A(_05200_),
    .B(_05242_),
    .Y(_05243_));
 sky130_fd_sc_hd__nand2_1 _24958_ (.A(_05145_),
    .B(_05147_),
    .Y(_05244_));
 sky130_fd_sc_hd__nor2_1 _24959_ (.A(_05145_),
    .B(_05147_),
    .Y(_05245_));
 sky130_fd_sc_hd__a21oi_2 _24960_ (.A1(_05091_),
    .A2(_05244_),
    .B1(_05245_),
    .Y(_05246_));
 sky130_fd_sc_hd__xnor2_1 _24961_ (.A(_05243_),
    .B(_05246_),
    .Y(_05247_));
 sky130_fd_sc_hd__xnor2_4 _24962_ (.A(_05199_),
    .B(_05247_),
    .Y(_05248_));
 sky130_fd_sc_hd__nor2_4 _24963_ (.A(_01698_),
    .B(_05248_),
    .Y(_05249_));
 sky130_fd_sc_hd__and2_0 _24964_ (.A(_01698_),
    .B(_03343_),
    .X(_05250_));
 sky130_fd_sc_hd__a21oi_1 _24965_ (.A1(net443),
    .A2(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[63] ),
    .B1(_02646_),
    .Y(_05251_));
 sky130_fd_sc_hd__o31a_4 _24966_ (.A1(net441),
    .A2(_05249_),
    .A3(_05250_),
    .B1(_05251_),
    .X(_05252_));
 sky130_fd_sc_hd__nor2_1 _24967_ (.A(_01733_),
    .B(_01770_),
    .Y(_05253_));
 sky130_fd_sc_hd__a21oi_1 _24968_ (.A1(_01733_),
    .A2(_01882_),
    .B1(_05253_),
    .Y(_05254_));
 sky130_fd_sc_hd__nor2_1 _24969_ (.A(_10724_),
    .B(_01898_),
    .Y(_05255_));
 sky130_fd_sc_hd__a22oi_1 _24970_ (.A1(_10724_),
    .A2(_01896_),
    .B1(_05255_),
    .B2(_10695_),
    .Y(_05256_));
 sky130_fd_sc_hd__nor2_1 _24971_ (.A(_10724_),
    .B(_01903_),
    .Y(_05257_));
 sky130_fd_sc_hd__o22ai_2 _24972_ (.A1(_01893_),
    .A2(_05256_),
    .B1(_05257_),
    .B2(_10695_),
    .Y(_05258_));
 sky130_fd_sc_hd__o221ai_4 _24973_ (.A1(net793),
    .A2(_01889_),
    .B1(_05254_),
    .B2(_01761_),
    .C1(_05258_),
    .Y(_05259_));
 sky130_fd_sc_hd__nand2_2 _24974_ (.A(net739),
    .B(_05259_),
    .Y(_05260_));
 sky130_fd_sc_hd__o211ai_4 _24975_ (.A1(_05193_),
    .A2(_05252_),
    .B1(_05260_),
    .C1(_11824_),
    .Y(_05261_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_245 ();
 sky130_fd_sc_hd__mux4_2 _24977_ (.A0(net51),
    .A1(net33),
    .A2(net56),
    .A3(net42),
    .S0(\load_store_unit_i.rdata_offset_q[1] ),
    .S1(\load_store_unit_i.rdata_offset_q[0] ),
    .X(_05263_));
 sky130_fd_sc_hd__a21oi_4 _24978_ (.A1(_01674_),
    .A2(_05263_),
    .B1(_03479_),
    .Y(_05264_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_244 ();
 sky130_fd_sc_hd__nor2_1 _24980_ (.A(_02123_),
    .B(_05264_),
    .Y(_05266_));
 sky130_fd_sc_hd__a22o_1 _24981_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[159] ),
    .A2(_02123_),
    .B1(_05261_),
    .B2(_05266_),
    .X(_00544_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_243 ();
 sky130_fd_sc_hd__nor3_4 _24983_ (.A(_02117_),
    .B(_01915_),
    .C(net448),
    .Y(_05268_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_242 ();
 sky130_fd_sc_hd__nand2_1 _24985_ (.A(_01909_),
    .B(net1479),
    .Y(_05270_));
 sky130_fd_sc_hd__nor2_8 _24986_ (.A(net448),
    .B(_01915_),
    .Y(_05271_));
 sky130_fd_sc_hd__nand2_8 _24987_ (.A(_02122_),
    .B(_05271_),
    .Y(_05272_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_241 ();
 sky130_fd_sc_hd__nand2_1 _24989_ (.A(\gen_regfile_ff.register_file_i.rf_reg[160] ),
    .B(_05272_),
    .Y(_05274_));
 sky130_fd_sc_hd__nand2_1 _24990_ (.A(_05270_),
    .B(_05274_),
    .Y(_00545_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_240 ();
 sky130_fd_sc_hd__and3_1 _24992_ (.A(_01670_),
    .B(\load_store_unit_i.rdata_offset_q[1] ),
    .C(net35),
    .X(_05276_));
 sky130_fd_sc_hd__a211oi_2 _24993_ (.A1(net58),
    .A2(_01672_),
    .B1(_01674_),
    .C1(_05276_),
    .Y(_05277_));
 sky130_fd_sc_hd__a221oi_2 _24994_ (.A1(\load_store_unit_i.rdata_q[9] ),
    .A2(_01672_),
    .B1(_01683_),
    .B2(\load_store_unit_i.rdata_q[17] ),
    .C1(_01684_),
    .Y(_05278_));
 sky130_fd_sc_hd__a22oi_2 _24995_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(net44),
    .B1(_01688_),
    .B2(\load_store_unit_i.rdata_q[25] ),
    .Y(_05279_));
 sky130_fd_sc_hd__nand3_1 _24996_ (.A(_01670_),
    .B(_01682_),
    .C(net38),
    .Y(_05280_));
 sky130_fd_sc_hd__o221ai_4 _24997_ (.A1(_05277_),
    .A2(_05278_),
    .B1(_05279_),
    .B2(_01693_),
    .C1(_05280_),
    .Y(_05281_));
 sky130_fd_sc_hd__nand2_1 _24998_ (.A(_01700_),
    .B(_03494_),
    .Y(_05282_));
 sky130_fd_sc_hd__o21ai_1 _24999_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[33] ),
    .A2(_01700_),
    .B1(_05282_),
    .Y(_05283_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_239 ();
 sky130_fd_sc_hd__nand2_1 _25001_ (.A(net295),
    .B(_05181_),
    .Y(_05285_));
 sky130_fd_sc_hd__nand2_1 _25002_ (.A(_01773_),
    .B(_05179_),
    .Y(_05286_));
 sky130_fd_sc_hd__a21oi_1 _25003_ (.A1(_05285_),
    .A2(_05286_),
    .B1(_01761_),
    .Y(_05287_));
 sky130_fd_sc_hd__nand2_1 _25004_ (.A(_08999_),
    .B(_02233_),
    .Y(_05288_));
 sky130_fd_sc_hd__nor2_1 _25005_ (.A(_09044_),
    .B(_01898_),
    .Y(_05289_));
 sky130_fd_sc_hd__nor2_1 _25006_ (.A(_08999_),
    .B(_01902_),
    .Y(_05290_));
 sky130_fd_sc_hd__a21oi_1 _25007_ (.A1(net722),
    .A2(_05289_),
    .B1(_05290_),
    .Y(_05291_));
 sky130_fd_sc_hd__nor2_1 _25008_ (.A(_01893_),
    .B(_05291_),
    .Y(_05292_));
 sky130_fd_sc_hd__a21oi_1 _25009_ (.A1(_09044_),
    .A2(_05288_),
    .B1(_05292_),
    .Y(_05293_));
 sky130_fd_sc_hd__a2111oi_0 _25010_ (.A1(_10970_),
    .A2(_01929_),
    .B1(_05287_),
    .C1(_05293_),
    .D1(net314),
    .Y(_05294_));
 sky130_fd_sc_hd__a21oi_1 _25011_ (.A1(_08272_),
    .A2(_05283_),
    .B1(_05294_),
    .Y(_05295_));
 sky130_fd_sc_hd__nand2_1 _25012_ (.A(_08632_),
    .B(_11580_),
    .Y(_05296_));
 sky130_fd_sc_hd__o21ai_0 _25013_ (.A1(_08632_),
    .A2(_05295_),
    .B1(_05296_),
    .Y(_05297_));
 sky130_fd_sc_hd__nand2_1 _25014_ (.A(net265),
    .B(_05297_),
    .Y(_05298_));
 sky130_fd_sc_hd__o21ai_4 _25015_ (.A1(net265),
    .A2(_05281_),
    .B1(_05298_),
    .Y(_05299_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_238 ();
 sky130_fd_sc_hd__nand2_1 _25017_ (.A(\gen_regfile_ff.register_file_i.rf_reg[161] ),
    .B(_05272_),
    .Y(_05301_));
 sky130_fd_sc_hd__o21ai_0 _25018_ (.A1(_05272_),
    .A2(_05299_),
    .B1(_05301_),
    .Y(_00546_));
 sky130_fd_sc_hd__nand2_1 _25019_ (.A(_01916_),
    .B(_02974_),
    .Y(_05302_));
 sky130_fd_sc_hd__nand2_1 _25020_ (.A(\gen_regfile_ff.register_file_i.rf_reg[44] ),
    .B(_01921_),
    .Y(_05303_));
 sky130_fd_sc_hd__nand2_1 _25021_ (.A(_05302_),
    .B(_05303_),
    .Y(_00547_));
 sky130_fd_sc_hd__or2_0 _25022_ (.A(_02284_),
    .B(_03619_),
    .X(_05304_));
 sky130_fd_sc_hd__o21ai_2 _25023_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[34] ),
    .A2(_01700_),
    .B1(_05304_),
    .Y(_05305_));
 sky130_fd_sc_hd__nand2_1 _25024_ (.A(net295),
    .B(_05073_),
    .Y(_05306_));
 sky130_fd_sc_hd__nand2_1 _25025_ (.A(_01773_),
    .B(_05071_),
    .Y(_05307_));
 sky130_fd_sc_hd__a21oi_1 _25026_ (.A1(_05306_),
    .A2(_05307_),
    .B1(_01761_),
    .Y(_05308_));
 sky130_fd_sc_hd__nor3_1 _25027_ (.A(net709),
    .B(_08850_),
    .C(_01898_),
    .Y(_05309_));
 sky130_fd_sc_hd__a21oi_1 _25028_ (.A1(_08850_),
    .A2(_01896_),
    .B1(_05309_),
    .Y(_05310_));
 sky130_fd_sc_hd__o21ai_0 _25029_ (.A1(_08850_),
    .A2(_01903_),
    .B1(net708),
    .Y(_05311_));
 sky130_fd_sc_hd__o21ai_0 _25030_ (.A1(_01893_),
    .A2(_05310_),
    .B1(_05311_),
    .Y(_05312_));
 sky130_fd_sc_hd__o21ai_0 _25031_ (.A1(_10974_),
    .A2(_01889_),
    .B1(_05312_),
    .Y(_05313_));
 sky130_fd_sc_hd__nor3_1 _25032_ (.A(net313),
    .B(_05308_),
    .C(_05313_),
    .Y(_05314_));
 sky130_fd_sc_hd__a21oi_1 _25033_ (.A1(_08272_),
    .A2(_05305_),
    .B1(_05314_),
    .Y(_05315_));
 sky130_fd_sc_hd__nand2_1 _25034_ (.A(_08632_),
    .B(_11307_),
    .Y(_05316_));
 sky130_fd_sc_hd__o21ai_1 _25035_ (.A1(_08632_),
    .A2(_05315_),
    .B1(_05316_),
    .Y(_05317_));
 sky130_fd_sc_hd__and3_1 _25036_ (.A(_01670_),
    .B(\load_store_unit_i.rdata_offset_q[1] ),
    .C(net36),
    .X(_05318_));
 sky130_fd_sc_hd__a21oi_1 _25037_ (.A1(net28),
    .A2(_01672_),
    .B1(_05318_),
    .Y(_05319_));
 sky130_fd_sc_hd__a221oi_1 _25038_ (.A1(\load_store_unit_i.rdata_q[10] ),
    .A2(_01672_),
    .B1(_01683_),
    .B2(\load_store_unit_i.rdata_q[18] ),
    .C1(_01684_),
    .Y(_05320_));
 sky130_fd_sc_hd__a21oi_1 _25039_ (.A1(_01684_),
    .A2(_05319_),
    .B1(_05320_),
    .Y(_05321_));
 sky130_fd_sc_hd__a22oi_1 _25040_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(net45),
    .B1(_01688_),
    .B2(\load_store_unit_i.rdata_q[26] ),
    .Y(_05322_));
 sky130_fd_sc_hd__nor2_1 _25041_ (.A(_01693_),
    .B(_05322_),
    .Y(_05323_));
 sky130_fd_sc_hd__a31o_1 _25042_ (.A1(_01670_),
    .A2(_01682_),
    .A3(net49),
    .B1(_05323_),
    .X(_05324_));
 sky130_fd_sc_hd__nor3_2 _25043_ (.A(net266),
    .B(_05321_),
    .C(_05324_),
    .Y(_05325_));
 sky130_fd_sc_hd__a21oi_4 _25044_ (.A1(net266),
    .A2(_05317_),
    .B1(_05325_),
    .Y(_05326_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_237 ();
 sky130_fd_sc_hd__nand2_1 _25046_ (.A(net1478),
    .B(_05326_),
    .Y(_05328_));
 sky130_fd_sc_hd__nand2_1 _25047_ (.A(\gen_regfile_ff.register_file_i.rf_reg[162] ),
    .B(_05272_),
    .Y(_05329_));
 sky130_fd_sc_hd__nand2_1 _25048_ (.A(_05328_),
    .B(_05329_),
    .Y(_00548_));
 sky130_fd_sc_hd__and3_1 _25049_ (.A(_01670_),
    .B(\load_store_unit_i.rdata_offset_q[1] ),
    .C(net37),
    .X(_05330_));
 sky130_fd_sc_hd__a211oi_2 _25050_ (.A1(net29),
    .A2(_01672_),
    .B1(_01674_),
    .C1(_05330_),
    .Y(_05331_));
 sky130_fd_sc_hd__a221oi_2 _25051_ (.A1(\load_store_unit_i.rdata_q[11] ),
    .A2(_01672_),
    .B1(_01683_),
    .B2(\load_store_unit_i.rdata_q[19] ),
    .C1(_01684_),
    .Y(_05332_));
 sky130_fd_sc_hd__a22oi_2 _25052_ (.A1(\load_store_unit_i.data_type_q[1] ),
    .A2(net46),
    .B1(_01688_),
    .B2(\load_store_unit_i.rdata_q[27] ),
    .Y(_05333_));
 sky130_fd_sc_hd__nand3_1 _25053_ (.A(_01670_),
    .B(_01682_),
    .C(net52),
    .Y(_05334_));
 sky130_fd_sc_hd__o221ai_4 _25054_ (.A1(_05331_),
    .A2(_05332_),
    .B1(_05333_),
    .B2(_01693_),
    .C1(_05334_),
    .Y(_05335_));
 sky130_fd_sc_hd__nand2_1 _25055_ (.A(_01762_),
    .B(_04885_),
    .Y(_05336_));
 sky130_fd_sc_hd__nand2_1 _25056_ (.A(_01773_),
    .B(_04882_),
    .Y(_05337_));
 sky130_fd_sc_hd__a21oi_2 _25057_ (.A1(_05336_),
    .A2(_05337_),
    .B1(_01761_),
    .Y(_05338_));
 sky130_fd_sc_hd__nand2_1 _25058_ (.A(net1131),
    .B(_02233_),
    .Y(_05339_));
 sky130_fd_sc_hd__nor2_1 _25059_ (.A(_08636_),
    .B(_01898_),
    .Y(_05340_));
 sky130_fd_sc_hd__nor2_1 _25060_ (.A(_08694_),
    .B(_01902_),
    .Y(_05341_));
 sky130_fd_sc_hd__a21oi_1 _25061_ (.A1(_08694_),
    .A2(_05340_),
    .B1(_05341_),
    .Y(_05342_));
 sky130_fd_sc_hd__nor2_1 _25062_ (.A(_01893_),
    .B(_05342_),
    .Y(_05343_));
 sky130_fd_sc_hd__a21oi_1 _25063_ (.A1(_08636_),
    .A2(_05339_),
    .B1(_05343_),
    .Y(_05344_));
 sky130_fd_sc_hd__a211oi_1 _25064_ (.A1(net174),
    .A2(_01929_),
    .B1(_05338_),
    .C1(_05344_),
    .Y(_05345_));
 sky130_fd_sc_hd__nand2_1 _25065_ (.A(_01700_),
    .B(_03751_),
    .Y(_05346_));
 sky130_fd_sc_hd__o211ai_4 _25066_ (.A1(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[35] ),
    .A2(_01700_),
    .B1(_05346_),
    .C1(net312),
    .Y(_05347_));
 sky130_fd_sc_hd__o211ai_1 _25067_ (.A1(net1101),
    .A2(_05345_),
    .B1(_05347_),
    .C1(_08581_),
    .Y(_05348_));
 sky130_fd_sc_hd__o21ai_0 _25068_ (.A1(_08581_),
    .A2(_11864_),
    .B1(_05348_),
    .Y(_05349_));
 sky130_fd_sc_hd__nand2_1 _25069_ (.A(net266),
    .B(_05349_),
    .Y(_05350_));
 sky130_fd_sc_hd__o21ai_4 _25070_ (.A1(net266),
    .A2(_05335_),
    .B1(_05350_),
    .Y(_05351_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_236 ();
 sky130_fd_sc_hd__nand2_1 _25072_ (.A(\gen_regfile_ff.register_file_i.rf_reg[163] ),
    .B(_05272_),
    .Y(_05353_));
 sky130_fd_sc_hd__o21ai_0 _25073_ (.A1(_05272_),
    .A2(_05351_),
    .B1(_05353_),
    .Y(_00549_));
 sky130_fd_sc_hd__nand2_1 _25074_ (.A(_02113_),
    .B(net257),
    .Y(_05354_));
 sky130_fd_sc_hd__nand2_1 _25075_ (.A(\gen_regfile_ff.register_file_i.rf_reg[164] ),
    .B(_05272_),
    .Y(_05355_));
 sky130_fd_sc_hd__nand2_1 _25076_ (.A(_05354_),
    .B(_05355_),
    .Y(_00550_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_235 ();
 sky130_fd_sc_hd__nand2_1 _25078_ (.A(_02250_),
    .B(net257),
    .Y(_05357_));
 sky130_fd_sc_hd__nand2_1 _25079_ (.A(\gen_regfile_ff.register_file_i.rf_reg[165] ),
    .B(_05272_),
    .Y(_05358_));
 sky130_fd_sc_hd__nand2_1 _25080_ (.A(_05357_),
    .B(_05358_),
    .Y(_00551_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_234 ();
 sky130_fd_sc_hd__nand2_1 _25082_ (.A(_02360_),
    .B(net257),
    .Y(_05360_));
 sky130_fd_sc_hd__nand2_1 _25083_ (.A(\gen_regfile_ff.register_file_i.rf_reg[166] ),
    .B(_05272_),
    .Y(_05361_));
 sky130_fd_sc_hd__nand2_1 _25084_ (.A(_05360_),
    .B(_05361_),
    .Y(_00552_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_233 ();
 sky130_fd_sc_hd__nand2_1 _25086_ (.A(_02468_),
    .B(net257),
    .Y(_05363_));
 sky130_fd_sc_hd__nand2_1 _25087_ (.A(\gen_regfile_ff.register_file_i.rf_reg[167] ),
    .B(_05272_),
    .Y(_05364_));
 sky130_fd_sc_hd__nand2_1 _25088_ (.A(_05363_),
    .B(_05364_),
    .Y(_00553_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_232 ();
 sky130_fd_sc_hd__nand2_1 _25090_ (.A(_02553_),
    .B(net1478),
    .Y(_05366_));
 sky130_fd_sc_hd__nand2_1 _25091_ (.A(\gen_regfile_ff.register_file_i.rf_reg[168] ),
    .B(_05272_),
    .Y(_05367_));
 sky130_fd_sc_hd__nand2_1 _25092_ (.A(_05366_),
    .B(_05367_),
    .Y(_00554_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_231 ();
 sky130_fd_sc_hd__nand2_1 _25094_ (.A(_02653_),
    .B(net1479),
    .Y(_05369_));
 sky130_fd_sc_hd__nand2_1 _25095_ (.A(\gen_regfile_ff.register_file_i.rf_reg[169] ),
    .B(_05272_),
    .Y(_05370_));
 sky130_fd_sc_hd__nand2_1 _25096_ (.A(_05369_),
    .B(_05370_),
    .Y(_00555_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_230 ();
 sky130_fd_sc_hd__nand2_1 _25098_ (.A(_02761_),
    .B(net257),
    .Y(_05372_));
 sky130_fd_sc_hd__nand2_1 _25099_ (.A(\gen_regfile_ff.register_file_i.rf_reg[170] ),
    .B(_05272_),
    .Y(_05373_));
 sky130_fd_sc_hd__nand2_1 _25100_ (.A(_05372_),
    .B(_05373_),
    .Y(_00556_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_229 ();
 sky130_fd_sc_hd__nand2_1 _25102_ (.A(_02849_),
    .B(net257),
    .Y(_05375_));
 sky130_fd_sc_hd__nand2_1 _25103_ (.A(\gen_regfile_ff.register_file_i.rf_reg[171] ),
    .B(_05272_),
    .Y(_05376_));
 sky130_fd_sc_hd__nand2_1 _25104_ (.A(_05375_),
    .B(_05376_),
    .Y(_00557_));
 sky130_fd_sc_hd__nand2_1 _25105_ (.A(_01916_),
    .B(_03080_),
    .Y(_05377_));
 sky130_fd_sc_hd__nand2_1 _25106_ (.A(\gen_regfile_ff.register_file_i.rf_reg[45] ),
    .B(_01921_),
    .Y(_05378_));
 sky130_fd_sc_hd__nand2_1 _25107_ (.A(_05377_),
    .B(_05378_),
    .Y(_00558_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_227 ();
 sky130_fd_sc_hd__nand2_1 _25110_ (.A(_02974_),
    .B(net257),
    .Y(_05381_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_226 ();
 sky130_fd_sc_hd__nand2_1 _25112_ (.A(\gen_regfile_ff.register_file_i.rf_reg[172] ),
    .B(_05272_),
    .Y(_05383_));
 sky130_fd_sc_hd__nand2_1 _25113_ (.A(_05381_),
    .B(_05383_),
    .Y(_00559_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_225 ();
 sky130_fd_sc_hd__nand2_1 _25115_ (.A(_03080_),
    .B(net1479),
    .Y(_05385_));
 sky130_fd_sc_hd__nand2_1 _25116_ (.A(\gen_regfile_ff.register_file_i.rf_reg[173] ),
    .B(_05272_),
    .Y(_05386_));
 sky130_fd_sc_hd__nand2_1 _25117_ (.A(_05385_),
    .B(_05386_),
    .Y(_00560_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_224 ();
 sky130_fd_sc_hd__nand2_1 _25119_ (.A(_03214_),
    .B(net257),
    .Y(_05388_));
 sky130_fd_sc_hd__nand2_1 _25120_ (.A(\gen_regfile_ff.register_file_i.rf_reg[174] ),
    .B(_05272_),
    .Y(_05389_));
 sky130_fd_sc_hd__nand2_1 _25121_ (.A(_05388_),
    .B(_05389_),
    .Y(_00561_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_223 ();
 sky130_fd_sc_hd__nand2_1 _25123_ (.A(_03348_),
    .B(net1479),
    .Y(_05391_));
 sky130_fd_sc_hd__nand2_1 _25124_ (.A(\gen_regfile_ff.register_file_i.rf_reg[175] ),
    .B(_05272_),
    .Y(_05392_));
 sky130_fd_sc_hd__nand2_1 _25125_ (.A(_05391_),
    .B(_05392_),
    .Y(_00562_));
 sky130_fd_sc_hd__nand2_1 _25126_ (.A(\gen_regfile_ff.register_file_i.rf_reg[176] ),
    .B(_05272_),
    .Y(_05393_));
 sky130_fd_sc_hd__o21ai_0 _25127_ (.A1(_03481_),
    .A2(_05272_),
    .B1(_05393_),
    .Y(_00563_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_222 ();
 sky130_fd_sc_hd__nand2_1 _25129_ (.A(_03614_),
    .B(net1479),
    .Y(_05395_));
 sky130_fd_sc_hd__nand2_1 _25130_ (.A(\gen_regfile_ff.register_file_i.rf_reg[177] ),
    .B(_05272_),
    .Y(_05396_));
 sky130_fd_sc_hd__nand2_1 _25131_ (.A(_05395_),
    .B(_05396_),
    .Y(_00564_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_221 ();
 sky130_fd_sc_hd__nand2_1 _25133_ (.A(_03739_),
    .B(net1478),
    .Y(_05398_));
 sky130_fd_sc_hd__nand2_1 _25134_ (.A(\gen_regfile_ff.register_file_i.rf_reg[178] ),
    .B(_05272_),
    .Y(_05399_));
 sky130_fd_sc_hd__nand2_1 _25135_ (.A(_05398_),
    .B(_05399_),
    .Y(_00565_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_220 ();
 sky130_fd_sc_hd__nand2_1 _25137_ (.A(_03866_),
    .B(net1478),
    .Y(_05401_));
 sky130_fd_sc_hd__nand2_1 _25138_ (.A(\gen_regfile_ff.register_file_i.rf_reg[179] ),
    .B(_05272_),
    .Y(_05402_));
 sky130_fd_sc_hd__nand2_1 _25139_ (.A(_05401_),
    .B(_05402_),
    .Y(_00566_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_219 ();
 sky130_fd_sc_hd__nand2_1 _25141_ (.A(net1544),
    .B(net257),
    .Y(_05404_));
 sky130_fd_sc_hd__nand2_1 _25142_ (.A(\gen_regfile_ff.register_file_i.rf_reg[180] ),
    .B(_05272_),
    .Y(_05405_));
 sky130_fd_sc_hd__nand2_1 _25143_ (.A(_05404_),
    .B(_05405_),
    .Y(_00567_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_218 ();
 sky130_fd_sc_hd__nand2_1 _25145_ (.A(net1585),
    .B(net257),
    .Y(_05407_));
 sky130_fd_sc_hd__nand2_1 _25146_ (.A(\gen_regfile_ff.register_file_i.rf_reg[181] ),
    .B(_05272_),
    .Y(_05408_));
 sky130_fd_sc_hd__nand2_1 _25147_ (.A(_05407_),
    .B(_05408_),
    .Y(_00568_));
 sky130_fd_sc_hd__nand2_1 _25148_ (.A(_01916_),
    .B(_03214_),
    .Y(_05409_));
 sky130_fd_sc_hd__nand2_1 _25149_ (.A(\gen_regfile_ff.register_file_i.rf_reg[46] ),
    .B(_01921_),
    .Y(_05410_));
 sky130_fd_sc_hd__nand2_1 _25150_ (.A(_05409_),
    .B(_05410_),
    .Y(_00569_));
 sky130_fd_sc_hd__mux2_4 _25151_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[182] ),
    .A1(_04252_),
    .S(net257),
    .X(_00570_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_217 ();
 sky130_fd_sc_hd__nand2_1 _25153_ (.A(_04390_),
    .B(net257),
    .Y(_05412_));
 sky130_fd_sc_hd__nand2_1 _25154_ (.A(\gen_regfile_ff.register_file_i.rf_reg[183] ),
    .B(_05272_),
    .Y(_05413_));
 sky130_fd_sc_hd__nand2_1 _25155_ (.A(_05412_),
    .B(_05413_),
    .Y(_00571_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_216 ();
 sky130_fd_sc_hd__nand2_2 _25157_ (.A(net1270),
    .B(net257),
    .Y(_05415_));
 sky130_fd_sc_hd__nand2_1 _25158_ (.A(\gen_regfile_ff.register_file_i.rf_reg[184] ),
    .B(_05272_),
    .Y(_05416_));
 sky130_fd_sc_hd__nand2_1 _25159_ (.A(_05415_),
    .B(_05416_),
    .Y(_00572_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_215 ();
 sky130_fd_sc_hd__nand2_1 _25161_ (.A(_04661_),
    .B(net1479),
    .Y(_05418_));
 sky130_fd_sc_hd__nand2_1 _25162_ (.A(\gen_regfile_ff.register_file_i.rf_reg[185] ),
    .B(_05272_),
    .Y(_05419_));
 sky130_fd_sc_hd__nand2_1 _25163_ (.A(_05418_),
    .B(_05419_),
    .Y(_00573_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_214 ();
 sky130_fd_sc_hd__nand2_2 _25165_ (.A(net1514),
    .B(net257),
    .Y(_05421_));
 sky130_fd_sc_hd__nand2_1 _25166_ (.A(\gen_regfile_ff.register_file_i.rf_reg[186] ),
    .B(_05272_),
    .Y(_05422_));
 sky130_fd_sc_hd__nand2_1 _25167_ (.A(_05421_),
    .B(_05422_),
    .Y(_00574_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_213 ();
 sky130_fd_sc_hd__nand2_4 _25169_ (.A(net1540),
    .B(net257),
    .Y(_05424_));
 sky130_fd_sc_hd__nand2_1 _25170_ (.A(\gen_regfile_ff.register_file_i.rf_reg[187] ),
    .B(_05272_),
    .Y(_05425_));
 sky130_fd_sc_hd__nand2_2 _25171_ (.A(_05424_),
    .B(_05425_),
    .Y(_00575_));
 sky130_fd_sc_hd__mux2_4 _25172_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[188] ),
    .A1(_04975_),
    .S(net257),
    .X(_00576_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_212 ();
 sky130_fd_sc_hd__nor2_1 _25174_ (.A(_05084_),
    .B(_05272_),
    .Y(_05427_));
 sky130_fd_sc_hd__a22o_1 _25175_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[189] ),
    .A2(_05272_),
    .B1(_05079_),
    .B2(_05427_),
    .X(_00577_));
 sky130_fd_sc_hd__mux2_4 _25176_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[190] ),
    .A1(_05191_),
    .S(net1477),
    .X(_00578_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_211 ();
 sky130_fd_sc_hd__nor2_1 _25178_ (.A(_05264_),
    .B(_05272_),
    .Y(_05429_));
 sky130_fd_sc_hd__a22o_1 _25179_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[191] ),
    .A2(_05272_),
    .B1(_05429_),
    .B2(_05261_),
    .X(_00579_));
 sky130_fd_sc_hd__nand2_1 _25180_ (.A(_01916_),
    .B(_03348_),
    .Y(_05430_));
 sky130_fd_sc_hd__nand2_1 _25181_ (.A(\gen_regfile_ff.register_file_i.rf_reg[47] ),
    .B(_01921_),
    .Y(_05431_));
 sky130_fd_sc_hd__nand2_1 _25182_ (.A(_05430_),
    .B(_05431_),
    .Y(_00580_));
 sky130_fd_sc_hd__nand2b_4 _25183_ (.A_N(net331),
    .B(net1021),
    .Y(_05432_));
 sky130_fd_sc_hd__nor3_4 _25184_ (.A(net447),
    .B(_02117_),
    .C(_05432_),
    .Y(_05433_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_210 ();
 sky130_fd_sc_hd__nand2_1 _25186_ (.A(_01909_),
    .B(_05433_),
    .Y(_05435_));
 sky130_fd_sc_hd__nor2_8 _25187_ (.A(net447),
    .B(_05432_),
    .Y(_05436_));
 sky130_fd_sc_hd__nand2_8 _25188_ (.A(_02122_),
    .B(_05436_),
    .Y(_05437_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_209 ();
 sky130_fd_sc_hd__nand2_1 _25190_ (.A(\gen_regfile_ff.register_file_i.rf_reg[192] ),
    .B(_05437_),
    .Y(_05439_));
 sky130_fd_sc_hd__nand2_1 _25191_ (.A(_05435_),
    .B(_05439_),
    .Y(_00581_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_208 ();
 sky130_fd_sc_hd__nand2_1 _25193_ (.A(\gen_regfile_ff.register_file_i.rf_reg[193] ),
    .B(_05437_),
    .Y(_05441_));
 sky130_fd_sc_hd__o21ai_0 _25194_ (.A1(_05299_),
    .A2(_05437_),
    .B1(_05441_),
    .Y(_00582_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_207 ();
 sky130_fd_sc_hd__nand2_1 _25196_ (.A(_05326_),
    .B(_05433_),
    .Y(_05443_));
 sky130_fd_sc_hd__nand2_1 _25197_ (.A(\gen_regfile_ff.register_file_i.rf_reg[194] ),
    .B(_05437_),
    .Y(_05444_));
 sky130_fd_sc_hd__nand2_1 _25198_ (.A(_05443_),
    .B(_05444_),
    .Y(_00583_));
 sky130_fd_sc_hd__nand2_1 _25199_ (.A(\gen_regfile_ff.register_file_i.rf_reg[195] ),
    .B(_05437_),
    .Y(_05445_));
 sky130_fd_sc_hd__o21ai_0 _25200_ (.A1(_05351_),
    .A2(_05437_),
    .B1(_05445_),
    .Y(_00584_));
 sky130_fd_sc_hd__nand2_1 _25201_ (.A(_02113_),
    .B(net256),
    .Y(_05446_));
 sky130_fd_sc_hd__nand2_1 _25202_ (.A(\gen_regfile_ff.register_file_i.rf_reg[196] ),
    .B(_05437_),
    .Y(_05447_));
 sky130_fd_sc_hd__nand2_1 _25203_ (.A(_05446_),
    .B(_05447_),
    .Y(_00585_));
 sky130_fd_sc_hd__nand2_1 _25204_ (.A(_02250_),
    .B(net256),
    .Y(_05448_));
 sky130_fd_sc_hd__nand2_1 _25205_ (.A(\gen_regfile_ff.register_file_i.rf_reg[197] ),
    .B(_05437_),
    .Y(_05449_));
 sky130_fd_sc_hd__nand2_1 _25206_ (.A(_05448_),
    .B(_05449_),
    .Y(_00586_));
 sky130_fd_sc_hd__nand2_1 _25207_ (.A(_02360_),
    .B(net256),
    .Y(_05450_));
 sky130_fd_sc_hd__nand2_1 _25208_ (.A(\gen_regfile_ff.register_file_i.rf_reg[198] ),
    .B(_05437_),
    .Y(_05451_));
 sky130_fd_sc_hd__nand2_1 _25209_ (.A(_05450_),
    .B(_05451_),
    .Y(_00587_));
 sky130_fd_sc_hd__nand2_1 _25210_ (.A(_02468_),
    .B(net256),
    .Y(_05452_));
 sky130_fd_sc_hd__nand2_1 _25211_ (.A(\gen_regfile_ff.register_file_i.rf_reg[199] ),
    .B(_05437_),
    .Y(_05453_));
 sky130_fd_sc_hd__nand2_1 _25212_ (.A(_05452_),
    .B(_05453_),
    .Y(_00588_));
 sky130_fd_sc_hd__nand2_1 _25213_ (.A(_02553_),
    .B(_05433_),
    .Y(_05454_));
 sky130_fd_sc_hd__nand2_1 _25214_ (.A(\gen_regfile_ff.register_file_i.rf_reg[200] ),
    .B(_05437_),
    .Y(_05455_));
 sky130_fd_sc_hd__nand2_1 _25215_ (.A(_05454_),
    .B(_05455_),
    .Y(_00589_));
 sky130_fd_sc_hd__nand2_1 _25216_ (.A(_02653_),
    .B(net256),
    .Y(_05456_));
 sky130_fd_sc_hd__nand2_1 _25217_ (.A(\gen_regfile_ff.register_file_i.rf_reg[201] ),
    .B(_05437_),
    .Y(_05457_));
 sky130_fd_sc_hd__nand2_1 _25218_ (.A(_05456_),
    .B(_05457_),
    .Y(_00590_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_206 ();
 sky130_fd_sc_hd__nand2_1 _25220_ (.A(\gen_regfile_ff.register_file_i.rf_reg[48] ),
    .B(_01921_),
    .Y(_05459_));
 sky130_fd_sc_hd__o21ai_0 _25221_ (.A1(_01921_),
    .A2(_03481_),
    .B1(_05459_),
    .Y(_00591_));
 sky130_fd_sc_hd__nand2_1 _25222_ (.A(_02761_),
    .B(net256),
    .Y(_05460_));
 sky130_fd_sc_hd__nand2_1 _25223_ (.A(\gen_regfile_ff.register_file_i.rf_reg[202] ),
    .B(_05437_),
    .Y(_05461_));
 sky130_fd_sc_hd__nand2_1 _25224_ (.A(_05460_),
    .B(_05461_),
    .Y(_00592_));
 sky130_fd_sc_hd__nand2_1 _25225_ (.A(_02849_),
    .B(net256),
    .Y(_05462_));
 sky130_fd_sc_hd__nand2_1 _25226_ (.A(\gen_regfile_ff.register_file_i.rf_reg[203] ),
    .B(_05437_),
    .Y(_05463_));
 sky130_fd_sc_hd__nand2_1 _25227_ (.A(_05462_),
    .B(_05463_),
    .Y(_00593_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_205 ();
 sky130_fd_sc_hd__nand2_1 _25229_ (.A(_02974_),
    .B(net256),
    .Y(_05465_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_204 ();
 sky130_fd_sc_hd__nand2_1 _25231_ (.A(\gen_regfile_ff.register_file_i.rf_reg[204] ),
    .B(_05437_),
    .Y(_05467_));
 sky130_fd_sc_hd__nand2_1 _25232_ (.A(_05465_),
    .B(_05467_),
    .Y(_00594_));
 sky130_fd_sc_hd__nand2_1 _25233_ (.A(_03080_),
    .B(_05433_),
    .Y(_05468_));
 sky130_fd_sc_hd__nand2_1 _25234_ (.A(\gen_regfile_ff.register_file_i.rf_reg[205] ),
    .B(_05437_),
    .Y(_05469_));
 sky130_fd_sc_hd__nand2_1 _25235_ (.A(_05468_),
    .B(_05469_),
    .Y(_00595_));
 sky130_fd_sc_hd__nand2_1 _25236_ (.A(_03214_),
    .B(net256),
    .Y(_05470_));
 sky130_fd_sc_hd__nand2_1 _25237_ (.A(\gen_regfile_ff.register_file_i.rf_reg[206] ),
    .B(_05437_),
    .Y(_05471_));
 sky130_fd_sc_hd__nand2_1 _25238_ (.A(_05470_),
    .B(_05471_),
    .Y(_00596_));
 sky130_fd_sc_hd__nand2_1 _25239_ (.A(_03348_),
    .B(_05433_),
    .Y(_05472_));
 sky130_fd_sc_hd__nand2_1 _25240_ (.A(\gen_regfile_ff.register_file_i.rf_reg[207] ),
    .B(_05437_),
    .Y(_05473_));
 sky130_fd_sc_hd__nand2_1 _25241_ (.A(_05472_),
    .B(_05473_),
    .Y(_00597_));
 sky130_fd_sc_hd__nand2_1 _25242_ (.A(\gen_regfile_ff.register_file_i.rf_reg[208] ),
    .B(_05437_),
    .Y(_05474_));
 sky130_fd_sc_hd__o21ai_0 _25243_ (.A1(_03481_),
    .A2(_05437_),
    .B1(_05474_),
    .Y(_00598_));
 sky130_fd_sc_hd__nand2_1 _25244_ (.A(_03614_),
    .B(_05433_),
    .Y(_05475_));
 sky130_fd_sc_hd__nand2_1 _25245_ (.A(\gen_regfile_ff.register_file_i.rf_reg[209] ),
    .B(_05437_),
    .Y(_05476_));
 sky130_fd_sc_hd__nand2_1 _25246_ (.A(_05475_),
    .B(_05476_),
    .Y(_00599_));
 sky130_fd_sc_hd__nand2_1 _25247_ (.A(_03739_),
    .B(_05433_),
    .Y(_05477_));
 sky130_fd_sc_hd__nand2_1 _25248_ (.A(\gen_regfile_ff.register_file_i.rf_reg[210] ),
    .B(_05437_),
    .Y(_05478_));
 sky130_fd_sc_hd__nand2_1 _25249_ (.A(_05477_),
    .B(_05478_),
    .Y(_00600_));
 sky130_fd_sc_hd__nand2_1 _25250_ (.A(_03866_),
    .B(_05433_),
    .Y(_05479_));
 sky130_fd_sc_hd__nand2_1 _25251_ (.A(\gen_regfile_ff.register_file_i.rf_reg[211] ),
    .B(_05437_),
    .Y(_05480_));
 sky130_fd_sc_hd__nand2_1 _25252_ (.A(_05479_),
    .B(_05480_),
    .Y(_00601_));
 sky130_fd_sc_hd__nand2_1 _25253_ (.A(_01916_),
    .B(_03614_),
    .Y(_05481_));
 sky130_fd_sc_hd__nand2_1 _25254_ (.A(\gen_regfile_ff.register_file_i.rf_reg[49] ),
    .B(_01921_),
    .Y(_05482_));
 sky130_fd_sc_hd__nand2_1 _25255_ (.A(_05481_),
    .B(_05482_),
    .Y(_00602_));
 sky130_fd_sc_hd__nand2_1 _25256_ (.A(_03982_),
    .B(net256),
    .Y(_05483_));
 sky130_fd_sc_hd__nand2_1 _25257_ (.A(\gen_regfile_ff.register_file_i.rf_reg[212] ),
    .B(_05437_),
    .Y(_05484_));
 sky130_fd_sc_hd__nand2_1 _25258_ (.A(_05483_),
    .B(_05484_),
    .Y(_00603_));
 sky130_fd_sc_hd__nand2_1 _25259_ (.A(net1017),
    .B(net256),
    .Y(_05485_));
 sky130_fd_sc_hd__nand2_1 _25260_ (.A(\gen_regfile_ff.register_file_i.rf_reg[213] ),
    .B(_05437_),
    .Y(_05486_));
 sky130_fd_sc_hd__nand2_1 _25261_ (.A(_05485_),
    .B(_05486_),
    .Y(_00604_));
 sky130_fd_sc_hd__mux2_1 _25262_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[214] ),
    .A1(_04252_),
    .S(net256),
    .X(_00605_));
 sky130_fd_sc_hd__nand2_1 _25263_ (.A(_04390_),
    .B(net256),
    .Y(_05487_));
 sky130_fd_sc_hd__nand2_1 _25264_ (.A(\gen_regfile_ff.register_file_i.rf_reg[215] ),
    .B(_05437_),
    .Y(_05488_));
 sky130_fd_sc_hd__nand2_1 _25265_ (.A(_05487_),
    .B(_05488_),
    .Y(_00606_));
 sky130_fd_sc_hd__nand2_2 _25266_ (.A(net1317),
    .B(net256),
    .Y(_05489_));
 sky130_fd_sc_hd__nand2_1 _25267_ (.A(\gen_regfile_ff.register_file_i.rf_reg[216] ),
    .B(_05437_),
    .Y(_05490_));
 sky130_fd_sc_hd__nand2_1 _25268_ (.A(_05489_),
    .B(_05490_),
    .Y(_00607_));
 sky130_fd_sc_hd__nand2_2 _25269_ (.A(net1564),
    .B(net256),
    .Y(_05491_));
 sky130_fd_sc_hd__nand2_1 _25270_ (.A(\gen_regfile_ff.register_file_i.rf_reg[217] ),
    .B(_05437_),
    .Y(_05492_));
 sky130_fd_sc_hd__nand2_1 _25271_ (.A(_05491_),
    .B(_05492_),
    .Y(_00608_));
 sky130_fd_sc_hd__nand2_1 _25272_ (.A(net1514),
    .B(net256),
    .Y(_05493_));
 sky130_fd_sc_hd__nand2_1 _25273_ (.A(\gen_regfile_ff.register_file_i.rf_reg[218] ),
    .B(_05437_),
    .Y(_05494_));
 sky130_fd_sc_hd__nand2_1 _25274_ (.A(_05493_),
    .B(_05494_),
    .Y(_00609_));
 sky130_fd_sc_hd__nand2_1 _25275_ (.A(net1540),
    .B(net256),
    .Y(_05495_));
 sky130_fd_sc_hd__nand2_1 _25276_ (.A(\gen_regfile_ff.register_file_i.rf_reg[219] ),
    .B(_05437_),
    .Y(_05496_));
 sky130_fd_sc_hd__nand2_1 _25277_ (.A(_05495_),
    .B(_05496_),
    .Y(_00610_));
 sky130_fd_sc_hd__mux2_4 _25278_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[220] ),
    .A1(_04975_),
    .S(net256),
    .X(_00611_));
 sky130_fd_sc_hd__nor2_1 _25279_ (.A(_05084_),
    .B(_05437_),
    .Y(_05497_));
 sky130_fd_sc_hd__a22o_1 _25280_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[221] ),
    .A2(_05437_),
    .B1(_05079_),
    .B2(_05497_),
    .X(_00612_));
 sky130_fd_sc_hd__nand2_1 _25281_ (.A(_01916_),
    .B(_03739_),
    .Y(_05498_));
 sky130_fd_sc_hd__nand2_1 _25282_ (.A(\gen_regfile_ff.register_file_i.rf_reg[50] ),
    .B(_01921_),
    .Y(_05499_));
 sky130_fd_sc_hd__nand2_1 _25283_ (.A(_05498_),
    .B(_05499_),
    .Y(_00613_));
 sky130_fd_sc_hd__mux2_4 _25284_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[222] ),
    .A1(net1237),
    .S(net256),
    .X(_00614_));
 sky130_fd_sc_hd__nor2_1 _25285_ (.A(_05264_),
    .B(_05437_),
    .Y(_05500_));
 sky130_fd_sc_hd__a22o_1 _25286_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[223] ),
    .A2(_05437_),
    .B1(net740),
    .B2(_05500_),
    .X(_00615_));
 sky130_fd_sc_hd__nand2_8 _25287_ (.A(net1021),
    .B(net331),
    .Y(_05501_));
 sky130_fd_sc_hd__nor3_4 _25288_ (.A(net448),
    .B(_02117_),
    .C(_05501_),
    .Y(_05502_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_203 ();
 sky130_fd_sc_hd__nand2_1 _25290_ (.A(_01909_),
    .B(_05502_),
    .Y(_05504_));
 sky130_fd_sc_hd__nor2_8 _25291_ (.A(net447),
    .B(_05501_),
    .Y(_05505_));
 sky130_fd_sc_hd__nand2_8 _25292_ (.A(_02122_),
    .B(_05505_),
    .Y(_05506_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_202 ();
 sky130_fd_sc_hd__nand2_1 _25294_ (.A(\gen_regfile_ff.register_file_i.rf_reg[224] ),
    .B(_05506_),
    .Y(_05508_));
 sky130_fd_sc_hd__nand2_1 _25295_ (.A(_05504_),
    .B(_05508_),
    .Y(_00616_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_201 ();
 sky130_fd_sc_hd__nand2_1 _25297_ (.A(\gen_regfile_ff.register_file_i.rf_reg[225] ),
    .B(_05506_),
    .Y(_05510_));
 sky130_fd_sc_hd__o21ai_0 _25298_ (.A1(_05299_),
    .A2(_05506_),
    .B1(_05510_),
    .Y(_00617_));
 sky130_fd_sc_hd__nand2_1 _25299_ (.A(_05326_),
    .B(_05502_),
    .Y(_05511_));
 sky130_fd_sc_hd__nand2_1 _25300_ (.A(\gen_regfile_ff.register_file_i.rf_reg[226] ),
    .B(_05506_),
    .Y(_05512_));
 sky130_fd_sc_hd__nand2_1 _25301_ (.A(_05511_),
    .B(_05512_),
    .Y(_00618_));
 sky130_fd_sc_hd__nand2_1 _25302_ (.A(\gen_regfile_ff.register_file_i.rf_reg[227] ),
    .B(_05506_),
    .Y(_05513_));
 sky130_fd_sc_hd__o21ai_0 _25303_ (.A1(_05351_),
    .A2(_05506_),
    .B1(_05513_),
    .Y(_00619_));
 sky130_fd_sc_hd__nand2_1 _25304_ (.A(_02113_),
    .B(net255),
    .Y(_05514_));
 sky130_fd_sc_hd__nand2_1 _25305_ (.A(\gen_regfile_ff.register_file_i.rf_reg[228] ),
    .B(_05506_),
    .Y(_05515_));
 sky130_fd_sc_hd__nand2_1 _25306_ (.A(_05514_),
    .B(_05515_),
    .Y(_00620_));
 sky130_fd_sc_hd__nand2_1 _25307_ (.A(_02250_),
    .B(net255),
    .Y(_05516_));
 sky130_fd_sc_hd__nand2_1 _25308_ (.A(\gen_regfile_ff.register_file_i.rf_reg[229] ),
    .B(_05506_),
    .Y(_05517_));
 sky130_fd_sc_hd__nand2_1 _25309_ (.A(_05516_),
    .B(_05517_),
    .Y(_00621_));
 sky130_fd_sc_hd__nand2_1 _25310_ (.A(_02360_),
    .B(net255),
    .Y(_05518_));
 sky130_fd_sc_hd__nand2_1 _25311_ (.A(\gen_regfile_ff.register_file_i.rf_reg[230] ),
    .B(_05506_),
    .Y(_05519_));
 sky130_fd_sc_hd__nand2_1 _25312_ (.A(_05518_),
    .B(_05519_),
    .Y(_00622_));
 sky130_fd_sc_hd__nand2_1 _25313_ (.A(_02468_),
    .B(net255),
    .Y(_05520_));
 sky130_fd_sc_hd__nand2_1 _25314_ (.A(\gen_regfile_ff.register_file_i.rf_reg[231] ),
    .B(_05506_),
    .Y(_05521_));
 sky130_fd_sc_hd__nand2_1 _25315_ (.A(_05520_),
    .B(_05521_),
    .Y(_00623_));
 sky130_fd_sc_hd__nand2_1 _25316_ (.A(_01916_),
    .B(_03866_),
    .Y(_05522_));
 sky130_fd_sc_hd__nand2_1 _25317_ (.A(\gen_regfile_ff.register_file_i.rf_reg[51] ),
    .B(_01921_),
    .Y(_05523_));
 sky130_fd_sc_hd__nand2_1 _25318_ (.A(_05522_),
    .B(_05523_),
    .Y(_00624_));
 sky130_fd_sc_hd__nand2_1 _25319_ (.A(\gen_regfile_ff.register_file_i.rf_reg[33] ),
    .B(_01921_),
    .Y(_05524_));
 sky130_fd_sc_hd__o21ai_0 _25320_ (.A1(_01921_),
    .A2(_05299_),
    .B1(_05524_),
    .Y(_00625_));
 sky130_fd_sc_hd__nand2_1 _25321_ (.A(_02553_),
    .B(_05502_),
    .Y(_05525_));
 sky130_fd_sc_hd__nand2_1 _25322_ (.A(\gen_regfile_ff.register_file_i.rf_reg[232] ),
    .B(_05506_),
    .Y(_05526_));
 sky130_fd_sc_hd__nand2_1 _25323_ (.A(_05525_),
    .B(_05526_),
    .Y(_00626_));
 sky130_fd_sc_hd__nand2_1 _25324_ (.A(_02653_),
    .B(_05502_),
    .Y(_05527_));
 sky130_fd_sc_hd__nand2_1 _25325_ (.A(\gen_regfile_ff.register_file_i.rf_reg[233] ),
    .B(_05506_),
    .Y(_05528_));
 sky130_fd_sc_hd__nand2_1 _25326_ (.A(_05527_),
    .B(_05528_),
    .Y(_00627_));
 sky130_fd_sc_hd__nand2_1 _25327_ (.A(_02761_),
    .B(net255),
    .Y(_05529_));
 sky130_fd_sc_hd__nand2_1 _25328_ (.A(\gen_regfile_ff.register_file_i.rf_reg[234] ),
    .B(_05506_),
    .Y(_05530_));
 sky130_fd_sc_hd__nand2_1 _25329_ (.A(_05529_),
    .B(_05530_),
    .Y(_00628_));
 sky130_fd_sc_hd__nand2_1 _25330_ (.A(_02849_),
    .B(net255),
    .Y(_05531_));
 sky130_fd_sc_hd__nand2_1 _25331_ (.A(\gen_regfile_ff.register_file_i.rf_reg[235] ),
    .B(_05506_),
    .Y(_05532_));
 sky130_fd_sc_hd__nand2_1 _25332_ (.A(_05531_),
    .B(_05532_),
    .Y(_00629_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_200 ();
 sky130_fd_sc_hd__nand2_1 _25334_ (.A(_02974_),
    .B(net255),
    .Y(_05534_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_199 ();
 sky130_fd_sc_hd__nand2_1 _25336_ (.A(\gen_regfile_ff.register_file_i.rf_reg[236] ),
    .B(_05506_),
    .Y(_05536_));
 sky130_fd_sc_hd__nand2_1 _25337_ (.A(_05534_),
    .B(_05536_),
    .Y(_00630_));
 sky130_fd_sc_hd__nand2_1 _25338_ (.A(_03080_),
    .B(_05502_),
    .Y(_05537_));
 sky130_fd_sc_hd__nand2_1 _25339_ (.A(\gen_regfile_ff.register_file_i.rf_reg[237] ),
    .B(_05506_),
    .Y(_05538_));
 sky130_fd_sc_hd__nand2_1 _25340_ (.A(_05537_),
    .B(_05538_),
    .Y(_00631_));
 sky130_fd_sc_hd__nand2_1 _25341_ (.A(_03214_),
    .B(net255),
    .Y(_05539_));
 sky130_fd_sc_hd__nand2_1 _25342_ (.A(\gen_regfile_ff.register_file_i.rf_reg[238] ),
    .B(_05506_),
    .Y(_05540_));
 sky130_fd_sc_hd__nand2_1 _25343_ (.A(_05539_),
    .B(_05540_),
    .Y(_00632_));
 sky130_fd_sc_hd__nand2_1 _25344_ (.A(_03348_),
    .B(_05502_),
    .Y(_05541_));
 sky130_fd_sc_hd__nand2_1 _25345_ (.A(\gen_regfile_ff.register_file_i.rf_reg[239] ),
    .B(_05506_),
    .Y(_05542_));
 sky130_fd_sc_hd__nand2_1 _25346_ (.A(_05541_),
    .B(_05542_),
    .Y(_00633_));
 sky130_fd_sc_hd__nand2_1 _25347_ (.A(\gen_regfile_ff.register_file_i.rf_reg[240] ),
    .B(_05506_),
    .Y(_05543_));
 sky130_fd_sc_hd__o21ai_0 _25348_ (.A1(_03481_),
    .A2(_05506_),
    .B1(_05543_),
    .Y(_00634_));
 sky130_fd_sc_hd__nand2_1 _25349_ (.A(_03614_),
    .B(_05502_),
    .Y(_05544_));
 sky130_fd_sc_hd__nand2_1 _25350_ (.A(\gen_regfile_ff.register_file_i.rf_reg[241] ),
    .B(_05506_),
    .Y(_05545_));
 sky130_fd_sc_hd__nand2_1 _25351_ (.A(_05544_),
    .B(_05545_),
    .Y(_00635_));
 sky130_fd_sc_hd__nand2_1 _25352_ (.A(_01916_),
    .B(_03982_),
    .Y(_05546_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_198 ();
 sky130_fd_sc_hd__nand2_1 _25354_ (.A(\gen_regfile_ff.register_file_i.rf_reg[52] ),
    .B(_01921_),
    .Y(_05548_));
 sky130_fd_sc_hd__nand2_1 _25355_ (.A(_05546_),
    .B(_05548_),
    .Y(_00636_));
 sky130_fd_sc_hd__nand2_1 _25356_ (.A(_03739_),
    .B(_05502_),
    .Y(_05549_));
 sky130_fd_sc_hd__nand2_1 _25357_ (.A(\gen_regfile_ff.register_file_i.rf_reg[242] ),
    .B(_05506_),
    .Y(_05550_));
 sky130_fd_sc_hd__nand2_1 _25358_ (.A(_05549_),
    .B(_05550_),
    .Y(_00637_));
 sky130_fd_sc_hd__nand2_1 _25359_ (.A(_03866_),
    .B(_05502_),
    .Y(_05551_));
 sky130_fd_sc_hd__nand2_1 _25360_ (.A(\gen_regfile_ff.register_file_i.rf_reg[243] ),
    .B(_05506_),
    .Y(_05552_));
 sky130_fd_sc_hd__nand2_1 _25361_ (.A(_05551_),
    .B(_05552_),
    .Y(_00638_));
 sky130_fd_sc_hd__nand2_1 _25362_ (.A(_03982_),
    .B(net255),
    .Y(_05553_));
 sky130_fd_sc_hd__nand2_1 _25363_ (.A(\gen_regfile_ff.register_file_i.rf_reg[244] ),
    .B(_05506_),
    .Y(_05554_));
 sky130_fd_sc_hd__nand2_1 _25364_ (.A(_05553_),
    .B(_05554_),
    .Y(_00639_));
 sky130_fd_sc_hd__nand2_1 _25365_ (.A(net1584),
    .B(net255),
    .Y(_05555_));
 sky130_fd_sc_hd__nand2_1 _25366_ (.A(\gen_regfile_ff.register_file_i.rf_reg[245] ),
    .B(_05506_),
    .Y(_05556_));
 sky130_fd_sc_hd__nand2_1 _25367_ (.A(_05555_),
    .B(_05556_),
    .Y(_00640_));
 sky130_fd_sc_hd__mux2_4 _25368_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[246] ),
    .A1(_04252_),
    .S(net255),
    .X(_00641_));
 sky130_fd_sc_hd__nand2_1 _25369_ (.A(_04390_),
    .B(net255),
    .Y(_05557_));
 sky130_fd_sc_hd__nand2_1 _25370_ (.A(\gen_regfile_ff.register_file_i.rf_reg[247] ),
    .B(_05506_),
    .Y(_05558_));
 sky130_fd_sc_hd__nand2_1 _25371_ (.A(_05557_),
    .B(_05558_),
    .Y(_00642_));
 sky130_fd_sc_hd__nand2_2 _25372_ (.A(net1270),
    .B(net255),
    .Y(_05559_));
 sky130_fd_sc_hd__nand2_1 _25373_ (.A(\gen_regfile_ff.register_file_i.rf_reg[248] ),
    .B(_05506_),
    .Y(_05560_));
 sky130_fd_sc_hd__nand2_1 _25374_ (.A(_05559_),
    .B(_05560_),
    .Y(_00643_));
 sky130_fd_sc_hd__nand2_1 _25375_ (.A(net1564),
    .B(_05502_),
    .Y(_05561_));
 sky130_fd_sc_hd__nand2_1 _25376_ (.A(\gen_regfile_ff.register_file_i.rf_reg[249] ),
    .B(_05506_),
    .Y(_05562_));
 sky130_fd_sc_hd__nand2_1 _25377_ (.A(_05561_),
    .B(_05562_),
    .Y(_00644_));
 sky130_fd_sc_hd__nand2_2 _25378_ (.A(net1514),
    .B(net255),
    .Y(_05563_));
 sky130_fd_sc_hd__nand2_1 _25379_ (.A(\gen_regfile_ff.register_file_i.rf_reg[250] ),
    .B(_05506_),
    .Y(_05564_));
 sky130_fd_sc_hd__nand2_1 _25380_ (.A(_05563_),
    .B(_05564_),
    .Y(_00645_));
 sky130_fd_sc_hd__nand2_1 _25381_ (.A(net1529),
    .B(net255),
    .Y(_05565_));
 sky130_fd_sc_hd__nand2_1 _25382_ (.A(\gen_regfile_ff.register_file_i.rf_reg[251] ),
    .B(_05506_),
    .Y(_05566_));
 sky130_fd_sc_hd__nand2_1 _25383_ (.A(_05565_),
    .B(_05566_),
    .Y(_00646_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_197 ();
 sky130_fd_sc_hd__nand2_1 _25385_ (.A(_01916_),
    .B(net1584),
    .Y(_05568_));
 sky130_fd_sc_hd__nand2_1 _25386_ (.A(\gen_regfile_ff.register_file_i.rf_reg[53] ),
    .B(_01921_),
    .Y(_05569_));
 sky130_fd_sc_hd__nand2_1 _25387_ (.A(_05568_),
    .B(_05569_),
    .Y(_00647_));
 sky130_fd_sc_hd__mux2_4 _25388_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[252] ),
    .A1(_04975_),
    .S(net255),
    .X(_00648_));
 sky130_fd_sc_hd__nor2_1 _25389_ (.A(_05084_),
    .B(_05506_),
    .Y(_05570_));
 sky130_fd_sc_hd__a22o_1 _25390_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[253] ),
    .A2(_05506_),
    .B1(_05079_),
    .B2(_05570_),
    .X(_00649_));
 sky130_fd_sc_hd__mux2_4 _25391_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[254] ),
    .A1(net1237),
    .S(_05502_),
    .X(_00650_));
 sky130_fd_sc_hd__nor2_1 _25392_ (.A(_05264_),
    .B(_05506_),
    .Y(_05571_));
 sky130_fd_sc_hd__a22o_1 _25393_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[255] ),
    .A2(_05506_),
    .B1(_05261_),
    .B2(_05571_),
    .X(_00651_));
 sky130_fd_sc_hd__nand3b_4 _25394_ (.A_N(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .B(_02115_),
    .C(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .Y(_05572_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_196 ();
 sky130_fd_sc_hd__nor2_8 _25396_ (.A(_08194_),
    .B(_05572_),
    .Y(_05574_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_195 ();
 sky130_fd_sc_hd__nand2_1 _25398_ (.A(_01909_),
    .B(_05574_),
    .Y(_05576_));
 sky130_fd_sc_hd__nor3b_4 _25399_ (.A(_01912_),
    .B(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .C_N(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .Y(_05577_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_194 ();
 sky130_fd_sc_hd__nand2_8 _25401_ (.A(_02121_),
    .B(_05577_),
    .Y(_05579_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_193 ();
 sky130_fd_sc_hd__nand2_1 _25403_ (.A(\gen_regfile_ff.register_file_i.rf_reg[256] ),
    .B(_05579_),
    .Y(_05581_));
 sky130_fd_sc_hd__nand2_1 _25404_ (.A(_05576_),
    .B(_05581_),
    .Y(_00652_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_192 ();
 sky130_fd_sc_hd__nand2_1 _25406_ (.A(\gen_regfile_ff.register_file_i.rf_reg[257] ),
    .B(_05579_),
    .Y(_05583_));
 sky130_fd_sc_hd__o21ai_0 _25407_ (.A1(_05299_),
    .A2(_05579_),
    .B1(_05583_),
    .Y(_00653_));
 sky130_fd_sc_hd__nand2_1 _25408_ (.A(_05326_),
    .B(_05574_),
    .Y(_05584_));
 sky130_fd_sc_hd__nand2_1 _25409_ (.A(\gen_regfile_ff.register_file_i.rf_reg[258] ),
    .B(_05579_),
    .Y(_05585_));
 sky130_fd_sc_hd__nand2_1 _25410_ (.A(_05584_),
    .B(_05585_),
    .Y(_00654_));
 sky130_fd_sc_hd__nand2_1 _25411_ (.A(\gen_regfile_ff.register_file_i.rf_reg[259] ),
    .B(_05579_),
    .Y(_05586_));
 sky130_fd_sc_hd__o21ai_0 _25412_ (.A1(_05351_),
    .A2(_05579_),
    .B1(_05586_),
    .Y(_00655_));
 sky130_fd_sc_hd__nand2_1 _25413_ (.A(_02113_),
    .B(_05574_),
    .Y(_05587_));
 sky130_fd_sc_hd__nand2_1 _25414_ (.A(\gen_regfile_ff.register_file_i.rf_reg[260] ),
    .B(_05579_),
    .Y(_05588_));
 sky130_fd_sc_hd__nand2_1 _25415_ (.A(_05587_),
    .B(_05588_),
    .Y(_00656_));
 sky130_fd_sc_hd__nand2_1 _25416_ (.A(_02250_),
    .B(_05574_),
    .Y(_05589_));
 sky130_fd_sc_hd__nand2_1 _25417_ (.A(\gen_regfile_ff.register_file_i.rf_reg[261] ),
    .B(_05579_),
    .Y(_05590_));
 sky130_fd_sc_hd__nand2_1 _25418_ (.A(_05589_),
    .B(_05590_),
    .Y(_00657_));
 sky130_fd_sc_hd__mux2_4 _25419_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[54] ),
    .A1(_04252_),
    .S(_01916_),
    .X(_00658_));
 sky130_fd_sc_hd__nand2_1 _25420_ (.A(_02360_),
    .B(_05574_),
    .Y(_05591_));
 sky130_fd_sc_hd__nand2_1 _25421_ (.A(\gen_regfile_ff.register_file_i.rf_reg[262] ),
    .B(_05579_),
    .Y(_05592_));
 sky130_fd_sc_hd__nand2_1 _25422_ (.A(_05591_),
    .B(_05592_),
    .Y(_00659_));
 sky130_fd_sc_hd__nand2_1 _25423_ (.A(_02468_),
    .B(_05574_),
    .Y(_05593_));
 sky130_fd_sc_hd__nand2_1 _25424_ (.A(\gen_regfile_ff.register_file_i.rf_reg[263] ),
    .B(_05579_),
    .Y(_05594_));
 sky130_fd_sc_hd__nand2_1 _25425_ (.A(_05593_),
    .B(_05594_),
    .Y(_00660_));
 sky130_fd_sc_hd__nand2_1 _25426_ (.A(_02553_),
    .B(_05574_),
    .Y(_05595_));
 sky130_fd_sc_hd__nand2_1 _25427_ (.A(\gen_regfile_ff.register_file_i.rf_reg[264] ),
    .B(_05579_),
    .Y(_05596_));
 sky130_fd_sc_hd__nand2_1 _25428_ (.A(_05595_),
    .B(_05596_),
    .Y(_00661_));
 sky130_fd_sc_hd__nand2_1 _25429_ (.A(_02653_),
    .B(_05574_),
    .Y(_05597_));
 sky130_fd_sc_hd__nand2_1 _25430_ (.A(\gen_regfile_ff.register_file_i.rf_reg[265] ),
    .B(_05579_),
    .Y(_05598_));
 sky130_fd_sc_hd__nand2_1 _25431_ (.A(_05597_),
    .B(_05598_),
    .Y(_00662_));
 sky130_fd_sc_hd__nand2_1 _25432_ (.A(_02761_),
    .B(_05574_),
    .Y(_05599_));
 sky130_fd_sc_hd__nand2_1 _25433_ (.A(\gen_regfile_ff.register_file_i.rf_reg[266] ),
    .B(_05579_),
    .Y(_05600_));
 sky130_fd_sc_hd__nand2_1 _25434_ (.A(_05599_),
    .B(_05600_),
    .Y(_00663_));
 sky130_fd_sc_hd__nand2_1 _25435_ (.A(_02849_),
    .B(_05574_),
    .Y(_05601_));
 sky130_fd_sc_hd__nand2_1 _25436_ (.A(\gen_regfile_ff.register_file_i.rf_reg[267] ),
    .B(_05579_),
    .Y(_05602_));
 sky130_fd_sc_hd__nand2_1 _25437_ (.A(_05601_),
    .B(_05602_),
    .Y(_00664_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_191 ();
 sky130_fd_sc_hd__nand2_1 _25439_ (.A(_02974_),
    .B(_05574_),
    .Y(_05604_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_190 ();
 sky130_fd_sc_hd__nand2_1 _25441_ (.A(\gen_regfile_ff.register_file_i.rf_reg[268] ),
    .B(_05579_),
    .Y(_05606_));
 sky130_fd_sc_hd__nand2_1 _25442_ (.A(_05604_),
    .B(_05606_),
    .Y(_00665_));
 sky130_fd_sc_hd__nand2_1 _25443_ (.A(_03080_),
    .B(_05574_),
    .Y(_05607_));
 sky130_fd_sc_hd__nand2_1 _25444_ (.A(\gen_regfile_ff.register_file_i.rf_reg[269] ),
    .B(_05579_),
    .Y(_05608_));
 sky130_fd_sc_hd__nand2_1 _25445_ (.A(_05607_),
    .B(_05608_),
    .Y(_00666_));
 sky130_fd_sc_hd__nand2_1 _25446_ (.A(_03214_),
    .B(_05574_),
    .Y(_05609_));
 sky130_fd_sc_hd__nand2_1 _25447_ (.A(\gen_regfile_ff.register_file_i.rf_reg[270] ),
    .B(_05579_),
    .Y(_05610_));
 sky130_fd_sc_hd__nand2_1 _25448_ (.A(_05609_),
    .B(_05610_),
    .Y(_00667_));
 sky130_fd_sc_hd__nand2_1 _25449_ (.A(_03348_),
    .B(_05574_),
    .Y(_05611_));
 sky130_fd_sc_hd__nand2_1 _25450_ (.A(\gen_regfile_ff.register_file_i.rf_reg[271] ),
    .B(_05579_),
    .Y(_05612_));
 sky130_fd_sc_hd__nand2_1 _25451_ (.A(_05611_),
    .B(_05612_),
    .Y(_00668_));
 sky130_fd_sc_hd__nand2_1 _25452_ (.A(_01916_),
    .B(_04390_),
    .Y(_05613_));
 sky130_fd_sc_hd__nand2_1 _25453_ (.A(\gen_regfile_ff.register_file_i.rf_reg[55] ),
    .B(_01921_),
    .Y(_05614_));
 sky130_fd_sc_hd__nand2_1 _25454_ (.A(_05613_),
    .B(_05614_),
    .Y(_00669_));
 sky130_fd_sc_hd__nand2_1 _25455_ (.A(\gen_regfile_ff.register_file_i.rf_reg[272] ),
    .B(_05579_),
    .Y(_05615_));
 sky130_fd_sc_hd__o21ai_0 _25456_ (.A1(_03481_),
    .A2(_05579_),
    .B1(_05615_),
    .Y(_00670_));
 sky130_fd_sc_hd__nand2_1 _25457_ (.A(net1575),
    .B(_05574_),
    .Y(_05616_));
 sky130_fd_sc_hd__nand2_1 _25458_ (.A(\gen_regfile_ff.register_file_i.rf_reg[273] ),
    .B(_05579_),
    .Y(_05617_));
 sky130_fd_sc_hd__nand2_1 _25459_ (.A(_05616_),
    .B(_05617_),
    .Y(_00671_));
 sky130_fd_sc_hd__nand2_1 _25460_ (.A(net1576),
    .B(_05574_),
    .Y(_05618_));
 sky130_fd_sc_hd__nand2_1 _25461_ (.A(\gen_regfile_ff.register_file_i.rf_reg[274] ),
    .B(_05579_),
    .Y(_05619_));
 sky130_fd_sc_hd__nand2_1 _25462_ (.A(_05618_),
    .B(_05619_),
    .Y(_00672_));
 sky130_fd_sc_hd__nand2_1 _25463_ (.A(net1551),
    .B(_05574_),
    .Y(_05620_));
 sky130_fd_sc_hd__nand2_1 _25464_ (.A(\gen_regfile_ff.register_file_i.rf_reg[275] ),
    .B(_05579_),
    .Y(_05621_));
 sky130_fd_sc_hd__nand2_1 _25465_ (.A(_05620_),
    .B(_05621_),
    .Y(_00673_));
 sky130_fd_sc_hd__nand2_1 _25466_ (.A(_03982_),
    .B(_05574_),
    .Y(_05622_));
 sky130_fd_sc_hd__nand2_1 _25467_ (.A(\gen_regfile_ff.register_file_i.rf_reg[276] ),
    .B(_05579_),
    .Y(_05623_));
 sky130_fd_sc_hd__nand2_1 _25468_ (.A(_05622_),
    .B(_05623_),
    .Y(_00674_));
 sky130_fd_sc_hd__nand2_1 _25469_ (.A(net1584),
    .B(_05574_),
    .Y(_05624_));
 sky130_fd_sc_hd__nand2_1 _25470_ (.A(\gen_regfile_ff.register_file_i.rf_reg[277] ),
    .B(_05579_),
    .Y(_05625_));
 sky130_fd_sc_hd__nand2_1 _25471_ (.A(_05624_),
    .B(_05625_),
    .Y(_00675_));
 sky130_fd_sc_hd__mux2_4 _25472_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[278] ),
    .A1(net1326),
    .S(_05574_),
    .X(_00676_));
 sky130_fd_sc_hd__nand2_2 _25473_ (.A(net1523),
    .B(_05574_),
    .Y(_05626_));
 sky130_fd_sc_hd__nand2_1 _25474_ (.A(\gen_regfile_ff.register_file_i.rf_reg[279] ),
    .B(_05579_),
    .Y(_05627_));
 sky130_fd_sc_hd__nand2_1 _25475_ (.A(_05626_),
    .B(_05627_),
    .Y(_00677_));
 sky130_fd_sc_hd__nand2_4 _25476_ (.A(net1270),
    .B(_05574_),
    .Y(_05628_));
 sky130_fd_sc_hd__nand2_1 _25477_ (.A(\gen_regfile_ff.register_file_i.rf_reg[280] ),
    .B(_05579_),
    .Y(_05629_));
 sky130_fd_sc_hd__nand2_2 _25478_ (.A(_05628_),
    .B(_05629_),
    .Y(_00678_));
 sky130_fd_sc_hd__nand2_1 _25479_ (.A(net1586),
    .B(_05574_),
    .Y(_05630_));
 sky130_fd_sc_hd__nand2_1 _25480_ (.A(\gen_regfile_ff.register_file_i.rf_reg[281] ),
    .B(_05579_),
    .Y(_05631_));
 sky130_fd_sc_hd__nand2_1 _25481_ (.A(_05630_),
    .B(_05631_),
    .Y(_00679_));
 sky130_fd_sc_hd__nand2_1 _25482_ (.A(_04535_),
    .B(_01916_),
    .Y(_05632_));
 sky130_fd_sc_hd__nand2_1 _25483_ (.A(\gen_regfile_ff.register_file_i.rf_reg[56] ),
    .B(_01921_),
    .Y(_05633_));
 sky130_fd_sc_hd__nand2_1 _25484_ (.A(_05632_),
    .B(_05633_),
    .Y(_00680_));
 sky130_fd_sc_hd__nand2_2 _25485_ (.A(net1536),
    .B(_05574_),
    .Y(_05634_));
 sky130_fd_sc_hd__nand2_1 _25486_ (.A(\gen_regfile_ff.register_file_i.rf_reg[282] ),
    .B(_05579_),
    .Y(_05635_));
 sky130_fd_sc_hd__nand2_1 _25487_ (.A(_05634_),
    .B(_05635_),
    .Y(_00681_));
 sky130_fd_sc_hd__nand2_2 _25488_ (.A(net1529),
    .B(_05574_),
    .Y(_05636_));
 sky130_fd_sc_hd__nand2_1 _25489_ (.A(\gen_regfile_ff.register_file_i.rf_reg[283] ),
    .B(_05579_),
    .Y(_05637_));
 sky130_fd_sc_hd__nand2_1 _25490_ (.A(_05636_),
    .B(_05637_),
    .Y(_00682_));
 sky130_fd_sc_hd__mux2_4 _25491_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[284] ),
    .A1(net250),
    .S(_05574_),
    .X(_00683_));
 sky130_fd_sc_hd__nor2_1 _25492_ (.A(_05084_),
    .B(_05579_),
    .Y(_05638_));
 sky130_fd_sc_hd__a22o_1 _25493_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[285] ),
    .A2(_05579_),
    .B1(net1254),
    .B2(_05638_),
    .X(_00684_));
 sky130_fd_sc_hd__mux2_4 _25494_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[286] ),
    .A1(net685),
    .S(_05574_),
    .X(_00685_));
 sky130_fd_sc_hd__nor2_1 _25495_ (.A(_05264_),
    .B(_05579_),
    .Y(_05639_));
 sky130_fd_sc_hd__a22o_1 _25496_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[287] ),
    .A2(_05579_),
    .B1(net957),
    .B2(_05639_),
    .X(_00686_));
 sky130_fd_sc_hd__nor3_4 _25497_ (.A(net448),
    .B(_01915_),
    .C(_05572_),
    .Y(_05640_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_189 ();
 sky130_fd_sc_hd__nand2_1 _25499_ (.A(_01909_),
    .B(net263),
    .Y(_05642_));
 sky130_fd_sc_hd__nand2_8 _25500_ (.A(_05271_),
    .B(net1250),
    .Y(_05643_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_188 ();
 sky130_fd_sc_hd__nand2_1 _25502_ (.A(\gen_regfile_ff.register_file_i.rf_reg[288] ),
    .B(_05643_),
    .Y(_05645_));
 sky130_fd_sc_hd__nand2_1 _25503_ (.A(_05642_),
    .B(_05645_),
    .Y(_00687_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_187 ();
 sky130_fd_sc_hd__nand2_1 _25505_ (.A(\gen_regfile_ff.register_file_i.rf_reg[289] ),
    .B(_05643_),
    .Y(_05647_));
 sky130_fd_sc_hd__o21ai_0 _25506_ (.A1(_05299_),
    .A2(_05643_),
    .B1(_05647_),
    .Y(_00688_));
 sky130_fd_sc_hd__nand2_1 _25507_ (.A(_05326_),
    .B(net263),
    .Y(_05648_));
 sky130_fd_sc_hd__nand2_1 _25508_ (.A(\gen_regfile_ff.register_file_i.rf_reg[290] ),
    .B(_05643_),
    .Y(_05649_));
 sky130_fd_sc_hd__nand2_1 _25509_ (.A(_05648_),
    .B(_05649_),
    .Y(_00689_));
 sky130_fd_sc_hd__nand2_1 _25510_ (.A(\gen_regfile_ff.register_file_i.rf_reg[291] ),
    .B(_05643_),
    .Y(_05650_));
 sky130_fd_sc_hd__o21ai_0 _25511_ (.A1(_05351_),
    .A2(_05643_),
    .B1(_05650_),
    .Y(_00690_));
 sky130_fd_sc_hd__nand2_4 _25512_ (.A(net1564),
    .B(_01916_),
    .Y(_05651_));
 sky130_fd_sc_hd__nand2_1 _25513_ (.A(\gen_regfile_ff.register_file_i.rf_reg[57] ),
    .B(_01921_),
    .Y(_05652_));
 sky130_fd_sc_hd__nand2_2 _25514_ (.A(_05651_),
    .B(_05652_),
    .Y(_00691_));
 sky130_fd_sc_hd__nand2_1 _25515_ (.A(_02113_),
    .B(net264),
    .Y(_05653_));
 sky130_fd_sc_hd__nand2_1 _25516_ (.A(\gen_regfile_ff.register_file_i.rf_reg[292] ),
    .B(_05643_),
    .Y(_05654_));
 sky130_fd_sc_hd__nand2_1 _25517_ (.A(_05653_),
    .B(_05654_),
    .Y(_00692_));
 sky130_fd_sc_hd__nand2_1 _25518_ (.A(_02250_),
    .B(net264),
    .Y(_05655_));
 sky130_fd_sc_hd__nand2_1 _25519_ (.A(\gen_regfile_ff.register_file_i.rf_reg[293] ),
    .B(_05643_),
    .Y(_05656_));
 sky130_fd_sc_hd__nand2_1 _25520_ (.A(_05655_),
    .B(_05656_),
    .Y(_00693_));
 sky130_fd_sc_hd__nand2_1 _25521_ (.A(_02360_),
    .B(net264),
    .Y(_05657_));
 sky130_fd_sc_hd__nand2_1 _25522_ (.A(\gen_regfile_ff.register_file_i.rf_reg[294] ),
    .B(_05643_),
    .Y(_05658_));
 sky130_fd_sc_hd__nand2_1 _25523_ (.A(_05657_),
    .B(_05658_),
    .Y(_00694_));
 sky130_fd_sc_hd__nand2_1 _25524_ (.A(_02468_),
    .B(net264),
    .Y(_05659_));
 sky130_fd_sc_hd__nand2_1 _25525_ (.A(\gen_regfile_ff.register_file_i.rf_reg[295] ),
    .B(_05643_),
    .Y(_05660_));
 sky130_fd_sc_hd__nand2_1 _25526_ (.A(_05659_),
    .B(_05660_),
    .Y(_00695_));
 sky130_fd_sc_hd__nand2_1 _25527_ (.A(_02553_),
    .B(net263),
    .Y(_05661_));
 sky130_fd_sc_hd__nand2_1 _25528_ (.A(\gen_regfile_ff.register_file_i.rf_reg[296] ),
    .B(_05643_),
    .Y(_05662_));
 sky130_fd_sc_hd__nand2_1 _25529_ (.A(_05661_),
    .B(_05662_),
    .Y(_00696_));
 sky130_fd_sc_hd__nand2_1 _25530_ (.A(_02653_),
    .B(_05640_),
    .Y(_05663_));
 sky130_fd_sc_hd__nand2_1 _25531_ (.A(\gen_regfile_ff.register_file_i.rf_reg[297] ),
    .B(_05643_),
    .Y(_05664_));
 sky130_fd_sc_hd__nand2_1 _25532_ (.A(_05663_),
    .B(_05664_),
    .Y(_00697_));
 sky130_fd_sc_hd__nand2_1 _25533_ (.A(_02761_),
    .B(net264),
    .Y(_05665_));
 sky130_fd_sc_hd__nand2_1 _25534_ (.A(\gen_regfile_ff.register_file_i.rf_reg[298] ),
    .B(_05643_),
    .Y(_05666_));
 sky130_fd_sc_hd__nand2_1 _25535_ (.A(_05665_),
    .B(_05666_),
    .Y(_00698_));
 sky130_fd_sc_hd__nand2_1 _25536_ (.A(_02849_),
    .B(net263),
    .Y(_05667_));
 sky130_fd_sc_hd__nand2_1 _25537_ (.A(\gen_regfile_ff.register_file_i.rf_reg[299] ),
    .B(_05643_),
    .Y(_05668_));
 sky130_fd_sc_hd__nand2_1 _25538_ (.A(_05667_),
    .B(_05668_),
    .Y(_00699_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_186 ();
 sky130_fd_sc_hd__nand2_1 _25540_ (.A(_02974_),
    .B(_05640_),
    .Y(_05670_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_185 ();
 sky130_fd_sc_hd__nand2_1 _25542_ (.A(\gen_regfile_ff.register_file_i.rf_reg[300] ),
    .B(_05643_),
    .Y(_05672_));
 sky130_fd_sc_hd__nand2_1 _25543_ (.A(_05670_),
    .B(_05672_),
    .Y(_00700_));
 sky130_fd_sc_hd__nand2_1 _25544_ (.A(_03080_),
    .B(net263),
    .Y(_05673_));
 sky130_fd_sc_hd__nand2_1 _25545_ (.A(\gen_regfile_ff.register_file_i.rf_reg[301] ),
    .B(_05643_),
    .Y(_05674_));
 sky130_fd_sc_hd__nand2_1 _25546_ (.A(_05673_),
    .B(_05674_),
    .Y(_00701_));
 sky130_fd_sc_hd__nand2_4 _25547_ (.A(net1515),
    .B(_01916_),
    .Y(_05675_));
 sky130_fd_sc_hd__nand2_1 _25548_ (.A(\gen_regfile_ff.register_file_i.rf_reg[58] ),
    .B(_01921_),
    .Y(_05676_));
 sky130_fd_sc_hd__nand2_2 _25549_ (.A(_05675_),
    .B(_05676_),
    .Y(_00702_));
 sky130_fd_sc_hd__nand2_1 _25550_ (.A(_03214_),
    .B(net264),
    .Y(_05677_));
 sky130_fd_sc_hd__nand2_1 _25551_ (.A(\gen_regfile_ff.register_file_i.rf_reg[302] ),
    .B(_05643_),
    .Y(_05678_));
 sky130_fd_sc_hd__nand2_1 _25552_ (.A(_05677_),
    .B(_05678_),
    .Y(_00703_));
 sky130_fd_sc_hd__nand2_1 _25553_ (.A(_03348_),
    .B(net263),
    .Y(_05679_));
 sky130_fd_sc_hd__nand2_1 _25554_ (.A(\gen_regfile_ff.register_file_i.rf_reg[303] ),
    .B(_05643_),
    .Y(_05680_));
 sky130_fd_sc_hd__nand2_1 _25555_ (.A(_05679_),
    .B(_05680_),
    .Y(_00704_));
 sky130_fd_sc_hd__nand2_1 _25556_ (.A(\gen_regfile_ff.register_file_i.rf_reg[304] ),
    .B(_05643_),
    .Y(_05681_));
 sky130_fd_sc_hd__o21ai_0 _25557_ (.A1(_03481_),
    .A2(_05643_),
    .B1(_05681_),
    .Y(_00705_));
 sky130_fd_sc_hd__nand2_1 _25558_ (.A(_03614_),
    .B(_05640_),
    .Y(_05682_));
 sky130_fd_sc_hd__nand2_1 _25559_ (.A(\gen_regfile_ff.register_file_i.rf_reg[305] ),
    .B(_05643_),
    .Y(_05683_));
 sky130_fd_sc_hd__nand2_1 _25560_ (.A(_05682_),
    .B(_05683_),
    .Y(_00706_));
 sky130_fd_sc_hd__nand2_1 _25561_ (.A(net1576),
    .B(net263),
    .Y(_05684_));
 sky130_fd_sc_hd__nand2_1 _25562_ (.A(\gen_regfile_ff.register_file_i.rf_reg[306] ),
    .B(_05643_),
    .Y(_05685_));
 sky130_fd_sc_hd__nand2_1 _25563_ (.A(_05684_),
    .B(_05685_),
    .Y(_00707_));
 sky130_fd_sc_hd__nand2_1 _25564_ (.A(net1551),
    .B(net263),
    .Y(_05686_));
 sky130_fd_sc_hd__nand2_1 _25565_ (.A(\gen_regfile_ff.register_file_i.rf_reg[307] ),
    .B(_05643_),
    .Y(_05687_));
 sky130_fd_sc_hd__nand2_1 _25566_ (.A(_05686_),
    .B(_05687_),
    .Y(_00708_));
 sky130_fd_sc_hd__nand2_1 _25567_ (.A(net1544),
    .B(net264),
    .Y(_05688_));
 sky130_fd_sc_hd__nand2_1 _25568_ (.A(\gen_regfile_ff.register_file_i.rf_reg[308] ),
    .B(_05643_),
    .Y(_05689_));
 sky130_fd_sc_hd__nand2_1 _25569_ (.A(_05688_),
    .B(_05689_),
    .Y(_00709_));
 sky130_fd_sc_hd__nand2_1 _25570_ (.A(net1584),
    .B(net263),
    .Y(_05690_));
 sky130_fd_sc_hd__nand2_1 _25571_ (.A(\gen_regfile_ff.register_file_i.rf_reg[309] ),
    .B(_05643_),
    .Y(_05691_));
 sky130_fd_sc_hd__nand2_1 _25572_ (.A(_05690_),
    .B(_05691_),
    .Y(_00710_));
 sky130_fd_sc_hd__mux2_4 _25573_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[310] ),
    .A1(net1517),
    .S(net264),
    .X(_00711_));
 sky130_fd_sc_hd__nand2_2 _25574_ (.A(net1523),
    .B(net264),
    .Y(_05692_));
 sky130_fd_sc_hd__nand2_1 _25575_ (.A(\gen_regfile_ff.register_file_i.rf_reg[311] ),
    .B(_05643_),
    .Y(_05693_));
 sky130_fd_sc_hd__nand2_1 _25576_ (.A(_05692_),
    .B(_05693_),
    .Y(_00712_));
 sky130_fd_sc_hd__nand2_2 _25577_ (.A(net1529),
    .B(_01916_),
    .Y(_05694_));
 sky130_fd_sc_hd__nand2_1 _25578_ (.A(\gen_regfile_ff.register_file_i.rf_reg[59] ),
    .B(_01921_),
    .Y(_05695_));
 sky130_fd_sc_hd__nand2_1 _25579_ (.A(_05694_),
    .B(_05695_),
    .Y(_00713_));
 sky130_fd_sc_hd__nand2_2 _25580_ (.A(net1270),
    .B(net264),
    .Y(_05696_));
 sky130_fd_sc_hd__nand2_1 _25581_ (.A(\gen_regfile_ff.register_file_i.rf_reg[312] ),
    .B(_05643_),
    .Y(_05697_));
 sky130_fd_sc_hd__nand2_2 _25582_ (.A(_05696_),
    .B(_05697_),
    .Y(_00714_));
 sky130_fd_sc_hd__nand2_1 _25583_ (.A(net252),
    .B(net263),
    .Y(_05698_));
 sky130_fd_sc_hd__nand2_1 _25584_ (.A(\gen_regfile_ff.register_file_i.rf_reg[313] ),
    .B(_05643_),
    .Y(_05699_));
 sky130_fd_sc_hd__nand2_1 _25585_ (.A(_05698_),
    .B(_05699_),
    .Y(_00715_));
 sky130_fd_sc_hd__nand2_2 _25586_ (.A(net1536),
    .B(net263),
    .Y(_05700_));
 sky130_fd_sc_hd__nand2_1 _25587_ (.A(\gen_regfile_ff.register_file_i.rf_reg[314] ),
    .B(_05643_),
    .Y(_05701_));
 sky130_fd_sc_hd__nand2_1 _25588_ (.A(_05700_),
    .B(_05701_),
    .Y(_00716_));
 sky130_fd_sc_hd__nand2_2 _25589_ (.A(net1542),
    .B(net263),
    .Y(_05702_));
 sky130_fd_sc_hd__nand2_1 _25590_ (.A(\gen_regfile_ff.register_file_i.rf_reg[315] ),
    .B(_05643_),
    .Y(_05703_));
 sky130_fd_sc_hd__nand2_1 _25591_ (.A(_05702_),
    .B(_05703_),
    .Y(_00717_));
 sky130_fd_sc_hd__mux2_4 _25592_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[316] ),
    .A1(net250),
    .S(_05640_),
    .X(_00718_));
 sky130_fd_sc_hd__nor2_1 _25593_ (.A(_05084_),
    .B(_05643_),
    .Y(_05704_));
 sky130_fd_sc_hd__a22o_1 _25594_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[317] ),
    .A2(_05643_),
    .B1(net1249),
    .B2(_05704_),
    .X(_00719_));
 sky130_fd_sc_hd__mux2_4 _25595_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[318] ),
    .A1(net685),
    .S(net263),
    .X(_00720_));
 sky130_fd_sc_hd__nor2_1 _25596_ (.A(_05264_),
    .B(_05643_),
    .Y(_05705_));
 sky130_fd_sc_hd__a22o_1 _25597_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[319] ),
    .A2(_05643_),
    .B1(_05705_),
    .B2(net652),
    .X(_00721_));
 sky130_fd_sc_hd__nor3_4 _25598_ (.A(net446),
    .B(_05432_),
    .C(_05572_),
    .Y(_05706_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_184 ();
 sky130_fd_sc_hd__nand2_1 _25600_ (.A(_01909_),
    .B(net261),
    .Y(_05708_));
 sky130_fd_sc_hd__nand2_8 _25601_ (.A(_05436_),
    .B(net1251),
    .Y(_05709_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_183 ();
 sky130_fd_sc_hd__nand2_1 _25603_ (.A(\gen_regfile_ff.register_file_i.rf_reg[320] ),
    .B(_05709_),
    .Y(_05711_));
 sky130_fd_sc_hd__nand2_1 _25604_ (.A(_05708_),
    .B(_05711_),
    .Y(_00722_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_182 ();
 sky130_fd_sc_hd__nand2_1 _25606_ (.A(\gen_regfile_ff.register_file_i.rf_reg[321] ),
    .B(_05709_),
    .Y(_05713_));
 sky130_fd_sc_hd__o21ai_0 _25607_ (.A1(_05299_),
    .A2(_05709_),
    .B1(_05713_),
    .Y(_00723_));
 sky130_fd_sc_hd__mux2_4 _25608_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[60] ),
    .A1(net885),
    .S(_01916_),
    .X(_00724_));
 sky130_fd_sc_hd__nand2_1 _25609_ (.A(_05326_),
    .B(net261),
    .Y(_05714_));
 sky130_fd_sc_hd__nand2_1 _25610_ (.A(\gen_regfile_ff.register_file_i.rf_reg[322] ),
    .B(_05709_),
    .Y(_05715_));
 sky130_fd_sc_hd__nand2_1 _25611_ (.A(_05714_),
    .B(_05715_),
    .Y(_00725_));
 sky130_fd_sc_hd__nand2_1 _25612_ (.A(\gen_regfile_ff.register_file_i.rf_reg[323] ),
    .B(_05709_),
    .Y(_05716_));
 sky130_fd_sc_hd__o21ai_0 _25613_ (.A1(_05351_),
    .A2(_05709_),
    .B1(_05716_),
    .Y(_00726_));
 sky130_fd_sc_hd__nand2_1 _25614_ (.A(_02113_),
    .B(net262),
    .Y(_05717_));
 sky130_fd_sc_hd__nand2_1 _25615_ (.A(\gen_regfile_ff.register_file_i.rf_reg[324] ),
    .B(_05709_),
    .Y(_05718_));
 sky130_fd_sc_hd__nand2_1 _25616_ (.A(_05717_),
    .B(_05718_),
    .Y(_00727_));
 sky130_fd_sc_hd__nand2_1 _25617_ (.A(_02250_),
    .B(net262),
    .Y(_05719_));
 sky130_fd_sc_hd__nand2_1 _25618_ (.A(\gen_regfile_ff.register_file_i.rf_reg[325] ),
    .B(_05709_),
    .Y(_05720_));
 sky130_fd_sc_hd__nand2_1 _25619_ (.A(_05719_),
    .B(_05720_),
    .Y(_00728_));
 sky130_fd_sc_hd__nand2_1 _25620_ (.A(_02360_),
    .B(net262),
    .Y(_05721_));
 sky130_fd_sc_hd__nand2_1 _25621_ (.A(\gen_regfile_ff.register_file_i.rf_reg[326] ),
    .B(_05709_),
    .Y(_05722_));
 sky130_fd_sc_hd__nand2_1 _25622_ (.A(_05721_),
    .B(_05722_),
    .Y(_00729_));
 sky130_fd_sc_hd__nand2_1 _25623_ (.A(_02468_),
    .B(net262),
    .Y(_05723_));
 sky130_fd_sc_hd__nand2_1 _25624_ (.A(\gen_regfile_ff.register_file_i.rf_reg[327] ),
    .B(_05709_),
    .Y(_05724_));
 sky130_fd_sc_hd__nand2_1 _25625_ (.A(_05723_),
    .B(_05724_),
    .Y(_00730_));
 sky130_fd_sc_hd__nand2_1 _25626_ (.A(_02553_),
    .B(net261),
    .Y(_05725_));
 sky130_fd_sc_hd__nand2_1 _25627_ (.A(\gen_regfile_ff.register_file_i.rf_reg[328] ),
    .B(_05709_),
    .Y(_05726_));
 sky130_fd_sc_hd__nand2_1 _25628_ (.A(_05725_),
    .B(_05726_),
    .Y(_00731_));
 sky130_fd_sc_hd__nand2_1 _25629_ (.A(_02653_),
    .B(_05706_),
    .Y(_05727_));
 sky130_fd_sc_hd__nand2_1 _25630_ (.A(\gen_regfile_ff.register_file_i.rf_reg[329] ),
    .B(_05709_),
    .Y(_05728_));
 sky130_fd_sc_hd__nand2_1 _25631_ (.A(_05727_),
    .B(_05728_),
    .Y(_00732_));
 sky130_fd_sc_hd__nand2_1 _25632_ (.A(_02761_),
    .B(net262),
    .Y(_05729_));
 sky130_fd_sc_hd__nand2_1 _25633_ (.A(\gen_regfile_ff.register_file_i.rf_reg[330] ),
    .B(_05709_),
    .Y(_05730_));
 sky130_fd_sc_hd__nand2_1 _25634_ (.A(_05729_),
    .B(_05730_),
    .Y(_00733_));
 sky130_fd_sc_hd__nand2_1 _25635_ (.A(_02849_),
    .B(net262),
    .Y(_05731_));
 sky130_fd_sc_hd__nand2_1 _25636_ (.A(\gen_regfile_ff.register_file_i.rf_reg[331] ),
    .B(_05709_),
    .Y(_05732_));
 sky130_fd_sc_hd__nand2_1 _25637_ (.A(_05731_),
    .B(_05732_),
    .Y(_00734_));
 sky130_fd_sc_hd__nor2_1 _25638_ (.A(_01921_),
    .B(_05084_),
    .Y(_05733_));
 sky130_fd_sc_hd__a22o_1 _25639_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[61] ),
    .A2(_01921_),
    .B1(_05079_),
    .B2(_05733_),
    .X(_00735_));
 sky130_fd_sc_hd__nand2_1 _25640_ (.A(_01916_),
    .B(_05326_),
    .Y(_05734_));
 sky130_fd_sc_hd__nand2_1 _25641_ (.A(\gen_regfile_ff.register_file_i.rf_reg[34] ),
    .B(_01921_),
    .Y(_05735_));
 sky130_fd_sc_hd__nand2_1 _25642_ (.A(_05734_),
    .B(_05735_),
    .Y(_00736_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_181 ();
 sky130_fd_sc_hd__nand2_1 _25644_ (.A(_02974_),
    .B(_05706_),
    .Y(_05737_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_180 ();
 sky130_fd_sc_hd__nand2_1 _25646_ (.A(\gen_regfile_ff.register_file_i.rf_reg[332] ),
    .B(_05709_),
    .Y(_05739_));
 sky130_fd_sc_hd__nand2_1 _25647_ (.A(_05737_),
    .B(_05739_),
    .Y(_00737_));
 sky130_fd_sc_hd__nand2_1 _25648_ (.A(_03080_),
    .B(net261),
    .Y(_05740_));
 sky130_fd_sc_hd__nand2_1 _25649_ (.A(\gen_regfile_ff.register_file_i.rf_reg[333] ),
    .B(_05709_),
    .Y(_05741_));
 sky130_fd_sc_hd__nand2_1 _25650_ (.A(_05740_),
    .B(_05741_),
    .Y(_00738_));
 sky130_fd_sc_hd__nand2_1 _25651_ (.A(_03214_),
    .B(net262),
    .Y(_05742_));
 sky130_fd_sc_hd__nand2_1 _25652_ (.A(\gen_regfile_ff.register_file_i.rf_reg[334] ),
    .B(_05709_),
    .Y(_05743_));
 sky130_fd_sc_hd__nand2_1 _25653_ (.A(_05742_),
    .B(_05743_),
    .Y(_00739_));
 sky130_fd_sc_hd__nand2_1 _25654_ (.A(_03348_),
    .B(net261),
    .Y(_05744_));
 sky130_fd_sc_hd__nand2_1 _25655_ (.A(\gen_regfile_ff.register_file_i.rf_reg[335] ),
    .B(_05709_),
    .Y(_05745_));
 sky130_fd_sc_hd__nand2_1 _25656_ (.A(_05744_),
    .B(_05745_),
    .Y(_00740_));
 sky130_fd_sc_hd__nand2_1 _25657_ (.A(\gen_regfile_ff.register_file_i.rf_reg[336] ),
    .B(_05709_),
    .Y(_05746_));
 sky130_fd_sc_hd__o21ai_0 _25658_ (.A1(_03481_),
    .A2(_05709_),
    .B1(_05746_),
    .Y(_00741_));
 sky130_fd_sc_hd__nand2_1 _25659_ (.A(_03614_),
    .B(_05706_),
    .Y(_05747_));
 sky130_fd_sc_hd__nand2_1 _25660_ (.A(\gen_regfile_ff.register_file_i.rf_reg[337] ),
    .B(_05709_),
    .Y(_05748_));
 sky130_fd_sc_hd__nand2_1 _25661_ (.A(_05747_),
    .B(_05748_),
    .Y(_00742_));
 sky130_fd_sc_hd__nand2_1 _25662_ (.A(net1576),
    .B(net261),
    .Y(_05749_));
 sky130_fd_sc_hd__nand2_1 _25663_ (.A(\gen_regfile_ff.register_file_i.rf_reg[338] ),
    .B(_05709_),
    .Y(_05750_));
 sky130_fd_sc_hd__nand2_1 _25664_ (.A(_05749_),
    .B(_05750_),
    .Y(_00743_));
 sky130_fd_sc_hd__nand2_1 _25665_ (.A(net1551),
    .B(net261),
    .Y(_05751_));
 sky130_fd_sc_hd__nand2_1 _25666_ (.A(\gen_regfile_ff.register_file_i.rf_reg[339] ),
    .B(_05709_),
    .Y(_05752_));
 sky130_fd_sc_hd__nand2_1 _25667_ (.A(_05751_),
    .B(_05752_),
    .Y(_00744_));
 sky130_fd_sc_hd__nand2_1 _25668_ (.A(_03982_),
    .B(net262),
    .Y(_05753_));
 sky130_fd_sc_hd__nand2_1 _25669_ (.A(\gen_regfile_ff.register_file_i.rf_reg[340] ),
    .B(_05709_),
    .Y(_05754_));
 sky130_fd_sc_hd__nand2_1 _25670_ (.A(_05753_),
    .B(_05754_),
    .Y(_00745_));
 sky130_fd_sc_hd__nand2_1 _25671_ (.A(net1584),
    .B(net261),
    .Y(_05755_));
 sky130_fd_sc_hd__nand2_1 _25672_ (.A(\gen_regfile_ff.register_file_i.rf_reg[341] ),
    .B(_05709_),
    .Y(_05756_));
 sky130_fd_sc_hd__nand2_1 _25673_ (.A(_05755_),
    .B(_05756_),
    .Y(_00746_));
 sky130_fd_sc_hd__mux2_4 _25674_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[62] ),
    .A1(net1237),
    .S(_01916_),
    .X(_00747_));
 sky130_fd_sc_hd__mux2_4 _25675_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[342] ),
    .A1(net1326),
    .S(net262),
    .X(_00748_));
 sky130_fd_sc_hd__nand2_2 _25676_ (.A(net1523),
    .B(net262),
    .Y(_05757_));
 sky130_fd_sc_hd__nand2_1 _25677_ (.A(\gen_regfile_ff.register_file_i.rf_reg[343] ),
    .B(_05709_),
    .Y(_05758_));
 sky130_fd_sc_hd__nand2_1 _25678_ (.A(_05757_),
    .B(_05758_),
    .Y(_00749_));
 sky130_fd_sc_hd__nand2_4 _25679_ (.A(net1315),
    .B(net262),
    .Y(_05759_));
 sky130_fd_sc_hd__nand2_1 _25680_ (.A(\gen_regfile_ff.register_file_i.rf_reg[344] ),
    .B(_05709_),
    .Y(_05760_));
 sky130_fd_sc_hd__nand2_2 _25681_ (.A(_05759_),
    .B(_05760_),
    .Y(_00750_));
 sky130_fd_sc_hd__nand2_1 _25682_ (.A(net1586),
    .B(net261),
    .Y(_05761_));
 sky130_fd_sc_hd__nand2_1 _25683_ (.A(\gen_regfile_ff.register_file_i.rf_reg[345] ),
    .B(_05709_),
    .Y(_05762_));
 sky130_fd_sc_hd__nand2_1 _25684_ (.A(_05761_),
    .B(_05762_),
    .Y(_00751_));
 sky130_fd_sc_hd__nand2_2 _25685_ (.A(net1536),
    .B(net261),
    .Y(_05763_));
 sky130_fd_sc_hd__nand2_1 _25686_ (.A(\gen_regfile_ff.register_file_i.rf_reg[346] ),
    .B(_05709_),
    .Y(_05764_));
 sky130_fd_sc_hd__nand2_1 _25687_ (.A(_05763_),
    .B(_05764_),
    .Y(_00752_));
 sky130_fd_sc_hd__nand2_2 _25688_ (.A(net261),
    .B(net1529),
    .Y(_05765_));
 sky130_fd_sc_hd__nand2_1 _25689_ (.A(\gen_regfile_ff.register_file_i.rf_reg[347] ),
    .B(_05709_),
    .Y(_05766_));
 sky130_fd_sc_hd__nand2_1 _25690_ (.A(_05765_),
    .B(_05766_),
    .Y(_00753_));
 sky130_fd_sc_hd__mux2_4 _25691_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[348] ),
    .A1(net250),
    .S(_05706_),
    .X(_00754_));
 sky130_fd_sc_hd__nor2_1 _25692_ (.A(_05084_),
    .B(_05709_),
    .Y(_05767_));
 sky130_fd_sc_hd__a22o_1 _25693_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[349] ),
    .A2(_05709_),
    .B1(net1249),
    .B2(_05767_),
    .X(_00755_));
 sky130_fd_sc_hd__mux2_4 _25694_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[350] ),
    .A1(net859),
    .S(net261),
    .X(_00756_));
 sky130_fd_sc_hd__nor2_1 _25695_ (.A(_05264_),
    .B(_05709_),
    .Y(_05768_));
 sky130_fd_sc_hd__a22o_1 _25696_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[351] ),
    .A2(_05709_),
    .B1(net957),
    .B2(_05768_),
    .X(_00757_));
 sky130_fd_sc_hd__nor2_1 _25697_ (.A(_01921_),
    .B(_05264_),
    .Y(_05769_));
 sky130_fd_sc_hd__a22o_1 _25698_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[63] ),
    .A2(_01921_),
    .B1(_05769_),
    .B2(net740),
    .X(_00758_));
 sky130_fd_sc_hd__nor3_4 _25699_ (.A(net447),
    .B(_05501_),
    .C(_05572_),
    .Y(_05770_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_179 ();
 sky130_fd_sc_hd__nand2_1 _25701_ (.A(_01909_),
    .B(net259),
    .Y(_05772_));
 sky130_fd_sc_hd__nand2_8 _25702_ (.A(_05505_),
    .B(net1252),
    .Y(_05773_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_178 ();
 sky130_fd_sc_hd__nand2_1 _25704_ (.A(\gen_regfile_ff.register_file_i.rf_reg[352] ),
    .B(_05773_),
    .Y(_05775_));
 sky130_fd_sc_hd__nand2_1 _25705_ (.A(_05772_),
    .B(_05775_),
    .Y(_00759_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_177 ();
 sky130_fd_sc_hd__nand2_1 _25707_ (.A(\gen_regfile_ff.register_file_i.rf_reg[353] ),
    .B(_05773_),
    .Y(_05777_));
 sky130_fd_sc_hd__o21ai_0 _25708_ (.A1(_05299_),
    .A2(_05773_),
    .B1(_05777_),
    .Y(_00760_));
 sky130_fd_sc_hd__nand2_1 _25709_ (.A(_05326_),
    .B(net259),
    .Y(_05778_));
 sky130_fd_sc_hd__nand2_1 _25710_ (.A(\gen_regfile_ff.register_file_i.rf_reg[354] ),
    .B(_05773_),
    .Y(_05779_));
 sky130_fd_sc_hd__nand2_1 _25711_ (.A(_05778_),
    .B(_05779_),
    .Y(_00761_));
 sky130_fd_sc_hd__nand2_1 _25712_ (.A(\gen_regfile_ff.register_file_i.rf_reg[355] ),
    .B(_05773_),
    .Y(_05780_));
 sky130_fd_sc_hd__o21ai_0 _25713_ (.A1(_05351_),
    .A2(_05773_),
    .B1(_05780_),
    .Y(_00762_));
 sky130_fd_sc_hd__nand2_1 _25714_ (.A(_02113_),
    .B(net260),
    .Y(_05781_));
 sky130_fd_sc_hd__nand2_1 _25715_ (.A(\gen_regfile_ff.register_file_i.rf_reg[356] ),
    .B(_05773_),
    .Y(_05782_));
 sky130_fd_sc_hd__nand2_1 _25716_ (.A(_05781_),
    .B(_05782_),
    .Y(_00763_));
 sky130_fd_sc_hd__nand2_1 _25717_ (.A(_02250_),
    .B(_05770_),
    .Y(_05783_));
 sky130_fd_sc_hd__nand2_1 _25718_ (.A(\gen_regfile_ff.register_file_i.rf_reg[357] ),
    .B(_05773_),
    .Y(_05784_));
 sky130_fd_sc_hd__nand2_1 _25719_ (.A(_05783_),
    .B(_05784_),
    .Y(_00764_));
 sky130_fd_sc_hd__nand2_1 _25720_ (.A(_02360_),
    .B(net260),
    .Y(_05785_));
 sky130_fd_sc_hd__nand2_1 _25721_ (.A(\gen_regfile_ff.register_file_i.rf_reg[358] ),
    .B(_05773_),
    .Y(_05786_));
 sky130_fd_sc_hd__nand2_1 _25722_ (.A(_05785_),
    .B(_05786_),
    .Y(_00765_));
 sky130_fd_sc_hd__nand2_1 _25723_ (.A(_02468_),
    .B(_05770_),
    .Y(_05787_));
 sky130_fd_sc_hd__nand2_1 _25724_ (.A(\gen_regfile_ff.register_file_i.rf_reg[359] ),
    .B(_05773_),
    .Y(_05788_));
 sky130_fd_sc_hd__nand2_1 _25725_ (.A(_05787_),
    .B(_05788_),
    .Y(_00766_));
 sky130_fd_sc_hd__nand2_1 _25726_ (.A(_02553_),
    .B(net259),
    .Y(_05789_));
 sky130_fd_sc_hd__nand2_1 _25727_ (.A(\gen_regfile_ff.register_file_i.rf_reg[360] ),
    .B(_05773_),
    .Y(_05790_));
 sky130_fd_sc_hd__nand2_1 _25728_ (.A(_05789_),
    .B(_05790_),
    .Y(_00767_));
 sky130_fd_sc_hd__nand2_1 _25729_ (.A(_02653_),
    .B(net260),
    .Y(_05791_));
 sky130_fd_sc_hd__nand2_1 _25730_ (.A(\gen_regfile_ff.register_file_i.rf_reg[361] ),
    .B(_05773_),
    .Y(_05792_));
 sky130_fd_sc_hd__nand2_1 _25731_ (.A(_05791_),
    .B(_05792_),
    .Y(_00768_));
 sky130_fd_sc_hd__nor2_8 _25732_ (.A(_01913_),
    .B(_05432_),
    .Y(_05793_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_176 ();
 sky130_fd_sc_hd__nand2_1 _25734_ (.A(_01909_),
    .B(_05793_),
    .Y(_05795_));
 sky130_fd_sc_hd__nor2b_4 _25735_ (.A(net331),
    .B_N(net1021),
    .Y(_05796_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_175 ();
 sky130_fd_sc_hd__nand2_8 _25737_ (.A(_01918_),
    .B(_05796_),
    .Y(_05798_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_174 ();
 sky130_fd_sc_hd__nand2_1 _25739_ (.A(\gen_regfile_ff.register_file_i.rf_reg[64] ),
    .B(_05798_),
    .Y(_05800_));
 sky130_fd_sc_hd__nand2_1 _25740_ (.A(_05795_),
    .B(_05800_),
    .Y(_00769_));
 sky130_fd_sc_hd__nand2_1 _25741_ (.A(_02761_),
    .B(net260),
    .Y(_05801_));
 sky130_fd_sc_hd__nand2_1 _25742_ (.A(\gen_regfile_ff.register_file_i.rf_reg[362] ),
    .B(_05773_),
    .Y(_05802_));
 sky130_fd_sc_hd__nand2_1 _25743_ (.A(_05801_),
    .B(_05802_),
    .Y(_00770_));
 sky130_fd_sc_hd__nand2_1 _25744_ (.A(_02849_),
    .B(net259),
    .Y(_05803_));
 sky130_fd_sc_hd__nand2_1 _25745_ (.A(\gen_regfile_ff.register_file_i.rf_reg[363] ),
    .B(_05773_),
    .Y(_05804_));
 sky130_fd_sc_hd__nand2_1 _25746_ (.A(_05803_),
    .B(_05804_),
    .Y(_00771_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_173 ();
 sky130_fd_sc_hd__nand2_1 _25748_ (.A(_02974_),
    .B(net260),
    .Y(_05806_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_172 ();
 sky130_fd_sc_hd__nand2_1 _25750_ (.A(\gen_regfile_ff.register_file_i.rf_reg[364] ),
    .B(_05773_),
    .Y(_05808_));
 sky130_fd_sc_hd__nand2_1 _25751_ (.A(_05806_),
    .B(_05808_),
    .Y(_00772_));
 sky130_fd_sc_hd__nand2_1 _25752_ (.A(_03080_),
    .B(net259),
    .Y(_05809_));
 sky130_fd_sc_hd__nand2_1 _25753_ (.A(\gen_regfile_ff.register_file_i.rf_reg[365] ),
    .B(_05773_),
    .Y(_05810_));
 sky130_fd_sc_hd__nand2_1 _25754_ (.A(_05809_),
    .B(_05810_),
    .Y(_00773_));
 sky130_fd_sc_hd__nand2_1 _25755_ (.A(_03214_),
    .B(_05770_),
    .Y(_05811_));
 sky130_fd_sc_hd__nand2_1 _25756_ (.A(\gen_regfile_ff.register_file_i.rf_reg[366] ),
    .B(_05773_),
    .Y(_05812_));
 sky130_fd_sc_hd__nand2_1 _25757_ (.A(_05811_),
    .B(_05812_),
    .Y(_00774_));
 sky130_fd_sc_hd__nand2_1 _25758_ (.A(_03348_),
    .B(net259),
    .Y(_05813_));
 sky130_fd_sc_hd__nand2_1 _25759_ (.A(\gen_regfile_ff.register_file_i.rf_reg[367] ),
    .B(_05773_),
    .Y(_05814_));
 sky130_fd_sc_hd__nand2_1 _25760_ (.A(_05813_),
    .B(_05814_),
    .Y(_00775_));
 sky130_fd_sc_hd__nand2_1 _25761_ (.A(\gen_regfile_ff.register_file_i.rf_reg[368] ),
    .B(_05773_),
    .Y(_05815_));
 sky130_fd_sc_hd__o21ai_0 _25762_ (.A1(_03481_),
    .A2(_05773_),
    .B1(_05815_),
    .Y(_00776_));
 sky130_fd_sc_hd__nand2_1 _25763_ (.A(_03614_),
    .B(net260),
    .Y(_05816_));
 sky130_fd_sc_hd__nand2_1 _25764_ (.A(\gen_regfile_ff.register_file_i.rf_reg[369] ),
    .B(_05773_),
    .Y(_05817_));
 sky130_fd_sc_hd__nand2_1 _25765_ (.A(_05816_),
    .B(_05817_),
    .Y(_00777_));
 sky130_fd_sc_hd__nand2_1 _25766_ (.A(net1576),
    .B(net259),
    .Y(_05818_));
 sky130_fd_sc_hd__nand2_1 _25767_ (.A(\gen_regfile_ff.register_file_i.rf_reg[370] ),
    .B(_05773_),
    .Y(_05819_));
 sky130_fd_sc_hd__nand2_1 _25768_ (.A(_05818_),
    .B(_05819_),
    .Y(_00778_));
 sky130_fd_sc_hd__nand2_1 _25769_ (.A(net1551),
    .B(net259),
    .Y(_05820_));
 sky130_fd_sc_hd__nand2_1 _25770_ (.A(\gen_regfile_ff.register_file_i.rf_reg[371] ),
    .B(_05773_),
    .Y(_05821_));
 sky130_fd_sc_hd__nand2_1 _25771_ (.A(_05820_),
    .B(_05821_),
    .Y(_00779_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_171 ();
 sky130_fd_sc_hd__nand2_1 _25773_ (.A(\gen_regfile_ff.register_file_i.rf_reg[65] ),
    .B(_05798_),
    .Y(_05823_));
 sky130_fd_sc_hd__o21ai_0 _25774_ (.A1(_05299_),
    .A2(_05798_),
    .B1(_05823_),
    .Y(_00780_));
 sky130_fd_sc_hd__nand2_1 _25775_ (.A(net1544),
    .B(_05770_),
    .Y(_05824_));
 sky130_fd_sc_hd__nand2_1 _25776_ (.A(\gen_regfile_ff.register_file_i.rf_reg[372] ),
    .B(_05773_),
    .Y(_05825_));
 sky130_fd_sc_hd__nand2_1 _25777_ (.A(_05824_),
    .B(_05825_),
    .Y(_00781_));
 sky130_fd_sc_hd__nand2_1 _25778_ (.A(net1584),
    .B(net259),
    .Y(_05826_));
 sky130_fd_sc_hd__nand2_1 _25779_ (.A(\gen_regfile_ff.register_file_i.rf_reg[373] ),
    .B(_05773_),
    .Y(_05827_));
 sky130_fd_sc_hd__nand2_1 _25780_ (.A(_05826_),
    .B(_05827_),
    .Y(_00782_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_170 ();
 sky130_fd_sc_hd__mux2_4 _25782_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[374] ),
    .A1(_04252_),
    .S(_05770_),
    .X(_00783_));
 sky130_fd_sc_hd__nand2_2 _25783_ (.A(net1523),
    .B(net259),
    .Y(_05829_));
 sky130_fd_sc_hd__nand2_1 _25784_ (.A(\gen_regfile_ff.register_file_i.rf_reg[375] ),
    .B(_05773_),
    .Y(_05830_));
 sky130_fd_sc_hd__nand2_1 _25785_ (.A(_05829_),
    .B(_05830_),
    .Y(_00784_));
 sky130_fd_sc_hd__nand2_2 _25786_ (.A(net1315),
    .B(_05770_),
    .Y(_05831_));
 sky130_fd_sc_hd__nand2_1 _25787_ (.A(\gen_regfile_ff.register_file_i.rf_reg[376] ),
    .B(_05773_),
    .Y(_05832_));
 sky130_fd_sc_hd__nand2_2 _25788_ (.A(_05832_),
    .B(_05831_),
    .Y(_00785_));
 sky130_fd_sc_hd__nand2_1 _25789_ (.A(net1586),
    .B(net259),
    .Y(_05833_));
 sky130_fd_sc_hd__nand2_1 _25790_ (.A(\gen_regfile_ff.register_file_i.rf_reg[377] ),
    .B(_05773_),
    .Y(_05834_));
 sky130_fd_sc_hd__nand2_1 _25791_ (.A(_05833_),
    .B(_05834_),
    .Y(_00786_));
 sky130_fd_sc_hd__nand2_2 _25792_ (.A(net1536),
    .B(net259),
    .Y(_05835_));
 sky130_fd_sc_hd__nand2_1 _25793_ (.A(\gen_regfile_ff.register_file_i.rf_reg[378] ),
    .B(_05773_),
    .Y(_05836_));
 sky130_fd_sc_hd__nand2_1 _25794_ (.A(_05835_),
    .B(_05836_),
    .Y(_00787_));
 sky130_fd_sc_hd__nand2_2 _25795_ (.A(net1542),
    .B(net260),
    .Y(_05837_));
 sky130_fd_sc_hd__nand2_1 _25796_ (.A(\gen_regfile_ff.register_file_i.rf_reg[379] ),
    .B(_05773_),
    .Y(_05838_));
 sky130_fd_sc_hd__nand2_1 _25797_ (.A(_05837_),
    .B(_05838_),
    .Y(_00788_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_169 ();
 sky130_fd_sc_hd__mux2_4 _25799_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[380] ),
    .A1(net250),
    .S(_05770_),
    .X(_00789_));
 sky130_fd_sc_hd__nor2_1 _25800_ (.A(_05084_),
    .B(_05773_),
    .Y(_05840_));
 sky130_fd_sc_hd__a22o_1 _25801_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[381] ),
    .A2(_05773_),
    .B1(net1254),
    .B2(_05840_),
    .X(_00790_));
 sky130_fd_sc_hd__nand2_1 _25802_ (.A(_05326_),
    .B(_05793_),
    .Y(_05841_));
 sky130_fd_sc_hd__nand2_1 _25803_ (.A(\gen_regfile_ff.register_file_i.rf_reg[66] ),
    .B(_05798_),
    .Y(_05842_));
 sky130_fd_sc_hd__nand2_1 _25804_ (.A(_05841_),
    .B(_05842_),
    .Y(_00791_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_168 ();
 sky130_fd_sc_hd__mux2_4 _25806_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[382] ),
    .A1(net859),
    .S(net259),
    .X(_00792_));
 sky130_fd_sc_hd__nor2_1 _25807_ (.A(_05264_),
    .B(_05773_),
    .Y(_05844_));
 sky130_fd_sc_hd__a22o_1 _25808_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[383] ),
    .A2(_05773_),
    .B1(_05844_),
    .B2(net500),
    .X(_00793_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_166 ();
 sky130_fd_sc_hd__and3_4 _25811_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .B(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .C(_02115_),
    .X(_05847_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_165 ();
 sky130_fd_sc_hd__nand2_8 _25813_ (.A(_02121_),
    .B(_05847_),
    .Y(_05849_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_163 ();
 sky130_fd_sc_hd__nand2_1 _25816_ (.A(\gen_regfile_ff.register_file_i.rf_reg[384] ),
    .B(_05849_),
    .Y(_05852_));
 sky130_fd_sc_hd__o31ai_1 _25817_ (.A1(_01732_),
    .A2(net258),
    .A3(_05849_),
    .B1(_05852_),
    .Y(_00794_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_162 ();
 sky130_fd_sc_hd__nand2_1 _25819_ (.A(\gen_regfile_ff.register_file_i.rf_reg[385] ),
    .B(_05849_),
    .Y(_05854_));
 sky130_fd_sc_hd__o21ai_0 _25820_ (.A1(_05299_),
    .A2(_05849_),
    .B1(_05854_),
    .Y(_00795_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_161 ();
 sky130_fd_sc_hd__mux2_1 _25822_ (.A0(_05326_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[386] ),
    .S(_05849_),
    .X(_00796_));
 sky130_fd_sc_hd__nand2_1 _25823_ (.A(\gen_regfile_ff.register_file_i.rf_reg[387] ),
    .B(_05849_),
    .Y(_05856_));
 sky130_fd_sc_hd__o21ai_0 _25824_ (.A1(_05351_),
    .A2(_05849_),
    .B1(_05856_),
    .Y(_00797_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_160 ();
 sky130_fd_sc_hd__mux2_1 _25826_ (.A0(_02113_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[388] ),
    .S(_05849_),
    .X(_00798_));
 sky130_fd_sc_hd__mux2_1 _25827_ (.A0(_02250_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[389] ),
    .S(_05849_),
    .X(_00799_));
 sky130_fd_sc_hd__mux2_1 _25828_ (.A0(_02360_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[390] ),
    .S(_05849_),
    .X(_00800_));
 sky130_fd_sc_hd__mux2_1 _25829_ (.A0(_02468_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[391] ),
    .S(_05849_),
    .X(_00801_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_159 ();
 sky130_fd_sc_hd__nand2_1 _25831_ (.A(\gen_regfile_ff.register_file_i.rf_reg[67] ),
    .B(_05798_),
    .Y(_05859_));
 sky130_fd_sc_hd__o21ai_0 _25832_ (.A1(_05351_),
    .A2(_05798_),
    .B1(_05859_),
    .Y(_00802_));
 sky130_fd_sc_hd__mux2_1 _25833_ (.A0(_02553_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[392] ),
    .S(_05849_),
    .X(_00803_));
 sky130_fd_sc_hd__mux2_1 _25834_ (.A0(_02653_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[393] ),
    .S(_05849_),
    .X(_00804_));
 sky130_fd_sc_hd__mux2_1 _25835_ (.A0(_02761_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[394] ),
    .S(_05849_),
    .X(_00805_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_158 ();
 sky130_fd_sc_hd__mux2_1 _25837_ (.A0(_02849_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[395] ),
    .S(_05849_),
    .X(_00806_));
 sky130_fd_sc_hd__mux2_1 _25838_ (.A0(_02974_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[396] ),
    .S(_05849_),
    .X(_00807_));
 sky130_fd_sc_hd__mux2_1 _25839_ (.A0(_03080_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[397] ),
    .S(_05849_),
    .X(_00808_));
 sky130_fd_sc_hd__mux2_1 _25840_ (.A0(_03214_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[398] ),
    .S(_05849_),
    .X(_00809_));
 sky130_fd_sc_hd__mux2_1 _25841_ (.A0(_03348_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[399] ),
    .S(_05849_),
    .X(_00810_));
 sky130_fd_sc_hd__nand2_1 _25842_ (.A(\gen_regfile_ff.register_file_i.rf_reg[400] ),
    .B(_05849_),
    .Y(_05861_));
 sky130_fd_sc_hd__o21ai_0 _25843_ (.A1(_03481_),
    .A2(_05849_),
    .B1(_05861_),
    .Y(_00811_));
 sky130_fd_sc_hd__mux2_1 _25844_ (.A0(_03614_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[401] ),
    .S(_05849_),
    .X(_00812_));
 sky130_fd_sc_hd__nand2_1 _25845_ (.A(_02113_),
    .B(_05793_),
    .Y(_05862_));
 sky130_fd_sc_hd__nand2_1 _25846_ (.A(\gen_regfile_ff.register_file_i.rf_reg[68] ),
    .B(_05798_),
    .Y(_05863_));
 sky130_fd_sc_hd__nand2_1 _25847_ (.A(_05862_),
    .B(_05863_),
    .Y(_00813_));
 sky130_fd_sc_hd__mux2_1 _25848_ (.A0(net1576),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[402] ),
    .S(_05849_),
    .X(_00814_));
 sky130_fd_sc_hd__mux2_1 _25849_ (.A0(net1551),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[403] ),
    .S(_05849_),
    .X(_00815_));
 sky130_fd_sc_hd__mux2_1 _25850_ (.A0(_03982_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[404] ),
    .S(_05849_),
    .X(_00816_));
 sky130_fd_sc_hd__mux2_1 _25851_ (.A0(net1017),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[405] ),
    .S(_05849_),
    .X(_00817_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_157 ();
 sky130_fd_sc_hd__mux2_4 _25853_ (.A0(net1326),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[406] ),
    .S(_05849_),
    .X(_00818_));
 sky130_fd_sc_hd__mux2_4 _25854_ (.A0(net1504),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[407] ),
    .S(_05849_),
    .X(_00819_));
 sky130_fd_sc_hd__mux2_4 _25855_ (.A0(net1315),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[408] ),
    .S(_05849_),
    .X(_00820_));
 sky130_fd_sc_hd__mux2_1 _25856_ (.A0(net252),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[409] ),
    .S(_05849_),
    .X(_00821_));
 sky130_fd_sc_hd__mux2_4 _25857_ (.A0(net1515),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[410] ),
    .S(_05849_),
    .X(_00822_));
 sky130_fd_sc_hd__mux2_4 _25858_ (.A0(_04865_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[411] ),
    .S(_05849_),
    .X(_00823_));
 sky130_fd_sc_hd__nand2_1 _25859_ (.A(_02250_),
    .B(_05793_),
    .Y(_05865_));
 sky130_fd_sc_hd__nand2_1 _25860_ (.A(\gen_regfile_ff.register_file_i.rf_reg[69] ),
    .B(_05798_),
    .Y(_05866_));
 sky130_fd_sc_hd__nand2_1 _25861_ (.A(_05865_),
    .B(_05866_),
    .Y(_00824_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_156 ();
 sky130_fd_sc_hd__mux2_4 _25863_ (.A0(net885),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[412] ),
    .S(_05849_),
    .X(_00825_));
 sky130_fd_sc_hd__nor2_1 _25864_ (.A(_05084_),
    .B(_05849_),
    .Y(_05868_));
 sky130_fd_sc_hd__a22o_1 _25865_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[413] ),
    .A2(_05849_),
    .B1(net1249),
    .B2(_05868_),
    .X(_00826_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_155 ();
 sky130_fd_sc_hd__mux2_4 _25867_ (.A0(net685),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[414] ),
    .S(_05849_),
    .X(_00827_));
 sky130_fd_sc_hd__nor2_1 _25868_ (.A(_05264_),
    .B(_05849_),
    .Y(_05870_));
 sky130_fd_sc_hd__a22o_1 _25869_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[415] ),
    .A2(_05849_),
    .B1(_05870_),
    .B2(net652),
    .X(_00828_));
 sky130_fd_sc_hd__nand2_8 _25870_ (.A(_05271_),
    .B(_05847_),
    .Y(_05871_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_153 ();
 sky130_fd_sc_hd__nand2_1 _25873_ (.A(\gen_regfile_ff.register_file_i.rf_reg[416] ),
    .B(_05871_),
    .Y(_05874_));
 sky130_fd_sc_hd__o31ai_1 _25874_ (.A1(_01732_),
    .A2(net258),
    .A3(_05871_),
    .B1(_05874_),
    .Y(_00829_));
 sky130_fd_sc_hd__nand2_1 _25875_ (.A(\gen_regfile_ff.register_file_i.rf_reg[417] ),
    .B(_05871_),
    .Y(_05875_));
 sky130_fd_sc_hd__o21ai_0 _25876_ (.A1(_05299_),
    .A2(_05871_),
    .B1(_05875_),
    .Y(_00830_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_151 ();
 sky130_fd_sc_hd__mux2_1 _25879_ (.A0(_05326_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[418] ),
    .S(_05871_),
    .X(_00831_));
 sky130_fd_sc_hd__nand2_1 _25880_ (.A(\gen_regfile_ff.register_file_i.rf_reg[419] ),
    .B(_05871_),
    .Y(_05878_));
 sky130_fd_sc_hd__o21ai_0 _25881_ (.A1(_05351_),
    .A2(_05871_),
    .B1(_05878_),
    .Y(_00832_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_150 ();
 sky130_fd_sc_hd__mux2_1 _25883_ (.A0(_02113_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[420] ),
    .S(_05871_),
    .X(_00833_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_149 ();
 sky130_fd_sc_hd__mux2_1 _25885_ (.A0(_02250_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[421] ),
    .S(_05871_),
    .X(_00834_));
 sky130_fd_sc_hd__nand2_1 _25886_ (.A(_02360_),
    .B(_05793_),
    .Y(_05881_));
 sky130_fd_sc_hd__nand2_1 _25887_ (.A(\gen_regfile_ff.register_file_i.rf_reg[70] ),
    .B(_05798_),
    .Y(_05882_));
 sky130_fd_sc_hd__nand2_1 _25888_ (.A(_05881_),
    .B(_05882_),
    .Y(_00835_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_148 ();
 sky130_fd_sc_hd__mux2_1 _25890_ (.A0(_02360_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[422] ),
    .S(_05871_),
    .X(_00836_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_147 ();
 sky130_fd_sc_hd__mux2_1 _25892_ (.A0(_02468_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[423] ),
    .S(_05871_),
    .X(_00837_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_146 ();
 sky130_fd_sc_hd__mux2_1 _25894_ (.A0(_02553_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[424] ),
    .S(_05871_),
    .X(_00838_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_145 ();
 sky130_fd_sc_hd__mux2_1 _25896_ (.A0(_02653_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[425] ),
    .S(_05871_),
    .X(_00839_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_144 ();
 sky130_fd_sc_hd__mux2_1 _25898_ (.A0(_02761_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[426] ),
    .S(_05871_),
    .X(_00840_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_142 ();
 sky130_fd_sc_hd__mux2_1 _25901_ (.A0(_02849_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[427] ),
    .S(_05871_),
    .X(_00841_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_141 ();
 sky130_fd_sc_hd__mux2_1 _25903_ (.A0(_02974_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[428] ),
    .S(_05871_),
    .X(_00842_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_140 ();
 sky130_fd_sc_hd__mux2_1 _25905_ (.A0(_03080_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[429] ),
    .S(_05871_),
    .X(_00843_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_139 ();
 sky130_fd_sc_hd__mux2_1 _25907_ (.A0(_03214_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[430] ),
    .S(_05871_),
    .X(_00844_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_138 ();
 sky130_fd_sc_hd__mux2_1 _25909_ (.A0(_03348_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[431] ),
    .S(_05871_),
    .X(_00845_));
 sky130_fd_sc_hd__nand2_1 _25910_ (.A(_02468_),
    .B(_05793_),
    .Y(_05894_));
 sky130_fd_sc_hd__nand2_1 _25911_ (.A(\gen_regfile_ff.register_file_i.rf_reg[71] ),
    .B(_05798_),
    .Y(_05895_));
 sky130_fd_sc_hd__nand2_1 _25912_ (.A(_05894_),
    .B(_05895_),
    .Y(_00846_));
 sky130_fd_sc_hd__nand2_1 _25913_ (.A(\gen_regfile_ff.register_file_i.rf_reg[35] ),
    .B(_01921_),
    .Y(_05896_));
 sky130_fd_sc_hd__o21ai_0 _25914_ (.A1(_01921_),
    .A2(_05351_),
    .B1(_05896_),
    .Y(_00847_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_137 ();
 sky130_fd_sc_hd__nand2_1 _25916_ (.A(\gen_regfile_ff.register_file_i.rf_reg[432] ),
    .B(_05871_),
    .Y(_05898_));
 sky130_fd_sc_hd__o21ai_0 _25917_ (.A1(_03481_),
    .A2(_05871_),
    .B1(_05898_),
    .Y(_00848_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_136 ();
 sky130_fd_sc_hd__mux2_1 _25919_ (.A0(_03614_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[433] ),
    .S(_05871_),
    .X(_00849_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_135 ();
 sky130_fd_sc_hd__mux2_1 _25921_ (.A0(net1576),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[434] ),
    .S(_05871_),
    .X(_00850_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_134 ();
 sky130_fd_sc_hd__mux2_1 _25923_ (.A0(_03866_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[435] ),
    .S(_05871_),
    .X(_00851_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_133 ();
 sky130_fd_sc_hd__mux2_1 _25925_ (.A0(_03982_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[436] ),
    .S(_05871_),
    .X(_00852_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_132 ();
 sky130_fd_sc_hd__mux2_1 _25927_ (.A0(net1017),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[437] ),
    .S(_05871_),
    .X(_00853_));
 sky130_fd_sc_hd__mux2_4 _25928_ (.A0(net1327),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[438] ),
    .S(_05871_),
    .X(_00854_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_131 ();
 sky130_fd_sc_hd__mux2_1 _25930_ (.A0(net1475),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[439] ),
    .S(_05871_),
    .X(_00855_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_130 ();
 sky130_fd_sc_hd__mux2_4 _25932_ (.A0(net1315),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[440] ),
    .S(_05871_),
    .X(_00856_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_129 ();
 sky130_fd_sc_hd__mux2_1 _25934_ (.A0(net252),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[441] ),
    .S(_05871_),
    .X(_00857_));
 sky130_fd_sc_hd__nand2_1 _25935_ (.A(_02553_),
    .B(_05793_),
    .Y(_05907_));
 sky130_fd_sc_hd__nand2_1 _25936_ (.A(\gen_regfile_ff.register_file_i.rf_reg[72] ),
    .B(_05798_),
    .Y(_05908_));
 sky130_fd_sc_hd__nand2_1 _25937_ (.A(_05907_),
    .B(_05908_),
    .Y(_00858_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_128 ();
 sky130_fd_sc_hd__mux2_4 _25939_ (.A0(net251),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[442] ),
    .S(_05871_),
    .X(_00859_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_127 ();
 sky130_fd_sc_hd__mux2_1 _25941_ (.A0(net1533),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[443] ),
    .S(_05871_),
    .X(_00860_));
 sky130_fd_sc_hd__mux2_4 _25942_ (.A0(net250),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[444] ),
    .S(_05871_),
    .X(_00861_));
 sky130_fd_sc_hd__nor2_1 _25943_ (.A(_05084_),
    .B(_05871_),
    .Y(_05911_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_126 ();
 sky130_fd_sc_hd__a22o_1 _25945_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[445] ),
    .A2(_05871_),
    .B1(net1249),
    .B2(_05911_),
    .X(_00862_));
 sky130_fd_sc_hd__mux2_4 _25946_ (.A0(net859),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[446] ),
    .S(_05871_),
    .X(_00863_));
 sky130_fd_sc_hd__nor2_1 _25947_ (.A(_05264_),
    .B(_05871_),
    .Y(_05913_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_125 ();
 sky130_fd_sc_hd__a22o_1 _25949_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[447] ),
    .A2(_05871_),
    .B1(_05913_),
    .B2(net500),
    .X(_00864_));
 sky130_fd_sc_hd__nand2_8 _25950_ (.A(_05436_),
    .B(_05847_),
    .Y(_05915_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_123 ();
 sky130_fd_sc_hd__nand2_1 _25953_ (.A(\gen_regfile_ff.register_file_i.rf_reg[448] ),
    .B(_05915_),
    .Y(_05918_));
 sky130_fd_sc_hd__o31ai_1 _25954_ (.A1(_01732_),
    .A2(net258),
    .A3(_05915_),
    .B1(_05918_),
    .Y(_00865_));
 sky130_fd_sc_hd__nand2_1 _25955_ (.A(\gen_regfile_ff.register_file_i.rf_reg[449] ),
    .B(_05915_),
    .Y(_05919_));
 sky130_fd_sc_hd__o21ai_0 _25956_ (.A1(_05299_),
    .A2(_05915_),
    .B1(_05919_),
    .Y(_00866_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_122 ();
 sky130_fd_sc_hd__mux2_1 _25958_ (.A0(_05326_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[450] ),
    .S(_05915_),
    .X(_00867_));
 sky130_fd_sc_hd__nand2_1 _25959_ (.A(\gen_regfile_ff.register_file_i.rf_reg[451] ),
    .B(_05915_),
    .Y(_05921_));
 sky130_fd_sc_hd__o21ai_0 _25960_ (.A1(_05351_),
    .A2(_05915_),
    .B1(_05921_),
    .Y(_00868_));
 sky130_fd_sc_hd__nand2_1 _25961_ (.A(_02653_),
    .B(_05793_),
    .Y(_05922_));
 sky130_fd_sc_hd__nand2_1 _25962_ (.A(\gen_regfile_ff.register_file_i.rf_reg[73] ),
    .B(_05798_),
    .Y(_05923_));
 sky130_fd_sc_hd__nand2_1 _25963_ (.A(_05922_),
    .B(_05923_),
    .Y(_00869_));
 sky130_fd_sc_hd__mux2_1 _25964_ (.A0(_02113_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[452] ),
    .S(_05915_),
    .X(_00870_));
 sky130_fd_sc_hd__mux2_1 _25965_ (.A0(_02250_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[453] ),
    .S(_05915_),
    .X(_00871_));
 sky130_fd_sc_hd__mux2_1 _25966_ (.A0(_02360_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[454] ),
    .S(_05915_),
    .X(_00872_));
 sky130_fd_sc_hd__mux2_1 _25967_ (.A0(_02468_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[455] ),
    .S(_05915_),
    .X(_00873_));
 sky130_fd_sc_hd__mux2_1 _25968_ (.A0(_02553_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[456] ),
    .S(_05915_),
    .X(_00874_));
 sky130_fd_sc_hd__mux2_1 _25969_ (.A0(_02653_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[457] ),
    .S(_05915_),
    .X(_00875_));
 sky130_fd_sc_hd__mux2_1 _25970_ (.A0(_02761_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[458] ),
    .S(_05915_),
    .X(_00876_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_121 ();
 sky130_fd_sc_hd__mux2_1 _25972_ (.A0(_02849_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[459] ),
    .S(_05915_),
    .X(_00877_));
 sky130_fd_sc_hd__mux2_1 _25973_ (.A0(_02974_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[460] ),
    .S(_05915_),
    .X(_00878_));
 sky130_fd_sc_hd__mux2_1 _25974_ (.A0(_03080_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[461] ),
    .S(_05915_),
    .X(_00879_));
 sky130_fd_sc_hd__nand2_1 _25975_ (.A(_02761_),
    .B(_05793_),
    .Y(_05925_));
 sky130_fd_sc_hd__nand2_1 _25976_ (.A(\gen_regfile_ff.register_file_i.rf_reg[74] ),
    .B(_05798_),
    .Y(_05926_));
 sky130_fd_sc_hd__nand2_1 _25977_ (.A(_05925_),
    .B(_05926_),
    .Y(_00880_));
 sky130_fd_sc_hd__mux2_1 _25978_ (.A0(_03214_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[462] ),
    .S(_05915_),
    .X(_00881_));
 sky130_fd_sc_hd__mux2_1 _25979_ (.A0(_03348_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[463] ),
    .S(_05915_),
    .X(_00882_));
 sky130_fd_sc_hd__nand2_1 _25980_ (.A(\gen_regfile_ff.register_file_i.rf_reg[464] ),
    .B(_05915_),
    .Y(_05927_));
 sky130_fd_sc_hd__o21ai_0 _25981_ (.A1(_03481_),
    .A2(_05915_),
    .B1(_05927_),
    .Y(_00883_));
 sky130_fd_sc_hd__mux2_1 _25982_ (.A0(_03614_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[465] ),
    .S(_05915_),
    .X(_00884_));
 sky130_fd_sc_hd__mux2_1 _25983_ (.A0(net1576),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[466] ),
    .S(_05915_),
    .X(_00885_));
 sky130_fd_sc_hd__mux2_1 _25984_ (.A0(net1551),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[467] ),
    .S(_05915_),
    .X(_00886_));
 sky130_fd_sc_hd__mux2_1 _25985_ (.A0(_03982_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[468] ),
    .S(_05915_),
    .X(_00887_));
 sky130_fd_sc_hd__mux2_1 _25986_ (.A0(net1017),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[469] ),
    .S(_05915_),
    .X(_00888_));
 sky130_fd_sc_hd__mux2_4 _25987_ (.A0(net1327),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[470] ),
    .S(_05915_),
    .X(_00889_));
 sky130_fd_sc_hd__mux2_4 _25988_ (.A0(net1475),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[471] ),
    .S(_05915_),
    .X(_00890_));
 sky130_fd_sc_hd__nand2_1 _25989_ (.A(_02849_),
    .B(_05793_),
    .Y(_05928_));
 sky130_fd_sc_hd__nand2_1 _25990_ (.A(\gen_regfile_ff.register_file_i.rf_reg[75] ),
    .B(_05798_),
    .Y(_05929_));
 sky130_fd_sc_hd__nand2_1 _25991_ (.A(_05928_),
    .B(_05929_),
    .Y(_00891_));
 sky130_fd_sc_hd__mux2_4 _25992_ (.A0(net1317),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[472] ),
    .S(_05915_),
    .X(_00892_));
 sky130_fd_sc_hd__mux2_1 _25993_ (.A0(net252),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[473] ),
    .S(_05915_),
    .X(_00893_));
 sky130_fd_sc_hd__mux2_4 _25994_ (.A0(net1515),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[474] ),
    .S(_05915_),
    .X(_00894_));
 sky130_fd_sc_hd__mux2_1 _25995_ (.A0(_04865_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[475] ),
    .S(_05915_),
    .X(_00895_));
 sky130_fd_sc_hd__mux2_4 _25996_ (.A0(net885),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[476] ),
    .S(_05915_),
    .X(_00896_));
 sky130_fd_sc_hd__nor2_1 _25997_ (.A(_05084_),
    .B(_05915_),
    .Y(_05930_));
 sky130_fd_sc_hd__a22o_1 _25998_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[477] ),
    .A2(_05915_),
    .B1(net1246),
    .B2(_05930_),
    .X(_00897_));
 sky130_fd_sc_hd__mux2_4 _25999_ (.A0(net685),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[478] ),
    .S(_05915_),
    .X(_00898_));
 sky130_fd_sc_hd__nor2_1 _26000_ (.A(_05264_),
    .B(_05915_),
    .Y(_05931_));
 sky130_fd_sc_hd__a22o_1 _26001_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[479] ),
    .A2(_05915_),
    .B1(_05931_),
    .B2(net652),
    .X(_00899_));
 sky130_fd_sc_hd__nand2_8 _26002_ (.A(_05505_),
    .B(_05847_),
    .Y(_05932_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_119 ();
 sky130_fd_sc_hd__nand2_1 _26005_ (.A(\gen_regfile_ff.register_file_i.rf_reg[480] ),
    .B(_05932_),
    .Y(_05935_));
 sky130_fd_sc_hd__o31ai_1 _26006_ (.A1(_01732_),
    .A2(net258),
    .A3(_05932_),
    .B1(_05935_),
    .Y(_00900_));
 sky130_fd_sc_hd__nand2_1 _26007_ (.A(\gen_regfile_ff.register_file_i.rf_reg[481] ),
    .B(_05932_),
    .Y(_05936_));
 sky130_fd_sc_hd__o21ai_0 _26008_ (.A1(_05299_),
    .A2(_05932_),
    .B1(_05936_),
    .Y(_00901_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_118 ();
 sky130_fd_sc_hd__nand2_1 _26010_ (.A(_02974_),
    .B(_05793_),
    .Y(_05938_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_117 ();
 sky130_fd_sc_hd__nand2_1 _26012_ (.A(\gen_regfile_ff.register_file_i.rf_reg[76] ),
    .B(_05798_),
    .Y(_05940_));
 sky130_fd_sc_hd__nand2_1 _26013_ (.A(_05938_),
    .B(_05940_),
    .Y(_00902_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_116 ();
 sky130_fd_sc_hd__mux2_1 _26015_ (.A0(_05326_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[482] ),
    .S(_05932_),
    .X(_00903_));
 sky130_fd_sc_hd__nand2_1 _26016_ (.A(\gen_regfile_ff.register_file_i.rf_reg[483] ),
    .B(_05932_),
    .Y(_05942_));
 sky130_fd_sc_hd__o21ai_0 _26017_ (.A1(_05351_),
    .A2(_05932_),
    .B1(_05942_),
    .Y(_00904_));
 sky130_fd_sc_hd__mux2_1 _26018_ (.A0(_02113_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[484] ),
    .S(_05932_),
    .X(_00905_));
 sky130_fd_sc_hd__mux2_1 _26019_ (.A0(_02250_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[485] ),
    .S(_05932_),
    .X(_00906_));
 sky130_fd_sc_hd__mux2_1 _26020_ (.A0(_02360_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[486] ),
    .S(_05932_),
    .X(_00907_));
 sky130_fd_sc_hd__mux2_1 _26021_ (.A0(_02468_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[487] ),
    .S(_05932_),
    .X(_00908_));
 sky130_fd_sc_hd__mux2_1 _26022_ (.A0(_02553_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[488] ),
    .S(_05932_),
    .X(_00909_));
 sky130_fd_sc_hd__mux2_1 _26023_ (.A0(_02653_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[489] ),
    .S(_05932_),
    .X(_00910_));
 sky130_fd_sc_hd__mux2_1 _26024_ (.A0(_02761_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[490] ),
    .S(_05932_),
    .X(_00911_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_115 ();
 sky130_fd_sc_hd__mux2_1 _26026_ (.A0(_02849_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[491] ),
    .S(_05932_),
    .X(_00912_));
 sky130_fd_sc_hd__nand2_1 _26027_ (.A(_03080_),
    .B(_05793_),
    .Y(_05944_));
 sky130_fd_sc_hd__nand2_1 _26028_ (.A(\gen_regfile_ff.register_file_i.rf_reg[77] ),
    .B(_05798_),
    .Y(_05945_));
 sky130_fd_sc_hd__nand2_1 _26029_ (.A(_05944_),
    .B(_05945_),
    .Y(_00913_));
 sky130_fd_sc_hd__mux2_1 _26030_ (.A0(_02974_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[492] ),
    .S(_05932_),
    .X(_00914_));
 sky130_fd_sc_hd__mux2_1 _26031_ (.A0(_03080_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[493] ),
    .S(_05932_),
    .X(_00915_));
 sky130_fd_sc_hd__mux2_1 _26032_ (.A0(_03214_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[494] ),
    .S(_05932_),
    .X(_00916_));
 sky130_fd_sc_hd__mux2_1 _26033_ (.A0(_03348_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[495] ),
    .S(_05932_),
    .X(_00917_));
 sky130_fd_sc_hd__nand2_1 _26034_ (.A(\gen_regfile_ff.register_file_i.rf_reg[496] ),
    .B(_05932_),
    .Y(_05946_));
 sky130_fd_sc_hd__o21ai_0 _26035_ (.A1(_03481_),
    .A2(_05932_),
    .B1(_05946_),
    .Y(_00918_));
 sky130_fd_sc_hd__mux2_1 _26036_ (.A0(_03614_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[497] ),
    .S(_05932_),
    .X(_00919_));
 sky130_fd_sc_hd__mux2_1 _26037_ (.A0(net1576),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[498] ),
    .S(_05932_),
    .X(_00920_));
 sky130_fd_sc_hd__mux2_1 _26038_ (.A0(net1551),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[499] ),
    .S(_05932_),
    .X(_00921_));
 sky130_fd_sc_hd__mux2_1 _26039_ (.A0(_03982_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[500] ),
    .S(_05932_),
    .X(_00922_));
 sky130_fd_sc_hd__mux2_1 _26040_ (.A0(net1017),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[501] ),
    .S(_05932_),
    .X(_00923_));
 sky130_fd_sc_hd__nand2_1 _26041_ (.A(_03214_),
    .B(_05793_),
    .Y(_05947_));
 sky130_fd_sc_hd__nand2_1 _26042_ (.A(\gen_regfile_ff.register_file_i.rf_reg[78] ),
    .B(_05798_),
    .Y(_05948_));
 sky130_fd_sc_hd__nand2_1 _26043_ (.A(_05947_),
    .B(_05948_),
    .Y(_00924_));
 sky130_fd_sc_hd__mux2_4 _26044_ (.A0(net1327),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[502] ),
    .S(_05932_),
    .X(_00925_));
 sky130_fd_sc_hd__mux2_1 _26045_ (.A0(net1290),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[503] ),
    .S(_05932_),
    .X(_00926_));
 sky130_fd_sc_hd__mux2_4 _26046_ (.A0(net1317),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[504] ),
    .S(_05932_),
    .X(_00927_));
 sky130_fd_sc_hd__mux2_1 _26047_ (.A0(net252),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[505] ),
    .S(_05932_),
    .X(_00928_));
 sky130_fd_sc_hd__mux2_4 _26048_ (.A0(net1515),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[506] ),
    .S(_05932_),
    .X(_00929_));
 sky130_fd_sc_hd__mux2_4 _26049_ (.A0(_04865_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[507] ),
    .S(_05932_),
    .X(_00930_));
 sky130_fd_sc_hd__mux2_4 _26050_ (.A0(net885),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[508] ),
    .S(_05932_),
    .X(_00931_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_114 ();
 sky130_fd_sc_hd__nor2_1 _26052_ (.A(_05084_),
    .B(_05932_),
    .Y(_05950_));
 sky130_fd_sc_hd__a22o_1 _26053_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[509] ),
    .A2(_05932_),
    .B1(net1254),
    .B2(_05950_),
    .X(_00932_));
 sky130_fd_sc_hd__mux2_4 _26054_ (.A0(net685),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[510] ),
    .S(_05932_),
    .X(_00933_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_113 ();
 sky130_fd_sc_hd__nor2_1 _26056_ (.A(_05264_),
    .B(_05932_),
    .Y(_05952_));
 sky130_fd_sc_hd__a22o_1 _26057_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[511] ),
    .A2(_05932_),
    .B1(net957),
    .B2(_05952_),
    .X(_00934_));
 sky130_fd_sc_hd__nand2_1 _26058_ (.A(_03348_),
    .B(_05793_),
    .Y(_05953_));
 sky130_fd_sc_hd__nand2_1 _26059_ (.A(\gen_regfile_ff.register_file_i.rf_reg[79] ),
    .B(_05798_),
    .Y(_05954_));
 sky130_fd_sc_hd__nand2_1 _26060_ (.A(_05953_),
    .B(_05954_),
    .Y(_00935_));
 sky130_fd_sc_hd__nor2_8 _26061_ (.A(net1021),
    .B(net331),
    .Y(_05955_));
 sky130_fd_sc_hd__nor4b_4 _26062_ (.A(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .B(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .C(_01912_),
    .D_N(net447),
    .Y(_05956_));
 sky130_fd_sc_hd__nand2_8 _26063_ (.A(_05955_),
    .B(net1323),
    .Y(_05957_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_111 ();
 sky130_fd_sc_hd__nand2_1 _26066_ (.A(\gen_regfile_ff.register_file_i.rf_reg[512] ),
    .B(_05957_),
    .Y(_05960_));
 sky130_fd_sc_hd__o31ai_1 _26067_ (.A1(_01732_),
    .A2(net258),
    .A3(_05957_),
    .B1(_05960_),
    .Y(_00936_));
 sky130_fd_sc_hd__nand2_1 _26068_ (.A(\gen_regfile_ff.register_file_i.rf_reg[513] ),
    .B(_05957_),
    .Y(_05961_));
 sky130_fd_sc_hd__o21ai_0 _26069_ (.A1(_05299_),
    .A2(_05957_),
    .B1(_05961_),
    .Y(_00937_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_110 ();
 sky130_fd_sc_hd__mux2_1 _26071_ (.A0(_05326_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[514] ),
    .S(_05957_),
    .X(_00938_));
 sky130_fd_sc_hd__nand2_1 _26072_ (.A(\gen_regfile_ff.register_file_i.rf_reg[515] ),
    .B(_05957_),
    .Y(_05963_));
 sky130_fd_sc_hd__o21ai_0 _26073_ (.A1(_05351_),
    .A2(_05957_),
    .B1(_05963_),
    .Y(_00939_));
 sky130_fd_sc_hd__mux2_1 _26074_ (.A0(_02113_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[516] ),
    .S(_05957_),
    .X(_00940_));
 sky130_fd_sc_hd__mux2_1 _26075_ (.A0(_02250_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[517] ),
    .S(_05957_),
    .X(_00941_));
 sky130_fd_sc_hd__mux2_1 _26076_ (.A0(_02360_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[518] ),
    .S(_05957_),
    .X(_00942_));
 sky130_fd_sc_hd__mux2_1 _26077_ (.A0(_02468_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[519] ),
    .S(_05957_),
    .X(_00943_));
 sky130_fd_sc_hd__mux2_1 _26078_ (.A0(_02553_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[520] ),
    .S(_05957_),
    .X(_00944_));
 sky130_fd_sc_hd__mux2_1 _26079_ (.A0(_02653_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[521] ),
    .S(_05957_),
    .X(_00945_));
 sky130_fd_sc_hd__nand2_1 _26080_ (.A(\gen_regfile_ff.register_file_i.rf_reg[80] ),
    .B(_05798_),
    .Y(_05964_));
 sky130_fd_sc_hd__o21ai_0 _26081_ (.A1(_03481_),
    .A2(_05798_),
    .B1(_05964_),
    .Y(_00946_));
 sky130_fd_sc_hd__mux2_1 _26082_ (.A0(_02761_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[522] ),
    .S(_05957_),
    .X(_00947_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_109 ();
 sky130_fd_sc_hd__mux2_1 _26084_ (.A0(_02849_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[523] ),
    .S(_05957_),
    .X(_00948_));
 sky130_fd_sc_hd__mux2_1 _26085_ (.A0(_02974_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[524] ),
    .S(_05957_),
    .X(_00949_));
 sky130_fd_sc_hd__mux2_1 _26086_ (.A0(_03080_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[525] ),
    .S(_05957_),
    .X(_00950_));
 sky130_fd_sc_hd__mux2_1 _26087_ (.A0(_03214_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[526] ),
    .S(_05957_),
    .X(_00951_));
 sky130_fd_sc_hd__mux2_1 _26088_ (.A0(_03348_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[527] ),
    .S(_05957_),
    .X(_00952_));
 sky130_fd_sc_hd__nand2_1 _26089_ (.A(\gen_regfile_ff.register_file_i.rf_reg[528] ),
    .B(_05957_),
    .Y(_05966_));
 sky130_fd_sc_hd__o21ai_0 _26090_ (.A1(_03481_),
    .A2(_05957_),
    .B1(_05966_),
    .Y(_00953_));
 sky130_fd_sc_hd__mux2_1 _26091_ (.A0(net1575),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[529] ),
    .S(_05957_),
    .X(_00954_));
 sky130_fd_sc_hd__mux2_1 _26092_ (.A0(_03739_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[530] ),
    .S(_05957_),
    .X(_00955_));
 sky130_fd_sc_hd__mux2_1 _26093_ (.A0(_03866_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[531] ),
    .S(_05957_),
    .X(_00956_));
 sky130_fd_sc_hd__nand2_1 _26094_ (.A(_03614_),
    .B(_05793_),
    .Y(_05967_));
 sky130_fd_sc_hd__nand2_1 _26095_ (.A(\gen_regfile_ff.register_file_i.rf_reg[81] ),
    .B(_05798_),
    .Y(_05968_));
 sky130_fd_sc_hd__nand2_1 _26096_ (.A(_05967_),
    .B(_05968_),
    .Y(_00957_));
 sky130_fd_sc_hd__nand2_1 _26097_ (.A(_01916_),
    .B(_02113_),
    .Y(_05969_));
 sky130_fd_sc_hd__nand2_1 _26098_ (.A(\gen_regfile_ff.register_file_i.rf_reg[36] ),
    .B(_01921_),
    .Y(_05970_));
 sky130_fd_sc_hd__nand2_1 _26099_ (.A(_05969_),
    .B(_05970_),
    .Y(_00958_));
 sky130_fd_sc_hd__mux2_4 _26100_ (.A0(net1537),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[532] ),
    .S(_05957_),
    .X(_00959_));
 sky130_fd_sc_hd__mux2_1 _26101_ (.A0(net1017),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[533] ),
    .S(_05957_),
    .X(_00960_));
 sky130_fd_sc_hd__mux2_4 _26102_ (.A0(net1326),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[534] ),
    .S(_05957_),
    .X(_00961_));
 sky130_fd_sc_hd__mux2_4 _26103_ (.A0(net1504),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[535] ),
    .S(_05957_),
    .X(_00962_));
 sky130_fd_sc_hd__mux2_4 _26104_ (.A0(net1271),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[536] ),
    .S(_05957_),
    .X(_00963_));
 sky130_fd_sc_hd__mux2_1 _26105_ (.A0(net252),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[537] ),
    .S(_05957_),
    .X(_00964_));
 sky130_fd_sc_hd__mux2_1 _26106_ (.A0(net251),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[538] ),
    .S(_05957_),
    .X(_00965_));
 sky130_fd_sc_hd__mux2_1 _26107_ (.A0(net1533),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[539] ),
    .S(_05957_),
    .X(_00966_));
 sky130_fd_sc_hd__mux2_4 _26108_ (.A0(net886),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[540] ),
    .S(_05957_),
    .X(_00967_));
 sky130_fd_sc_hd__nor2_1 _26109_ (.A(_05084_),
    .B(_05957_),
    .Y(_05971_));
 sky130_fd_sc_hd__a22o_1 _26110_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[541] ),
    .A2(_05957_),
    .B1(net1246),
    .B2(_05971_),
    .X(_00968_));
 sky130_fd_sc_hd__nand2_1 _26111_ (.A(_03739_),
    .B(_05793_),
    .Y(_05972_));
 sky130_fd_sc_hd__nand2_1 _26112_ (.A(\gen_regfile_ff.register_file_i.rf_reg[82] ),
    .B(_05798_),
    .Y(_05973_));
 sky130_fd_sc_hd__nand2_1 _26113_ (.A(_05972_),
    .B(_05973_),
    .Y(_00969_));
 sky130_fd_sc_hd__mux2_4 _26114_ (.A0(net1237),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[542] ),
    .S(_05957_),
    .X(_00970_));
 sky130_fd_sc_hd__nor2_1 _26115_ (.A(_05264_),
    .B(_05957_),
    .Y(_05974_));
 sky130_fd_sc_hd__a22o_1 _26116_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[543] ),
    .A2(_05957_),
    .B1(_05974_),
    .B2(net500),
    .X(_00971_));
 sky130_fd_sc_hd__nand2_8 _26117_ (.A(_01919_),
    .B(net1324),
    .Y(_05975_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_107 ();
 sky130_fd_sc_hd__nand2_1 _26120_ (.A(\gen_regfile_ff.register_file_i.rf_reg[544] ),
    .B(_05975_),
    .Y(_05978_));
 sky130_fd_sc_hd__o31ai_1 _26121_ (.A1(_01732_),
    .A2(net258),
    .A3(_05975_),
    .B1(_05978_),
    .Y(_00972_));
 sky130_fd_sc_hd__nand2_1 _26122_ (.A(\gen_regfile_ff.register_file_i.rf_reg[545] ),
    .B(_05975_),
    .Y(_05979_));
 sky130_fd_sc_hd__o21ai_0 _26123_ (.A1(_05299_),
    .A2(_05975_),
    .B1(_05979_),
    .Y(_00973_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_106 ();
 sky130_fd_sc_hd__mux2_1 _26125_ (.A0(_05326_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[546] ),
    .S(_05975_),
    .X(_00974_));
 sky130_fd_sc_hd__nand2_1 _26126_ (.A(\gen_regfile_ff.register_file_i.rf_reg[547] ),
    .B(_05975_),
    .Y(_05981_));
 sky130_fd_sc_hd__o21ai_0 _26127_ (.A1(_05351_),
    .A2(_05975_),
    .B1(_05981_),
    .Y(_00975_));
 sky130_fd_sc_hd__mux2_1 _26128_ (.A0(_02113_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[548] ),
    .S(_05975_),
    .X(_00976_));
 sky130_fd_sc_hd__mux2_1 _26129_ (.A0(_02250_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[549] ),
    .S(_05975_),
    .X(_00977_));
 sky130_fd_sc_hd__mux2_1 _26130_ (.A0(_02360_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[550] ),
    .S(_05975_),
    .X(_00978_));
 sky130_fd_sc_hd__mux2_1 _26131_ (.A0(_02468_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[551] ),
    .S(_05975_),
    .X(_00979_));
 sky130_fd_sc_hd__nand2_1 _26132_ (.A(_03866_),
    .B(_05793_),
    .Y(_05982_));
 sky130_fd_sc_hd__nand2_1 _26133_ (.A(\gen_regfile_ff.register_file_i.rf_reg[83] ),
    .B(_05798_),
    .Y(_05983_));
 sky130_fd_sc_hd__nand2_1 _26134_ (.A(_05982_),
    .B(_05983_),
    .Y(_00980_));
 sky130_fd_sc_hd__mux2_1 _26135_ (.A0(_02553_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[552] ),
    .S(_05975_),
    .X(_00981_));
 sky130_fd_sc_hd__mux2_1 _26136_ (.A0(_02653_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[553] ),
    .S(_05975_),
    .X(_00982_));
 sky130_fd_sc_hd__mux2_1 _26137_ (.A0(_02761_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[554] ),
    .S(_05975_),
    .X(_00983_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_105 ();
 sky130_fd_sc_hd__mux2_1 _26139_ (.A0(_02849_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[555] ),
    .S(_05975_),
    .X(_00984_));
 sky130_fd_sc_hd__mux2_1 _26140_ (.A0(_02974_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[556] ),
    .S(_05975_),
    .X(_00985_));
 sky130_fd_sc_hd__mux2_1 _26141_ (.A0(_03080_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[557] ),
    .S(_05975_),
    .X(_00986_));
 sky130_fd_sc_hd__mux2_1 _26142_ (.A0(_03214_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[558] ),
    .S(_05975_),
    .X(_00987_));
 sky130_fd_sc_hd__mux2_1 _26143_ (.A0(_03348_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[559] ),
    .S(_05975_),
    .X(_00988_));
 sky130_fd_sc_hd__nand2_1 _26144_ (.A(\gen_regfile_ff.register_file_i.rf_reg[560] ),
    .B(_05975_),
    .Y(_05985_));
 sky130_fd_sc_hd__o21ai_0 _26145_ (.A1(_03481_),
    .A2(_05975_),
    .B1(_05985_),
    .Y(_00989_));
 sky130_fd_sc_hd__mux2_1 _26146_ (.A0(net1575),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[561] ),
    .S(_05975_),
    .X(_00990_));
 sky130_fd_sc_hd__nand2_1 _26147_ (.A(_03982_),
    .B(_05793_),
    .Y(_05986_));
 sky130_fd_sc_hd__o21ai_0 _26148_ (.A1(_10020_),
    .A2(_05793_),
    .B1(_05986_),
    .Y(_00991_));
 sky130_fd_sc_hd__mux2_1 _26149_ (.A0(_03739_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[562] ),
    .S(_05975_),
    .X(_00992_));
 sky130_fd_sc_hd__mux2_1 _26150_ (.A0(net1551),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[563] ),
    .S(_05975_),
    .X(_00993_));
 sky130_fd_sc_hd__mux2_4 _26151_ (.A0(net1537),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[564] ),
    .S(_05975_),
    .X(_00994_));
 sky130_fd_sc_hd__mux2_1 _26152_ (.A0(net1017),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[565] ),
    .S(_05975_),
    .X(_00995_));
 sky130_fd_sc_hd__mux2_4 _26153_ (.A0(net1327),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[566] ),
    .S(_05975_),
    .X(_00996_));
 sky130_fd_sc_hd__mux2_1 _26154_ (.A0(net1475),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[567] ),
    .S(_05975_),
    .X(_00997_));
 sky130_fd_sc_hd__mux2_1 _26155_ (.A0(net1271),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[568] ),
    .S(_05975_),
    .X(_00998_));
 sky130_fd_sc_hd__mux2_1 _26156_ (.A0(net252),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[569] ),
    .S(_05975_),
    .X(_00999_));
 sky130_fd_sc_hd__mux2_4 _26157_ (.A0(net251),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[570] ),
    .S(_05975_),
    .X(_01000_));
 sky130_fd_sc_hd__mux2_1 _26158_ (.A0(net1533),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[571] ),
    .S(_05975_),
    .X(_01001_));
 sky130_fd_sc_hd__nand2_1 _26159_ (.A(net1017),
    .B(_05793_),
    .Y(_05987_));
 sky130_fd_sc_hd__nand2_1 _26160_ (.A(\gen_regfile_ff.register_file_i.rf_reg[85] ),
    .B(_05798_),
    .Y(_05988_));
 sky130_fd_sc_hd__nand2_1 _26161_ (.A(_05987_),
    .B(_05988_),
    .Y(_01002_));
 sky130_fd_sc_hd__mux2_4 _26162_ (.A0(net886),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[572] ),
    .S(_05975_),
    .X(_01003_));
 sky130_fd_sc_hd__nor2_1 _26163_ (.A(_05084_),
    .B(_05975_),
    .Y(_05989_));
 sky130_fd_sc_hd__a22o_1 _26164_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[573] ),
    .A2(_05975_),
    .B1(net1254),
    .B2(_05989_),
    .X(_01004_));
 sky130_fd_sc_hd__mux2_4 _26165_ (.A0(net1238),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[574] ),
    .S(_05975_),
    .X(_01005_));
 sky130_fd_sc_hd__nor2_1 _26166_ (.A(_05264_),
    .B(_05975_),
    .Y(_05990_));
 sky130_fd_sc_hd__a22o_1 _26167_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[575] ),
    .A2(_05975_),
    .B1(_05990_),
    .B2(net652),
    .X(_01006_));
 sky130_fd_sc_hd__nand2_8 _26168_ (.A(_05796_),
    .B(net1323),
    .Y(_05991_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_103 ();
 sky130_fd_sc_hd__nand2_1 _26171_ (.A(\gen_regfile_ff.register_file_i.rf_reg[576] ),
    .B(_05991_),
    .Y(_05994_));
 sky130_fd_sc_hd__o31ai_1 _26172_ (.A1(_01732_),
    .A2(net258),
    .A3(_05991_),
    .B1(_05994_),
    .Y(_01007_));
 sky130_fd_sc_hd__nand2_1 _26173_ (.A(\gen_regfile_ff.register_file_i.rf_reg[577] ),
    .B(_05991_),
    .Y(_05995_));
 sky130_fd_sc_hd__o21ai_0 _26174_ (.A1(_05299_),
    .A2(_05991_),
    .B1(_05995_),
    .Y(_01008_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_102 ();
 sky130_fd_sc_hd__mux2_1 _26176_ (.A0(_05326_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[578] ),
    .S(_05991_),
    .X(_01009_));
 sky130_fd_sc_hd__nand2_1 _26177_ (.A(\gen_regfile_ff.register_file_i.rf_reg[579] ),
    .B(_05991_),
    .Y(_05997_));
 sky130_fd_sc_hd__o21ai_0 _26178_ (.A1(_05351_),
    .A2(_05991_),
    .B1(_05997_),
    .Y(_01010_));
 sky130_fd_sc_hd__mux2_1 _26179_ (.A0(_02113_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[580] ),
    .S(_05991_),
    .X(_01011_));
 sky130_fd_sc_hd__mux2_1 _26180_ (.A0(_02250_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[581] ),
    .S(_05991_),
    .X(_01012_));
 sky130_fd_sc_hd__mux2_4 _26181_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[86] ),
    .A1(_04252_),
    .S(_05793_),
    .X(_01013_));
 sky130_fd_sc_hd__mux2_1 _26182_ (.A0(_02360_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[582] ),
    .S(_05991_),
    .X(_01014_));
 sky130_fd_sc_hd__mux2_1 _26183_ (.A0(_02468_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[583] ),
    .S(_05991_),
    .X(_01015_));
 sky130_fd_sc_hd__mux2_1 _26184_ (.A0(_02553_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[584] ),
    .S(_05991_),
    .X(_01016_));
 sky130_fd_sc_hd__mux2_1 _26185_ (.A0(_02653_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[585] ),
    .S(_05991_),
    .X(_01017_));
 sky130_fd_sc_hd__mux2_1 _26186_ (.A0(_02761_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[586] ),
    .S(_05991_),
    .X(_01018_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_101 ();
 sky130_fd_sc_hd__mux2_1 _26188_ (.A0(_02849_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[587] ),
    .S(_05991_),
    .X(_01019_));
 sky130_fd_sc_hd__mux2_1 _26189_ (.A0(_02974_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[588] ),
    .S(_05991_),
    .X(_01020_));
 sky130_fd_sc_hd__mux2_1 _26190_ (.A0(_03080_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[589] ),
    .S(_05991_),
    .X(_01021_));
 sky130_fd_sc_hd__mux2_1 _26191_ (.A0(_03214_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[590] ),
    .S(_05991_),
    .X(_01022_));
 sky130_fd_sc_hd__mux2_1 _26192_ (.A0(_03348_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[591] ),
    .S(_05991_),
    .X(_01023_));
 sky130_fd_sc_hd__nand2_1 _26193_ (.A(_05793_),
    .B(_04390_),
    .Y(_05999_));
 sky130_fd_sc_hd__nand2_1 _26194_ (.A(\gen_regfile_ff.register_file_i.rf_reg[87] ),
    .B(_05798_),
    .Y(_06000_));
 sky130_fd_sc_hd__nand2_1 _26195_ (.A(_05999_),
    .B(_06000_),
    .Y(_01024_));
 sky130_fd_sc_hd__nand2_1 _26196_ (.A(\gen_regfile_ff.register_file_i.rf_reg[592] ),
    .B(_05991_),
    .Y(_06001_));
 sky130_fd_sc_hd__o21ai_0 _26197_ (.A1(_03481_),
    .A2(_05991_),
    .B1(_06001_),
    .Y(_01025_));
 sky130_fd_sc_hd__mux2_1 _26198_ (.A0(_03614_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[593] ),
    .S(_05991_),
    .X(_01026_));
 sky130_fd_sc_hd__mux2_1 _26199_ (.A0(net1576),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[594] ),
    .S(_05991_),
    .X(_01027_));
 sky130_fd_sc_hd__mux2_1 _26200_ (.A0(_03866_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[595] ),
    .S(_05991_),
    .X(_01028_));
 sky130_fd_sc_hd__mux2_4 _26201_ (.A0(net1537),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[596] ),
    .S(_05991_),
    .X(_01029_));
 sky130_fd_sc_hd__mux2_1 _26202_ (.A0(net1017),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[597] ),
    .S(_05991_),
    .X(_01030_));
 sky130_fd_sc_hd__mux2_4 _26203_ (.A0(net1517),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[598] ),
    .S(_05991_),
    .X(_01031_));
 sky130_fd_sc_hd__mux2_4 _26204_ (.A0(net1504),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[599] ),
    .S(_05991_),
    .X(_01032_));
 sky130_fd_sc_hd__mux2_4 _26205_ (.A0(net1316),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[600] ),
    .S(_05991_),
    .X(_01033_));
 sky130_fd_sc_hd__mux2_1 _26206_ (.A0(net252),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[601] ),
    .S(_05991_),
    .X(_01034_));
 sky130_fd_sc_hd__nand2_1 _26207_ (.A(_04535_),
    .B(_05793_),
    .Y(_06002_));
 sky130_fd_sc_hd__nand2_1 _26208_ (.A(\gen_regfile_ff.register_file_i.rf_reg[88] ),
    .B(_05798_),
    .Y(_06003_));
 sky130_fd_sc_hd__nand2_1 _26209_ (.A(_06002_),
    .B(_06003_),
    .Y(_01035_));
 sky130_fd_sc_hd__mux2_4 _26210_ (.A0(net251),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[602] ),
    .S(_05991_),
    .X(_01036_));
 sky130_fd_sc_hd__mux2_4 _26211_ (.A0(_04865_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[603] ),
    .S(_05991_),
    .X(_01037_));
 sky130_fd_sc_hd__mux2_4 _26212_ (.A0(net886),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[604] ),
    .S(_05991_),
    .X(_01038_));
 sky130_fd_sc_hd__nor2_1 _26213_ (.A(_05084_),
    .B(_05991_),
    .Y(_06004_));
 sky130_fd_sc_hd__a22o_1 _26214_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[605] ),
    .A2(_05991_),
    .B1(net1246),
    .B2(_06004_),
    .X(_01039_));
 sky130_fd_sc_hd__mux2_4 _26215_ (.A0(net1238),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[606] ),
    .S(_05991_),
    .X(_01040_));
 sky130_fd_sc_hd__nor2_1 _26216_ (.A(_05264_),
    .B(_05991_),
    .Y(_06005_));
 sky130_fd_sc_hd__a22o_1 _26217_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[607] ),
    .A2(_05991_),
    .B1(net957),
    .B2(_06005_),
    .X(_01041_));
 sky130_fd_sc_hd__nand3_4 _26218_ (.A(net1020),
    .B(net331),
    .C(net1324),
    .Y(_06006_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_99 ();
 sky130_fd_sc_hd__nand2_1 _26221_ (.A(\gen_regfile_ff.register_file_i.rf_reg[608] ),
    .B(net1300),
    .Y(_06009_));
 sky130_fd_sc_hd__o31ai_1 _26222_ (.A1(_01732_),
    .A2(net258),
    .A3(net1300),
    .B1(_06009_),
    .Y(_01042_));
 sky130_fd_sc_hd__nand2_1 _26223_ (.A(\gen_regfile_ff.register_file_i.rf_reg[609] ),
    .B(net1300),
    .Y(_06010_));
 sky130_fd_sc_hd__o21ai_0 _26224_ (.A1(_05299_),
    .A2(net1300),
    .B1(_06010_),
    .Y(_01043_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_98 ();
 sky130_fd_sc_hd__mux2_1 _26226_ (.A0(_05326_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[610] ),
    .S(_06006_),
    .X(_01044_));
 sky130_fd_sc_hd__nand2_1 _26227_ (.A(\gen_regfile_ff.register_file_i.rf_reg[611] ),
    .B(net1300),
    .Y(_06012_));
 sky130_fd_sc_hd__o21ai_0 _26228_ (.A1(_05351_),
    .A2(net1300),
    .B1(_06012_),
    .Y(_01045_));
 sky130_fd_sc_hd__nand2_2 _26229_ (.A(net1564),
    .B(_05793_),
    .Y(_06013_));
 sky130_fd_sc_hd__nand2_1 _26230_ (.A(\gen_regfile_ff.register_file_i.rf_reg[89] ),
    .B(_05798_),
    .Y(_06014_));
 sky130_fd_sc_hd__nand2_1 _26231_ (.A(_06013_),
    .B(_06014_),
    .Y(_01046_));
 sky130_fd_sc_hd__mux2_1 _26232_ (.A0(_02113_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[612] ),
    .S(_06006_),
    .X(_01047_));
 sky130_fd_sc_hd__mux2_1 _26233_ (.A0(_02250_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[613] ),
    .S(_06006_),
    .X(_01048_));
 sky130_fd_sc_hd__mux2_1 _26234_ (.A0(_02360_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[614] ),
    .S(_06006_),
    .X(_01049_));
 sky130_fd_sc_hd__mux2_1 _26235_ (.A0(_02468_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[615] ),
    .S(_06006_),
    .X(_01050_));
 sky130_fd_sc_hd__mux2_1 _26236_ (.A0(_02553_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[616] ),
    .S(_06006_),
    .X(_01051_));
 sky130_fd_sc_hd__mux2_1 _26237_ (.A0(_02653_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[617] ),
    .S(_06006_),
    .X(_01052_));
 sky130_fd_sc_hd__mux2_1 _26238_ (.A0(_02761_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[618] ),
    .S(net1300),
    .X(_01053_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_97 ();
 sky130_fd_sc_hd__mux2_1 _26240_ (.A0(_02849_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[619] ),
    .S(net1300),
    .X(_01054_));
 sky130_fd_sc_hd__mux2_1 _26241_ (.A0(_02974_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[620] ),
    .S(_06006_),
    .X(_01055_));
 sky130_fd_sc_hd__mux2_1 _26242_ (.A0(_03080_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[621] ),
    .S(net1300),
    .X(_01056_));
 sky130_fd_sc_hd__nand2_4 _26243_ (.A(net1515),
    .B(_05793_),
    .Y(_06016_));
 sky130_fd_sc_hd__nand2_1 _26244_ (.A(\gen_regfile_ff.register_file_i.rf_reg[90] ),
    .B(_05798_),
    .Y(_06017_));
 sky130_fd_sc_hd__nand2_2 _26245_ (.A(_06016_),
    .B(_06017_),
    .Y(_01057_));
 sky130_fd_sc_hd__mux2_1 _26246_ (.A0(_03214_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[622] ),
    .S(_06006_),
    .X(_01058_));
 sky130_fd_sc_hd__mux2_1 _26247_ (.A0(_03348_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[623] ),
    .S(_06006_),
    .X(_01059_));
 sky130_fd_sc_hd__nand2_1 _26248_ (.A(\gen_regfile_ff.register_file_i.rf_reg[624] ),
    .B(net1300),
    .Y(_06018_));
 sky130_fd_sc_hd__o21ai_0 _26249_ (.A1(_03481_),
    .A2(net1300),
    .B1(_06018_),
    .Y(_01060_));
 sky130_fd_sc_hd__mux2_1 _26250_ (.A0(_03614_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[625] ),
    .S(_06006_),
    .X(_01061_));
 sky130_fd_sc_hd__mux2_1 _26251_ (.A0(_03739_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[626] ),
    .S(_06006_),
    .X(_01062_));
 sky130_fd_sc_hd__mux2_1 _26252_ (.A0(_03866_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[627] ),
    .S(_06006_),
    .X(_01063_));
 sky130_fd_sc_hd__mux2_4 _26253_ (.A0(net1537),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[628] ),
    .S(_06006_),
    .X(_01064_));
 sky130_fd_sc_hd__mux2_1 _26254_ (.A0(net1017),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[629] ),
    .S(net1300),
    .X(_01065_));
 sky130_fd_sc_hd__mux2_4 _26255_ (.A0(net1517),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[630] ),
    .S(_06006_),
    .X(_01066_));
 sky130_fd_sc_hd__mux2_4 _26256_ (.A0(net1504),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[631] ),
    .S(net1300),
    .X(_01067_));
 sky130_fd_sc_hd__nand2_2 _26257_ (.A(net1529),
    .B(_05793_),
    .Y(_06019_));
 sky130_fd_sc_hd__nand2_1 _26258_ (.A(\gen_regfile_ff.register_file_i.rf_reg[91] ),
    .B(_05798_),
    .Y(_06020_));
 sky130_fd_sc_hd__nand2_1 _26259_ (.A(_06019_),
    .B(_06020_),
    .Y(_01068_));
 sky130_fd_sc_hd__nand2_1 _26260_ (.A(_01916_),
    .B(_02250_),
    .Y(_06021_));
 sky130_fd_sc_hd__nand2_1 _26261_ (.A(\gen_regfile_ff.register_file_i.rf_reg[37] ),
    .B(_01921_),
    .Y(_06022_));
 sky130_fd_sc_hd__nand2_1 _26262_ (.A(_06021_),
    .B(_06022_),
    .Y(_01069_));
 sky130_fd_sc_hd__mux2_4 _26263_ (.A0(net1316),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[632] ),
    .S(_06006_),
    .X(_01070_));
 sky130_fd_sc_hd__mux2_1 _26264_ (.A0(net252),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[633] ),
    .S(_06006_),
    .X(_01071_));
 sky130_fd_sc_hd__mux2_1 _26265_ (.A0(net251),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[634] ),
    .S(_06006_),
    .X(_01072_));
 sky130_fd_sc_hd__mux2_1 _26266_ (.A0(net1533),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[635] ),
    .S(net1300),
    .X(_01073_));
 sky130_fd_sc_hd__mux2_4 _26267_ (.A0(net886),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[636] ),
    .S(_06006_),
    .X(_01074_));
 sky130_fd_sc_hd__nor2_1 _26268_ (.A(_05084_),
    .B(net1300),
    .Y(_06023_));
 sky130_fd_sc_hd__a22o_1 _26269_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[637] ),
    .A2(net1300),
    .B1(net1246),
    .B2(_06023_),
    .X(_01075_));
 sky130_fd_sc_hd__mux2_4 _26270_ (.A0(net1238),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[638] ),
    .S(net1300),
    .X(_01076_));
 sky130_fd_sc_hd__nor2_1 _26271_ (.A(_05264_),
    .B(net1300),
    .Y(_06024_));
 sky130_fd_sc_hd__a22o_1 _26272_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[639] ),
    .A2(net1300),
    .B1(_06024_),
    .B2(net652),
    .X(_01077_));
 sky130_fd_sc_hd__nand2_4 _26273_ (.A(net446),
    .B(_05955_),
    .Y(_06025_));
 sky130_fd_sc_hd__nor2_8 _26274_ (.A(_02117_),
    .B(_06025_),
    .Y(_06026_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_96 ();
 sky130_fd_sc_hd__nand2_1 _26276_ (.A(_01909_),
    .B(_06026_),
    .Y(_06028_));
 sky130_fd_sc_hd__nand3_4 _26277_ (.A(net446),
    .B(_05955_),
    .C(_02122_),
    .Y(_06029_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_95 ();
 sky130_fd_sc_hd__nand2_1 _26279_ (.A(\gen_regfile_ff.register_file_i.rf_reg[640] ),
    .B(_06029_),
    .Y(_06031_));
 sky130_fd_sc_hd__nand2_1 _26280_ (.A(_06028_),
    .B(_06031_),
    .Y(_01078_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_94 ();
 sky130_fd_sc_hd__nand2_1 _26282_ (.A(\gen_regfile_ff.register_file_i.rf_reg[641] ),
    .B(_06029_),
    .Y(_06033_));
 sky130_fd_sc_hd__o21ai_0 _26283_ (.A1(_05299_),
    .A2(_06029_),
    .B1(_06033_),
    .Y(_01079_));
 sky130_fd_sc_hd__mux2_4 _26284_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[92] ),
    .A1(net250),
    .S(_05793_),
    .X(_01080_));
 sky130_fd_sc_hd__nand2_1 _26285_ (.A(_05326_),
    .B(_06026_),
    .Y(_06034_));
 sky130_fd_sc_hd__nand2_1 _26286_ (.A(\gen_regfile_ff.register_file_i.rf_reg[642] ),
    .B(_06029_),
    .Y(_06035_));
 sky130_fd_sc_hd__nand2_1 _26287_ (.A(_06034_),
    .B(_06035_),
    .Y(_01081_));
 sky130_fd_sc_hd__nand2_1 _26288_ (.A(\gen_regfile_ff.register_file_i.rf_reg[643] ),
    .B(_06029_),
    .Y(_06036_));
 sky130_fd_sc_hd__o21ai_0 _26289_ (.A1(_05351_),
    .A2(_06029_),
    .B1(_06036_),
    .Y(_01082_));
 sky130_fd_sc_hd__nand2_1 _26290_ (.A(_02113_),
    .B(_06026_),
    .Y(_06037_));
 sky130_fd_sc_hd__nand2_1 _26291_ (.A(\gen_regfile_ff.register_file_i.rf_reg[644] ),
    .B(_06029_),
    .Y(_06038_));
 sky130_fd_sc_hd__nand2_1 _26292_ (.A(_06037_),
    .B(_06038_),
    .Y(_01083_));
 sky130_fd_sc_hd__nand2_1 _26293_ (.A(_02250_),
    .B(_06026_),
    .Y(_06039_));
 sky130_fd_sc_hd__nand2_1 _26294_ (.A(\gen_regfile_ff.register_file_i.rf_reg[645] ),
    .B(_06029_),
    .Y(_06040_));
 sky130_fd_sc_hd__nand2_1 _26295_ (.A(_06039_),
    .B(_06040_),
    .Y(_01084_));
 sky130_fd_sc_hd__nand2_1 _26296_ (.A(_02360_),
    .B(_06026_),
    .Y(_06041_));
 sky130_fd_sc_hd__nand2_1 _26297_ (.A(\gen_regfile_ff.register_file_i.rf_reg[646] ),
    .B(_06029_),
    .Y(_06042_));
 sky130_fd_sc_hd__nand2_1 _26298_ (.A(_06041_),
    .B(_06042_),
    .Y(_01085_));
 sky130_fd_sc_hd__nand2_1 _26299_ (.A(_02468_),
    .B(_06026_),
    .Y(_06043_));
 sky130_fd_sc_hd__nand2_1 _26300_ (.A(\gen_regfile_ff.register_file_i.rf_reg[647] ),
    .B(_06029_),
    .Y(_06044_));
 sky130_fd_sc_hd__nand2_1 _26301_ (.A(_06043_),
    .B(_06044_),
    .Y(_01086_));
 sky130_fd_sc_hd__nand2_1 _26302_ (.A(_02553_),
    .B(_06026_),
    .Y(_06045_));
 sky130_fd_sc_hd__nand2_1 _26303_ (.A(\gen_regfile_ff.register_file_i.rf_reg[648] ),
    .B(_06029_),
    .Y(_06046_));
 sky130_fd_sc_hd__nand2_1 _26304_ (.A(_06045_),
    .B(_06046_),
    .Y(_01087_));
 sky130_fd_sc_hd__nand2_1 _26305_ (.A(_02653_),
    .B(_06026_),
    .Y(_06047_));
 sky130_fd_sc_hd__nand2_1 _26306_ (.A(\gen_regfile_ff.register_file_i.rf_reg[649] ),
    .B(_06029_),
    .Y(_06048_));
 sky130_fd_sc_hd__nand2_1 _26307_ (.A(_06047_),
    .B(_06048_),
    .Y(_01088_));
 sky130_fd_sc_hd__nand2_1 _26308_ (.A(_02761_),
    .B(_06026_),
    .Y(_06049_));
 sky130_fd_sc_hd__nand2_1 _26309_ (.A(\gen_regfile_ff.register_file_i.rf_reg[650] ),
    .B(_06029_),
    .Y(_06050_));
 sky130_fd_sc_hd__nand2_1 _26310_ (.A(_06049_),
    .B(_06050_),
    .Y(_01089_));
 sky130_fd_sc_hd__nand2_1 _26311_ (.A(_02849_),
    .B(_06026_),
    .Y(_06051_));
 sky130_fd_sc_hd__nand2_1 _26312_ (.A(\gen_regfile_ff.register_file_i.rf_reg[651] ),
    .B(_06029_),
    .Y(_06052_));
 sky130_fd_sc_hd__nand2_1 _26313_ (.A(_06051_),
    .B(_06052_),
    .Y(_01090_));
 sky130_fd_sc_hd__nor2_1 _26314_ (.A(_05084_),
    .B(_05798_),
    .Y(_06053_));
 sky130_fd_sc_hd__a22o_1 _26315_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[93] ),
    .A2(_05798_),
    .B1(_05079_),
    .B2(_06053_),
    .X(_01091_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_93 ();
 sky130_fd_sc_hd__nand2_1 _26317_ (.A(_02974_),
    .B(_06026_),
    .Y(_06055_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_92 ();
 sky130_fd_sc_hd__nand2_1 _26319_ (.A(\gen_regfile_ff.register_file_i.rf_reg[652] ),
    .B(_06029_),
    .Y(_06057_));
 sky130_fd_sc_hd__nand2_1 _26320_ (.A(_06055_),
    .B(_06057_),
    .Y(_01092_));
 sky130_fd_sc_hd__nand2_1 _26321_ (.A(_03080_),
    .B(_06026_),
    .Y(_06058_));
 sky130_fd_sc_hd__nand2_1 _26322_ (.A(\gen_regfile_ff.register_file_i.rf_reg[653] ),
    .B(_06029_),
    .Y(_06059_));
 sky130_fd_sc_hd__nand2_1 _26323_ (.A(_06058_),
    .B(_06059_),
    .Y(_01093_));
 sky130_fd_sc_hd__nand2_1 _26324_ (.A(_03214_),
    .B(_06026_),
    .Y(_06060_));
 sky130_fd_sc_hd__nand2_1 _26325_ (.A(\gen_regfile_ff.register_file_i.rf_reg[654] ),
    .B(_06029_),
    .Y(_06061_));
 sky130_fd_sc_hd__nand2_1 _26326_ (.A(_06060_),
    .B(_06061_),
    .Y(_01094_));
 sky130_fd_sc_hd__nand2_1 _26327_ (.A(_03348_),
    .B(_06026_),
    .Y(_06062_));
 sky130_fd_sc_hd__nand2_1 _26328_ (.A(\gen_regfile_ff.register_file_i.rf_reg[655] ),
    .B(_06029_),
    .Y(_06063_));
 sky130_fd_sc_hd__nand2_1 _26329_ (.A(_06062_),
    .B(_06063_),
    .Y(_01095_));
 sky130_fd_sc_hd__nand2_1 _26330_ (.A(\gen_regfile_ff.register_file_i.rf_reg[656] ),
    .B(_06029_),
    .Y(_06064_));
 sky130_fd_sc_hd__o21ai_0 _26331_ (.A1(_03481_),
    .A2(_06029_),
    .B1(_06064_),
    .Y(_01096_));
 sky130_fd_sc_hd__nand2_1 _26332_ (.A(net1575),
    .B(_06026_),
    .Y(_06065_));
 sky130_fd_sc_hd__nand2_1 _26333_ (.A(\gen_regfile_ff.register_file_i.rf_reg[657] ),
    .B(_06029_),
    .Y(_06066_));
 sky130_fd_sc_hd__nand2_1 _26334_ (.A(_06065_),
    .B(_06066_),
    .Y(_01097_));
 sky130_fd_sc_hd__nand2_1 _26335_ (.A(_03739_),
    .B(_06026_),
    .Y(_06067_));
 sky130_fd_sc_hd__nand2_1 _26336_ (.A(\gen_regfile_ff.register_file_i.rf_reg[658] ),
    .B(_06029_),
    .Y(_06068_));
 sky130_fd_sc_hd__nand2_1 _26337_ (.A(_06067_),
    .B(_06068_),
    .Y(_01098_));
 sky130_fd_sc_hd__nand2_1 _26338_ (.A(net1551),
    .B(_06026_),
    .Y(_06069_));
 sky130_fd_sc_hd__nand2_1 _26339_ (.A(\gen_regfile_ff.register_file_i.rf_reg[659] ),
    .B(_06029_),
    .Y(_06070_));
 sky130_fd_sc_hd__nand2_1 _26340_ (.A(_06069_),
    .B(_06070_),
    .Y(_01099_));
 sky130_fd_sc_hd__nand2_1 _26341_ (.A(net1544),
    .B(_06026_),
    .Y(_06071_));
 sky130_fd_sc_hd__nand2_1 _26342_ (.A(\gen_regfile_ff.register_file_i.rf_reg[660] ),
    .B(_06029_),
    .Y(_06072_));
 sky130_fd_sc_hd__nand2_1 _26343_ (.A(_06071_),
    .B(_06072_),
    .Y(_01100_));
 sky130_fd_sc_hd__nand2_1 _26344_ (.A(net1584),
    .B(_06026_),
    .Y(_06073_));
 sky130_fd_sc_hd__nand2_1 _26345_ (.A(\gen_regfile_ff.register_file_i.rf_reg[661] ),
    .B(_06029_),
    .Y(_06074_));
 sky130_fd_sc_hd__nand2_1 _26346_ (.A(_06073_),
    .B(_06074_),
    .Y(_01101_));
 sky130_fd_sc_hd__mux2_4 _26347_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[94] ),
    .A1(net1237),
    .S(_05793_),
    .X(_01102_));
 sky130_fd_sc_hd__mux2_4 _26348_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[662] ),
    .A1(net1517),
    .S(_06026_),
    .X(_01103_));
 sky130_fd_sc_hd__nand2_2 _26349_ (.A(net1291),
    .B(_06026_),
    .Y(_06075_));
 sky130_fd_sc_hd__nand2_1 _26350_ (.A(\gen_regfile_ff.register_file_i.rf_reg[663] ),
    .B(_06029_),
    .Y(_06076_));
 sky130_fd_sc_hd__nand2_1 _26351_ (.A(_06075_),
    .B(_06076_),
    .Y(_01104_));
 sky130_fd_sc_hd__nand2_1 _26352_ (.A(net1541),
    .B(_06026_),
    .Y(_06077_));
 sky130_fd_sc_hd__nand2_1 _26353_ (.A(\gen_regfile_ff.register_file_i.rf_reg[664] ),
    .B(_06029_),
    .Y(_06078_));
 sky130_fd_sc_hd__nand2_1 _26354_ (.A(_06077_),
    .B(_06078_),
    .Y(_01105_));
 sky130_fd_sc_hd__nand2_1 _26355_ (.A(net1586),
    .B(_06026_),
    .Y(_06079_));
 sky130_fd_sc_hd__nand2_1 _26356_ (.A(\gen_regfile_ff.register_file_i.rf_reg[665] ),
    .B(_06029_),
    .Y(_06080_));
 sky130_fd_sc_hd__nand2_1 _26357_ (.A(_06079_),
    .B(_06080_),
    .Y(_01106_));
 sky130_fd_sc_hd__nand2_1 _26358_ (.A(net1536),
    .B(_06026_),
    .Y(_06081_));
 sky130_fd_sc_hd__nand2_1 _26359_ (.A(\gen_regfile_ff.register_file_i.rf_reg[666] ),
    .B(_06029_),
    .Y(_06082_));
 sky130_fd_sc_hd__nand2_1 _26360_ (.A(_06081_),
    .B(_06082_),
    .Y(_01107_));
 sky130_fd_sc_hd__nand2_2 _26361_ (.A(net1542),
    .B(_06026_),
    .Y(_06083_));
 sky130_fd_sc_hd__nand2_1 _26362_ (.A(\gen_regfile_ff.register_file_i.rf_reg[667] ),
    .B(_06029_),
    .Y(_06084_));
 sky130_fd_sc_hd__nand2_1 _26363_ (.A(_06083_),
    .B(_06084_),
    .Y(_01108_));
 sky130_fd_sc_hd__mux2_4 _26364_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[668] ),
    .A1(net886),
    .S(_06026_),
    .X(_01109_));
 sky130_fd_sc_hd__nor2_1 _26365_ (.A(_05084_),
    .B(_06029_),
    .Y(_06085_));
 sky130_fd_sc_hd__a22o_1 _26366_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[669] ),
    .A2(_06029_),
    .B1(net1246),
    .B2(_06085_),
    .X(_01110_));
 sky130_fd_sc_hd__mux2_4 _26367_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[670] ),
    .A1(net1238),
    .S(_06026_),
    .X(_01111_));
 sky130_fd_sc_hd__nor2_1 _26368_ (.A(_05264_),
    .B(_06029_),
    .Y(_06086_));
 sky130_fd_sc_hd__a22o_1 _26369_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[671] ),
    .A2(_06029_),
    .B1(_06086_),
    .B2(net740),
    .X(_01112_));
 sky130_fd_sc_hd__nor2_1 _26370_ (.A(_05264_),
    .B(_05798_),
    .Y(_06087_));
 sky130_fd_sc_hd__a22o_1 _26371_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[95] ),
    .A2(_05798_),
    .B1(net740),
    .B2(_06087_),
    .X(_01113_));
 sky130_fd_sc_hd__nand2_4 _26372_ (.A(net446),
    .B(_01919_),
    .Y(_06088_));
 sky130_fd_sc_hd__nor2_8 _26373_ (.A(_02117_),
    .B(_06088_),
    .Y(_06089_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_91 ();
 sky130_fd_sc_hd__nand2_1 _26375_ (.A(_01909_),
    .B(_06089_),
    .Y(_06091_));
 sky130_fd_sc_hd__nand3_4 _26376_ (.A(net446),
    .B(_01919_),
    .C(_02122_),
    .Y(_06092_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_90 ();
 sky130_fd_sc_hd__nand2_1 _26378_ (.A(\gen_regfile_ff.register_file_i.rf_reg[672] ),
    .B(_06092_),
    .Y(_06094_));
 sky130_fd_sc_hd__nand2_1 _26379_ (.A(_06091_),
    .B(_06094_),
    .Y(_01114_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_89 ();
 sky130_fd_sc_hd__nand2_1 _26381_ (.A(\gen_regfile_ff.register_file_i.rf_reg[673] ),
    .B(_06092_),
    .Y(_06096_));
 sky130_fd_sc_hd__o21ai_0 _26382_ (.A1(_05299_),
    .A2(_06092_),
    .B1(_06096_),
    .Y(_01115_));
 sky130_fd_sc_hd__nand2_1 _26383_ (.A(_05326_),
    .B(_06089_),
    .Y(_06097_));
 sky130_fd_sc_hd__nand2_1 _26384_ (.A(\gen_regfile_ff.register_file_i.rf_reg[674] ),
    .B(_06092_),
    .Y(_06098_));
 sky130_fd_sc_hd__nand2_1 _26385_ (.A(_06097_),
    .B(_06098_),
    .Y(_01116_));
 sky130_fd_sc_hd__nand2_1 _26386_ (.A(\gen_regfile_ff.register_file_i.rf_reg[675] ),
    .B(_06092_),
    .Y(_06099_));
 sky130_fd_sc_hd__o21ai_0 _26387_ (.A1(_05351_),
    .A2(_06092_),
    .B1(_06099_),
    .Y(_01117_));
 sky130_fd_sc_hd__nand2_1 _26388_ (.A(_02113_),
    .B(_06089_),
    .Y(_06100_));
 sky130_fd_sc_hd__nand2_1 _26389_ (.A(\gen_regfile_ff.register_file_i.rf_reg[676] ),
    .B(_06092_),
    .Y(_06101_));
 sky130_fd_sc_hd__nand2_1 _26390_ (.A(_06100_),
    .B(_06101_),
    .Y(_01118_));
 sky130_fd_sc_hd__nand2_1 _26391_ (.A(_02250_),
    .B(_06089_),
    .Y(_06102_));
 sky130_fd_sc_hd__nand2_1 _26392_ (.A(\gen_regfile_ff.register_file_i.rf_reg[677] ),
    .B(_06092_),
    .Y(_06103_));
 sky130_fd_sc_hd__nand2_1 _26393_ (.A(_06102_),
    .B(_06103_),
    .Y(_01119_));
 sky130_fd_sc_hd__nand2_1 _26394_ (.A(_02360_),
    .B(_06089_),
    .Y(_06104_));
 sky130_fd_sc_hd__nand2_1 _26395_ (.A(\gen_regfile_ff.register_file_i.rf_reg[678] ),
    .B(_06092_),
    .Y(_06105_));
 sky130_fd_sc_hd__nand2_1 _26396_ (.A(_06104_),
    .B(_06105_),
    .Y(_01120_));
 sky130_fd_sc_hd__nand2_1 _26397_ (.A(_02468_),
    .B(_06089_),
    .Y(_06106_));
 sky130_fd_sc_hd__nand2_1 _26398_ (.A(\gen_regfile_ff.register_file_i.rf_reg[679] ),
    .B(_06092_),
    .Y(_06107_));
 sky130_fd_sc_hd__nand2_1 _26399_ (.A(_06106_),
    .B(_06107_),
    .Y(_01121_));
 sky130_fd_sc_hd__nand2_1 _26400_ (.A(_02553_),
    .B(_06089_),
    .Y(_06108_));
 sky130_fd_sc_hd__nand2_1 _26401_ (.A(\gen_regfile_ff.register_file_i.rf_reg[680] ),
    .B(_06092_),
    .Y(_06109_));
 sky130_fd_sc_hd__nand2_1 _26402_ (.A(_06108_),
    .B(_06109_),
    .Y(_01122_));
 sky130_fd_sc_hd__nand2_1 _26403_ (.A(_02653_),
    .B(_06089_),
    .Y(_06110_));
 sky130_fd_sc_hd__nand2_1 _26404_ (.A(\gen_regfile_ff.register_file_i.rf_reg[681] ),
    .B(_06092_),
    .Y(_06111_));
 sky130_fd_sc_hd__nand2_1 _26405_ (.A(_06110_),
    .B(_06111_),
    .Y(_01123_));
 sky130_fd_sc_hd__nor2_8 _26406_ (.A(_01913_),
    .B(_05501_),
    .Y(_06112_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_88 ();
 sky130_fd_sc_hd__nand2_1 _26408_ (.A(_01909_),
    .B(_06112_),
    .Y(_06114_));
 sky130_fd_sc_hd__nand3_4 _26409_ (.A(net1021),
    .B(net331),
    .C(_01918_),
    .Y(_06115_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_87 ();
 sky130_fd_sc_hd__nand2_1 _26411_ (.A(\gen_regfile_ff.register_file_i.rf_reg[96] ),
    .B(_06115_),
    .Y(_06117_));
 sky130_fd_sc_hd__nand2_1 _26412_ (.A(_06114_),
    .B(_06117_),
    .Y(_01124_));
 sky130_fd_sc_hd__nand2_1 _26413_ (.A(_02761_),
    .B(_06089_),
    .Y(_06118_));
 sky130_fd_sc_hd__nand2_1 _26414_ (.A(\gen_regfile_ff.register_file_i.rf_reg[682] ),
    .B(_06092_),
    .Y(_06119_));
 sky130_fd_sc_hd__nand2_1 _26415_ (.A(_06118_),
    .B(_06119_),
    .Y(_01125_));
 sky130_fd_sc_hd__nand2_1 _26416_ (.A(_02849_),
    .B(_06089_),
    .Y(_06120_));
 sky130_fd_sc_hd__nand2_1 _26417_ (.A(\gen_regfile_ff.register_file_i.rf_reg[683] ),
    .B(_06092_),
    .Y(_06121_));
 sky130_fd_sc_hd__nand2_1 _26418_ (.A(_06120_),
    .B(_06121_),
    .Y(_01126_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_86 ();
 sky130_fd_sc_hd__nand2_1 _26420_ (.A(_02974_),
    .B(_06089_),
    .Y(_06123_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_85 ();
 sky130_fd_sc_hd__nand2_1 _26422_ (.A(\gen_regfile_ff.register_file_i.rf_reg[684] ),
    .B(_06092_),
    .Y(_06125_));
 sky130_fd_sc_hd__nand2_1 _26423_ (.A(_06123_),
    .B(_06125_),
    .Y(_01127_));
 sky130_fd_sc_hd__nand2_1 _26424_ (.A(_03080_),
    .B(_06089_),
    .Y(_06126_));
 sky130_fd_sc_hd__nand2_1 _26425_ (.A(\gen_regfile_ff.register_file_i.rf_reg[685] ),
    .B(_06092_),
    .Y(_06127_));
 sky130_fd_sc_hd__nand2_1 _26426_ (.A(_06126_),
    .B(_06127_),
    .Y(_01128_));
 sky130_fd_sc_hd__nand2_1 _26427_ (.A(_03214_),
    .B(_06089_),
    .Y(_06128_));
 sky130_fd_sc_hd__nand2_1 _26428_ (.A(\gen_regfile_ff.register_file_i.rf_reg[686] ),
    .B(_06092_),
    .Y(_06129_));
 sky130_fd_sc_hd__nand2_1 _26429_ (.A(_06128_),
    .B(_06129_),
    .Y(_01129_));
 sky130_fd_sc_hd__nand2_1 _26430_ (.A(_03348_),
    .B(_06089_),
    .Y(_06130_));
 sky130_fd_sc_hd__nand2_1 _26431_ (.A(\gen_regfile_ff.register_file_i.rf_reg[687] ),
    .B(_06092_),
    .Y(_06131_));
 sky130_fd_sc_hd__nand2_1 _26432_ (.A(_06130_),
    .B(_06131_),
    .Y(_01130_));
 sky130_fd_sc_hd__nand2_1 _26433_ (.A(\gen_regfile_ff.register_file_i.rf_reg[688] ),
    .B(_06092_),
    .Y(_06132_));
 sky130_fd_sc_hd__o21ai_0 _26434_ (.A1(_03481_),
    .A2(_06092_),
    .B1(_06132_),
    .Y(_01131_));
 sky130_fd_sc_hd__nand2_1 _26435_ (.A(net1575),
    .B(_06089_),
    .Y(_06133_));
 sky130_fd_sc_hd__nand2_1 _26436_ (.A(\gen_regfile_ff.register_file_i.rf_reg[689] ),
    .B(_06092_),
    .Y(_06134_));
 sky130_fd_sc_hd__nand2_1 _26437_ (.A(_06133_),
    .B(_06134_),
    .Y(_01132_));
 sky130_fd_sc_hd__nand2_1 _26438_ (.A(_03739_),
    .B(_06089_),
    .Y(_06135_));
 sky130_fd_sc_hd__nand2_1 _26439_ (.A(\gen_regfile_ff.register_file_i.rf_reg[690] ),
    .B(_06092_),
    .Y(_06136_));
 sky130_fd_sc_hd__nand2_1 _26440_ (.A(_06135_),
    .B(_06136_),
    .Y(_01133_));
 sky130_fd_sc_hd__nand2_1 _26441_ (.A(_03866_),
    .B(_06089_),
    .Y(_06137_));
 sky130_fd_sc_hd__nand2_1 _26442_ (.A(\gen_regfile_ff.register_file_i.rf_reg[691] ),
    .B(_06092_),
    .Y(_06138_));
 sky130_fd_sc_hd__nand2_1 _26443_ (.A(_06137_),
    .B(_06138_),
    .Y(_01134_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_83 ();
 sky130_fd_sc_hd__nand2_1 _26446_ (.A(\gen_regfile_ff.register_file_i.rf_reg[97] ),
    .B(_06115_),
    .Y(_06141_));
 sky130_fd_sc_hd__o21ai_0 _26447_ (.A1(_05299_),
    .A2(_06115_),
    .B1(_06141_),
    .Y(_01135_));
 sky130_fd_sc_hd__nand2_1 _26448_ (.A(_03982_),
    .B(_06089_),
    .Y(_06142_));
 sky130_fd_sc_hd__nand2_1 _26449_ (.A(\gen_regfile_ff.register_file_i.rf_reg[692] ),
    .B(_06092_),
    .Y(_06143_));
 sky130_fd_sc_hd__nand2_1 _26450_ (.A(_06142_),
    .B(_06143_),
    .Y(_01136_));
 sky130_fd_sc_hd__nand2_1 _26451_ (.A(net1584),
    .B(_06089_),
    .Y(_06144_));
 sky130_fd_sc_hd__nand2_1 _26452_ (.A(\gen_regfile_ff.register_file_i.rf_reg[693] ),
    .B(_06092_),
    .Y(_06145_));
 sky130_fd_sc_hd__nand2_1 _26453_ (.A(_06144_),
    .B(_06145_),
    .Y(_01137_));
 sky130_fd_sc_hd__mux2_4 _26454_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[694] ),
    .A1(net1517),
    .S(_06089_),
    .X(_01138_));
 sky130_fd_sc_hd__nand2_4 _26455_ (.A(net1291),
    .B(_06089_),
    .Y(_06146_));
 sky130_fd_sc_hd__nand2_1 _26456_ (.A(\gen_regfile_ff.register_file_i.rf_reg[695] ),
    .B(_06092_),
    .Y(_06147_));
 sky130_fd_sc_hd__nand2_2 _26457_ (.A(_06147_),
    .B(_06146_),
    .Y(_01139_));
 sky130_fd_sc_hd__nand2_1 _26458_ (.A(net1541),
    .B(_06089_),
    .Y(_06148_));
 sky130_fd_sc_hd__nand2_1 _26459_ (.A(\gen_regfile_ff.register_file_i.rf_reg[696] ),
    .B(_06092_),
    .Y(_06149_));
 sky130_fd_sc_hd__nand2_1 _26460_ (.A(_06148_),
    .B(_06149_),
    .Y(_01140_));
 sky130_fd_sc_hd__nand2_1 _26461_ (.A(net1586),
    .B(_06089_),
    .Y(_06150_));
 sky130_fd_sc_hd__nand2_1 _26462_ (.A(\gen_regfile_ff.register_file_i.rf_reg[697] ),
    .B(_06092_),
    .Y(_06151_));
 sky130_fd_sc_hd__nand2_1 _26463_ (.A(_06150_),
    .B(_06151_),
    .Y(_01141_));
 sky130_fd_sc_hd__nand2_4 _26464_ (.A(net1514),
    .B(_06089_),
    .Y(_06152_));
 sky130_fd_sc_hd__nand2_1 _26465_ (.A(\gen_regfile_ff.register_file_i.rf_reg[698] ),
    .B(_06092_),
    .Y(_06153_));
 sky130_fd_sc_hd__nand2_2 _26466_ (.A(_06152_),
    .B(_06153_),
    .Y(_01142_));
 sky130_fd_sc_hd__nand2_2 _26467_ (.A(net1542),
    .B(_06089_),
    .Y(_06154_));
 sky130_fd_sc_hd__nand2_1 _26468_ (.A(\gen_regfile_ff.register_file_i.rf_reg[699] ),
    .B(_06092_),
    .Y(_06155_));
 sky130_fd_sc_hd__nand2_1 _26469_ (.A(_06154_),
    .B(_06155_),
    .Y(_01143_));
 sky130_fd_sc_hd__mux2_4 _26470_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[700] ),
    .A1(net885),
    .S(_06089_),
    .X(_01144_));
 sky130_fd_sc_hd__nor2_1 _26471_ (.A(_05084_),
    .B(_06092_),
    .Y(_06156_));
 sky130_fd_sc_hd__a22o_1 _26472_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[701] ),
    .A2(_06092_),
    .B1(net1254),
    .B2(_06156_),
    .X(_01145_));
 sky130_fd_sc_hd__nand2_1 _26473_ (.A(_05326_),
    .B(_06112_),
    .Y(_06157_));
 sky130_fd_sc_hd__nand2_1 _26474_ (.A(\gen_regfile_ff.register_file_i.rf_reg[98] ),
    .B(_06115_),
    .Y(_06158_));
 sky130_fd_sc_hd__nand2_1 _26475_ (.A(_06157_),
    .B(_06158_),
    .Y(_01146_));
 sky130_fd_sc_hd__mux2_4 _26476_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[702] ),
    .A1(net1238),
    .S(_06089_),
    .X(_01147_));
 sky130_fd_sc_hd__nor2_1 _26477_ (.A(_05264_),
    .B(_06092_),
    .Y(_06159_));
 sky130_fd_sc_hd__a22o_1 _26478_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[703] ),
    .A2(_06092_),
    .B1(_06159_),
    .B2(net652),
    .X(_01148_));
 sky130_fd_sc_hd__nand2_4 _26479_ (.A(net446),
    .B(_05796_),
    .Y(_06160_));
 sky130_fd_sc_hd__nor2_8 _26480_ (.A(_02117_),
    .B(_06160_),
    .Y(_06161_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_82 ();
 sky130_fd_sc_hd__nand2_1 _26482_ (.A(_01909_),
    .B(_06161_),
    .Y(_06163_));
 sky130_fd_sc_hd__nand3_4 _26483_ (.A(net446),
    .B(_02122_),
    .C(_05796_),
    .Y(_06164_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_81 ();
 sky130_fd_sc_hd__nand2_1 _26485_ (.A(\gen_regfile_ff.register_file_i.rf_reg[704] ),
    .B(_06164_),
    .Y(_06166_));
 sky130_fd_sc_hd__nand2_1 _26486_ (.A(_06163_),
    .B(_06166_),
    .Y(_01149_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_80 ();
 sky130_fd_sc_hd__nand2_1 _26488_ (.A(\gen_regfile_ff.register_file_i.rf_reg[705] ),
    .B(_06164_),
    .Y(_06168_));
 sky130_fd_sc_hd__o21ai_0 _26489_ (.A1(_05299_),
    .A2(_06164_),
    .B1(_06168_),
    .Y(_01150_));
 sky130_fd_sc_hd__nand2_1 _26490_ (.A(_05326_),
    .B(_06161_),
    .Y(_06169_));
 sky130_fd_sc_hd__nand2_1 _26491_ (.A(\gen_regfile_ff.register_file_i.rf_reg[706] ),
    .B(_06164_),
    .Y(_06170_));
 sky130_fd_sc_hd__nand2_1 _26492_ (.A(_06169_),
    .B(_06170_),
    .Y(_01151_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_79 ();
 sky130_fd_sc_hd__nand2_1 _26494_ (.A(\gen_regfile_ff.register_file_i.rf_reg[707] ),
    .B(_06164_),
    .Y(_06172_));
 sky130_fd_sc_hd__o21ai_0 _26495_ (.A1(_05351_),
    .A2(_06164_),
    .B1(_06172_),
    .Y(_01152_));
 sky130_fd_sc_hd__nand2_1 _26496_ (.A(_02113_),
    .B(_06161_),
    .Y(_06173_));
 sky130_fd_sc_hd__nand2_1 _26497_ (.A(\gen_regfile_ff.register_file_i.rf_reg[708] ),
    .B(_06164_),
    .Y(_06174_));
 sky130_fd_sc_hd__nand2_1 _26498_ (.A(_06173_),
    .B(_06174_),
    .Y(_01153_));
 sky130_fd_sc_hd__nand2_1 _26499_ (.A(_02250_),
    .B(_06161_),
    .Y(_06175_));
 sky130_fd_sc_hd__nand2_1 _26500_ (.A(\gen_regfile_ff.register_file_i.rf_reg[709] ),
    .B(_06164_),
    .Y(_06176_));
 sky130_fd_sc_hd__nand2_1 _26501_ (.A(_06175_),
    .B(_06176_),
    .Y(_01154_));
 sky130_fd_sc_hd__nand2_1 _26502_ (.A(_02360_),
    .B(_06161_),
    .Y(_06177_));
 sky130_fd_sc_hd__nand2_1 _26503_ (.A(\gen_regfile_ff.register_file_i.rf_reg[710] ),
    .B(_06164_),
    .Y(_06178_));
 sky130_fd_sc_hd__nand2_1 _26504_ (.A(_06177_),
    .B(_06178_),
    .Y(_01155_));
 sky130_fd_sc_hd__nand2_1 _26505_ (.A(_02468_),
    .B(_06161_),
    .Y(_06179_));
 sky130_fd_sc_hd__nand2_1 _26506_ (.A(\gen_regfile_ff.register_file_i.rf_reg[711] ),
    .B(_06164_),
    .Y(_06180_));
 sky130_fd_sc_hd__nand2_1 _26507_ (.A(_06179_),
    .B(_06180_),
    .Y(_01156_));
 sky130_fd_sc_hd__nand2_1 _26508_ (.A(\gen_regfile_ff.register_file_i.rf_reg[99] ),
    .B(_06115_),
    .Y(_06181_));
 sky130_fd_sc_hd__o21ai_0 _26509_ (.A1(_05351_),
    .A2(_06115_),
    .B1(_06181_),
    .Y(_01157_));
 sky130_fd_sc_hd__nand2_1 _26510_ (.A(_02553_),
    .B(_06161_),
    .Y(_06182_));
 sky130_fd_sc_hd__nand2_1 _26511_ (.A(\gen_regfile_ff.register_file_i.rf_reg[712] ),
    .B(_06164_),
    .Y(_06183_));
 sky130_fd_sc_hd__nand2_1 _26512_ (.A(_06182_),
    .B(_06183_),
    .Y(_01158_));
 sky130_fd_sc_hd__nand2_1 _26513_ (.A(_02653_),
    .B(_06161_),
    .Y(_06184_));
 sky130_fd_sc_hd__nand2_1 _26514_ (.A(\gen_regfile_ff.register_file_i.rf_reg[713] ),
    .B(_06164_),
    .Y(_06185_));
 sky130_fd_sc_hd__nand2_1 _26515_ (.A(_06184_),
    .B(_06185_),
    .Y(_01159_));
 sky130_fd_sc_hd__nand2_1 _26516_ (.A(_02761_),
    .B(_06161_),
    .Y(_06186_));
 sky130_fd_sc_hd__nand2_1 _26517_ (.A(\gen_regfile_ff.register_file_i.rf_reg[714] ),
    .B(_06164_),
    .Y(_06187_));
 sky130_fd_sc_hd__nand2_1 _26518_ (.A(_06186_),
    .B(_06187_),
    .Y(_01160_));
 sky130_fd_sc_hd__nand2_1 _26519_ (.A(_02849_),
    .B(_06161_),
    .Y(_06188_));
 sky130_fd_sc_hd__nand2_1 _26520_ (.A(\gen_regfile_ff.register_file_i.rf_reg[715] ),
    .B(_06164_),
    .Y(_06189_));
 sky130_fd_sc_hd__nand2_1 _26521_ (.A(_06188_),
    .B(_06189_),
    .Y(_01161_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_78 ();
 sky130_fd_sc_hd__nand2_1 _26523_ (.A(_02974_),
    .B(_06161_),
    .Y(_06191_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_77 ();
 sky130_fd_sc_hd__nand2_1 _26525_ (.A(\gen_regfile_ff.register_file_i.rf_reg[716] ),
    .B(_06164_),
    .Y(_06193_));
 sky130_fd_sc_hd__nand2_1 _26526_ (.A(_06191_),
    .B(_06193_),
    .Y(_01162_));
 sky130_fd_sc_hd__nand2_1 _26527_ (.A(_03080_),
    .B(_06161_),
    .Y(_06194_));
 sky130_fd_sc_hd__nand2_1 _26528_ (.A(\gen_regfile_ff.register_file_i.rf_reg[717] ),
    .B(_06164_),
    .Y(_06195_));
 sky130_fd_sc_hd__nand2_1 _26529_ (.A(_06194_),
    .B(_06195_),
    .Y(_01163_));
 sky130_fd_sc_hd__nand2_1 _26530_ (.A(_03214_),
    .B(_06161_),
    .Y(_06196_));
 sky130_fd_sc_hd__nand2_1 _26531_ (.A(\gen_regfile_ff.register_file_i.rf_reg[718] ),
    .B(_06164_),
    .Y(_06197_));
 sky130_fd_sc_hd__nand2_1 _26532_ (.A(_06196_),
    .B(_06197_),
    .Y(_01164_));
 sky130_fd_sc_hd__nand2_1 _26533_ (.A(_03348_),
    .B(_06161_),
    .Y(_06198_));
 sky130_fd_sc_hd__nand2_1 _26534_ (.A(\gen_regfile_ff.register_file_i.rf_reg[719] ),
    .B(_06164_),
    .Y(_06199_));
 sky130_fd_sc_hd__nand2_1 _26535_ (.A(_06198_),
    .B(_06199_),
    .Y(_01165_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_76 ();
 sky130_fd_sc_hd__nand2_1 _26537_ (.A(\gen_regfile_ff.register_file_i.rf_reg[720] ),
    .B(_06164_),
    .Y(_06201_));
 sky130_fd_sc_hd__o21ai_0 _26538_ (.A1(_03481_),
    .A2(_06164_),
    .B1(_06201_),
    .Y(_01166_));
 sky130_fd_sc_hd__nand2_1 _26539_ (.A(net1575),
    .B(_06161_),
    .Y(_06202_));
 sky130_fd_sc_hd__nand2_1 _26540_ (.A(\gen_regfile_ff.register_file_i.rf_reg[721] ),
    .B(_06164_),
    .Y(_06203_));
 sky130_fd_sc_hd__nand2_1 _26541_ (.A(_06202_),
    .B(_06203_),
    .Y(_01167_));
 sky130_fd_sc_hd__nand2_1 _26542_ (.A(_02113_),
    .B(_06112_),
    .Y(_06204_));
 sky130_fd_sc_hd__nand2_1 _26543_ (.A(\gen_regfile_ff.register_file_i.rf_reg[100] ),
    .B(_06115_),
    .Y(_06205_));
 sky130_fd_sc_hd__nand2_1 _26544_ (.A(_06204_),
    .B(_06205_),
    .Y(_01168_));
 sky130_fd_sc_hd__nand2_1 _26545_ (.A(net1576),
    .B(_06161_),
    .Y(_06206_));
 sky130_fd_sc_hd__nand2_1 _26546_ (.A(\gen_regfile_ff.register_file_i.rf_reg[722] ),
    .B(_06164_),
    .Y(_06207_));
 sky130_fd_sc_hd__nand2_1 _26547_ (.A(_06206_),
    .B(_06207_),
    .Y(_01169_));
 sky130_fd_sc_hd__nand2_1 _26548_ (.A(net1551),
    .B(_06161_),
    .Y(_06208_));
 sky130_fd_sc_hd__nand2_1 _26549_ (.A(\gen_regfile_ff.register_file_i.rf_reg[723] ),
    .B(_06164_),
    .Y(_06209_));
 sky130_fd_sc_hd__nand2_1 _26550_ (.A(_06208_),
    .B(_06209_),
    .Y(_01170_));
 sky130_fd_sc_hd__nand2_1 _26551_ (.A(net1544),
    .B(_06161_),
    .Y(_06210_));
 sky130_fd_sc_hd__nand2_1 _26552_ (.A(\gen_regfile_ff.register_file_i.rf_reg[724] ),
    .B(_06164_),
    .Y(_06211_));
 sky130_fd_sc_hd__nand2_1 _26553_ (.A(_06210_),
    .B(_06211_),
    .Y(_01171_));
 sky130_fd_sc_hd__nand2_1 _26554_ (.A(net1584),
    .B(_06161_),
    .Y(_06212_));
 sky130_fd_sc_hd__nand2_1 _26555_ (.A(\gen_regfile_ff.register_file_i.rf_reg[725] ),
    .B(_06164_),
    .Y(_06213_));
 sky130_fd_sc_hd__nand2_1 _26556_ (.A(_06212_),
    .B(_06213_),
    .Y(_01172_));
 sky130_fd_sc_hd__mux2_4 _26557_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[726] ),
    .A1(net1326),
    .S(_06161_),
    .X(_01173_));
 sky130_fd_sc_hd__nand2_2 _26558_ (.A(net1291),
    .B(_06161_),
    .Y(_06214_));
 sky130_fd_sc_hd__nand2_1 _26559_ (.A(\gen_regfile_ff.register_file_i.rf_reg[727] ),
    .B(_06164_),
    .Y(_06215_));
 sky130_fd_sc_hd__nand2_1 _26560_ (.A(_06214_),
    .B(_06215_),
    .Y(_01174_));
 sky130_fd_sc_hd__nand2_1 _26561_ (.A(net1541),
    .B(_06161_),
    .Y(_06216_));
 sky130_fd_sc_hd__nand2_1 _26562_ (.A(\gen_regfile_ff.register_file_i.rf_reg[728] ),
    .B(_06164_),
    .Y(_06217_));
 sky130_fd_sc_hd__nand2_1 _26563_ (.A(_06216_),
    .B(_06217_),
    .Y(_01175_));
 sky130_fd_sc_hd__nand2_1 _26564_ (.A(net1586),
    .B(_06161_),
    .Y(_06218_));
 sky130_fd_sc_hd__nand2_1 _26565_ (.A(\gen_regfile_ff.register_file_i.rf_reg[729] ),
    .B(_06164_),
    .Y(_06219_));
 sky130_fd_sc_hd__nand2_1 _26566_ (.A(_06218_),
    .B(_06219_),
    .Y(_01176_));
 sky130_fd_sc_hd__nand2_2 _26567_ (.A(net1514),
    .B(_06161_),
    .Y(_06220_));
 sky130_fd_sc_hd__nand2_1 _26568_ (.A(\gen_regfile_ff.register_file_i.rf_reg[730] ),
    .B(_06164_),
    .Y(_06221_));
 sky130_fd_sc_hd__nand2_1 _26569_ (.A(_06220_),
    .B(_06221_),
    .Y(_01177_));
 sky130_fd_sc_hd__nand2_2 _26570_ (.A(net1542),
    .B(_06161_),
    .Y(_06222_));
 sky130_fd_sc_hd__nand2_1 _26571_ (.A(\gen_regfile_ff.register_file_i.rf_reg[731] ),
    .B(_06164_),
    .Y(_06223_));
 sky130_fd_sc_hd__nand2_1 _26572_ (.A(_06222_),
    .B(_06223_),
    .Y(_01178_));
 sky130_fd_sc_hd__nand2_1 _26573_ (.A(_02250_),
    .B(_06112_),
    .Y(_06224_));
 sky130_fd_sc_hd__nand2_1 _26574_ (.A(\gen_regfile_ff.register_file_i.rf_reg[101] ),
    .B(_06115_),
    .Y(_06225_));
 sky130_fd_sc_hd__nand2_1 _26575_ (.A(_06224_),
    .B(_06225_),
    .Y(_01179_));
 sky130_fd_sc_hd__nand2_1 _26576_ (.A(_01916_),
    .B(_02360_),
    .Y(_06226_));
 sky130_fd_sc_hd__nand2_1 _26577_ (.A(\gen_regfile_ff.register_file_i.rf_reg[38] ),
    .B(_01921_),
    .Y(_06227_));
 sky130_fd_sc_hd__nand2_1 _26578_ (.A(_06226_),
    .B(_06227_),
    .Y(_01180_));
 sky130_fd_sc_hd__mux2_4 _26579_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[732] ),
    .A1(net1294),
    .S(_06161_),
    .X(_01181_));
 sky130_fd_sc_hd__nor2_1 _26580_ (.A(_05084_),
    .B(_06164_),
    .Y(_06228_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_75 ();
 sky130_fd_sc_hd__a22o_1 _26582_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[733] ),
    .A2(_06164_),
    .B1(net1249),
    .B2(_06228_),
    .X(_01182_));
 sky130_fd_sc_hd__mux2_4 _26583_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[734] ),
    .A1(net1237),
    .S(_06161_),
    .X(_01183_));
 sky130_fd_sc_hd__nor2_1 _26584_ (.A(_05264_),
    .B(_06164_),
    .Y(_06230_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_74 ();
 sky130_fd_sc_hd__a22o_1 _26586_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[735] ),
    .A2(_06164_),
    .B1(_06230_),
    .B2(net500),
    .X(_01184_));
 sky130_fd_sc_hd__nand3_4 _26587_ (.A(net1020),
    .B(net331),
    .C(net446),
    .Y(_06232_));
 sky130_fd_sc_hd__nor2_8 _26588_ (.A(_02117_),
    .B(_06232_),
    .Y(_06233_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_73 ();
 sky130_fd_sc_hd__nand2_1 _26590_ (.A(_01909_),
    .B(_06233_),
    .Y(_06235_));
 sky130_fd_sc_hd__and3_4 _26591_ (.A(net1021),
    .B(net331),
    .C(net446),
    .X(_06236_));
 sky130_fd_sc_hd__nand2_8 _26592_ (.A(_02122_),
    .B(_06236_),
    .Y(_06237_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_72 ();
 sky130_fd_sc_hd__nand2_1 _26594_ (.A(\gen_regfile_ff.register_file_i.rf_reg[736] ),
    .B(_06237_),
    .Y(_06239_));
 sky130_fd_sc_hd__nand2_1 _26595_ (.A(_06235_),
    .B(_06239_),
    .Y(_01185_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_71 ();
 sky130_fd_sc_hd__nand2_1 _26597_ (.A(\gen_regfile_ff.register_file_i.rf_reg[737] ),
    .B(_06237_),
    .Y(_06241_));
 sky130_fd_sc_hd__o21ai_0 _26598_ (.A1(_05299_),
    .A2(_06237_),
    .B1(_06241_),
    .Y(_01186_));
 sky130_fd_sc_hd__nand2_1 _26599_ (.A(_05326_),
    .B(_06233_),
    .Y(_06242_));
 sky130_fd_sc_hd__nand2_1 _26600_ (.A(\gen_regfile_ff.register_file_i.rf_reg[738] ),
    .B(_06237_),
    .Y(_06243_));
 sky130_fd_sc_hd__nand2_1 _26601_ (.A(_06242_),
    .B(_06243_),
    .Y(_01187_));
 sky130_fd_sc_hd__nand2_1 _26602_ (.A(\gen_regfile_ff.register_file_i.rf_reg[739] ),
    .B(_06237_),
    .Y(_06244_));
 sky130_fd_sc_hd__o21ai_0 _26603_ (.A1(_05351_),
    .A2(_06237_),
    .B1(_06244_),
    .Y(_01188_));
 sky130_fd_sc_hd__nand2_1 _26604_ (.A(_02113_),
    .B(_06233_),
    .Y(_06245_));
 sky130_fd_sc_hd__nand2_1 _26605_ (.A(\gen_regfile_ff.register_file_i.rf_reg[740] ),
    .B(_06237_),
    .Y(_06246_));
 sky130_fd_sc_hd__nand2_1 _26606_ (.A(_06245_),
    .B(_06246_),
    .Y(_01189_));
 sky130_fd_sc_hd__nand2_1 _26607_ (.A(_02250_),
    .B(_06233_),
    .Y(_06247_));
 sky130_fd_sc_hd__nand2_1 _26608_ (.A(\gen_regfile_ff.register_file_i.rf_reg[741] ),
    .B(_06237_),
    .Y(_06248_));
 sky130_fd_sc_hd__nand2_1 _26609_ (.A(_06247_),
    .B(_06248_),
    .Y(_01190_));
 sky130_fd_sc_hd__nand2_1 _26610_ (.A(_02360_),
    .B(_06112_),
    .Y(_06249_));
 sky130_fd_sc_hd__nand2_1 _26611_ (.A(\gen_regfile_ff.register_file_i.rf_reg[102] ),
    .B(_06115_),
    .Y(_06250_));
 sky130_fd_sc_hd__nand2_1 _26612_ (.A(_06249_),
    .B(_06250_),
    .Y(_01191_));
 sky130_fd_sc_hd__nand2_1 _26613_ (.A(_02360_),
    .B(_06233_),
    .Y(_06251_));
 sky130_fd_sc_hd__nand2_1 _26614_ (.A(\gen_regfile_ff.register_file_i.rf_reg[742] ),
    .B(_06237_),
    .Y(_06252_));
 sky130_fd_sc_hd__nand2_1 _26615_ (.A(_06251_),
    .B(_06252_),
    .Y(_01192_));
 sky130_fd_sc_hd__nand2_1 _26616_ (.A(_02468_),
    .B(_06233_),
    .Y(_06253_));
 sky130_fd_sc_hd__nand2_1 _26617_ (.A(\gen_regfile_ff.register_file_i.rf_reg[743] ),
    .B(_06237_),
    .Y(_06254_));
 sky130_fd_sc_hd__nand2_1 _26618_ (.A(_06253_),
    .B(_06254_),
    .Y(_01193_));
 sky130_fd_sc_hd__nand2_1 _26619_ (.A(_02553_),
    .B(_06233_),
    .Y(_06255_));
 sky130_fd_sc_hd__nand2_1 _26620_ (.A(\gen_regfile_ff.register_file_i.rf_reg[744] ),
    .B(_06237_),
    .Y(_06256_));
 sky130_fd_sc_hd__nand2_1 _26621_ (.A(_06255_),
    .B(_06256_),
    .Y(_01194_));
 sky130_fd_sc_hd__nand2_1 _26622_ (.A(_02653_),
    .B(_06233_),
    .Y(_06257_));
 sky130_fd_sc_hd__nand2_1 _26623_ (.A(\gen_regfile_ff.register_file_i.rf_reg[745] ),
    .B(_06237_),
    .Y(_06258_));
 sky130_fd_sc_hd__nand2_1 _26624_ (.A(_06257_),
    .B(_06258_),
    .Y(_01195_));
 sky130_fd_sc_hd__nand2_1 _26625_ (.A(_02761_),
    .B(_06233_),
    .Y(_06259_));
 sky130_fd_sc_hd__nand2_1 _26626_ (.A(\gen_regfile_ff.register_file_i.rf_reg[746] ),
    .B(_06237_),
    .Y(_06260_));
 sky130_fd_sc_hd__nand2_1 _26627_ (.A(_06259_),
    .B(_06260_),
    .Y(_01196_));
 sky130_fd_sc_hd__nand2_1 _26628_ (.A(_02849_),
    .B(_06233_),
    .Y(_06261_));
 sky130_fd_sc_hd__nand2_1 _26629_ (.A(\gen_regfile_ff.register_file_i.rf_reg[747] ),
    .B(_06237_),
    .Y(_06262_));
 sky130_fd_sc_hd__nand2_1 _26630_ (.A(_06261_),
    .B(_06262_),
    .Y(_01197_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_70 ();
 sky130_fd_sc_hd__nand2_1 _26632_ (.A(_02974_),
    .B(_06233_),
    .Y(_06264_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_69 ();
 sky130_fd_sc_hd__nand2_1 _26634_ (.A(\gen_regfile_ff.register_file_i.rf_reg[748] ),
    .B(_06237_),
    .Y(_06266_));
 sky130_fd_sc_hd__nand2_1 _26635_ (.A(_06264_),
    .B(_06266_),
    .Y(_01198_));
 sky130_fd_sc_hd__nand2_1 _26636_ (.A(_03080_),
    .B(_06233_),
    .Y(_06267_));
 sky130_fd_sc_hd__nand2_1 _26637_ (.A(\gen_regfile_ff.register_file_i.rf_reg[749] ),
    .B(_06237_),
    .Y(_06268_));
 sky130_fd_sc_hd__nand2_1 _26638_ (.A(_06267_),
    .B(_06268_),
    .Y(_01199_));
 sky130_fd_sc_hd__nand2_1 _26639_ (.A(_03214_),
    .B(_06233_),
    .Y(_06269_));
 sky130_fd_sc_hd__nand2_1 _26640_ (.A(\gen_regfile_ff.register_file_i.rf_reg[750] ),
    .B(_06237_),
    .Y(_06270_));
 sky130_fd_sc_hd__nand2_1 _26641_ (.A(_06269_),
    .B(_06270_),
    .Y(_01200_));
 sky130_fd_sc_hd__nand2_1 _26642_ (.A(_03348_),
    .B(_06233_),
    .Y(_06271_));
 sky130_fd_sc_hd__nand2_1 _26643_ (.A(\gen_regfile_ff.register_file_i.rf_reg[751] ),
    .B(_06237_),
    .Y(_06272_));
 sky130_fd_sc_hd__nand2_1 _26644_ (.A(_06271_),
    .B(_06272_),
    .Y(_01201_));
 sky130_fd_sc_hd__nand2_1 _26645_ (.A(_02468_),
    .B(_06112_),
    .Y(_06273_));
 sky130_fd_sc_hd__nand2_1 _26646_ (.A(\gen_regfile_ff.register_file_i.rf_reg[103] ),
    .B(_06115_),
    .Y(_06274_));
 sky130_fd_sc_hd__nand2_1 _26647_ (.A(_06273_),
    .B(_06274_),
    .Y(_01202_));
 sky130_fd_sc_hd__nand2_1 _26648_ (.A(\gen_regfile_ff.register_file_i.rf_reg[752] ),
    .B(_06237_),
    .Y(_06275_));
 sky130_fd_sc_hd__o21ai_0 _26649_ (.A1(_03481_),
    .A2(_06237_),
    .B1(_06275_),
    .Y(_01203_));
 sky130_fd_sc_hd__nand2_1 _26650_ (.A(net1575),
    .B(_06233_),
    .Y(_06276_));
 sky130_fd_sc_hd__nand2_1 _26651_ (.A(\gen_regfile_ff.register_file_i.rf_reg[753] ),
    .B(_06237_),
    .Y(_06277_));
 sky130_fd_sc_hd__nand2_1 _26652_ (.A(_06276_),
    .B(_06277_),
    .Y(_01204_));
 sky130_fd_sc_hd__nand2_1 _26653_ (.A(net1576),
    .B(_06233_),
    .Y(_06278_));
 sky130_fd_sc_hd__nand2_1 _26654_ (.A(\gen_regfile_ff.register_file_i.rf_reg[754] ),
    .B(_06237_),
    .Y(_06279_));
 sky130_fd_sc_hd__nand2_1 _26655_ (.A(_06278_),
    .B(_06279_),
    .Y(_01205_));
 sky130_fd_sc_hd__nand2_1 _26656_ (.A(net1551),
    .B(_06233_),
    .Y(_06280_));
 sky130_fd_sc_hd__nand2_1 _26657_ (.A(\gen_regfile_ff.register_file_i.rf_reg[755] ),
    .B(_06237_),
    .Y(_06281_));
 sky130_fd_sc_hd__nand2_1 _26658_ (.A(_06280_),
    .B(_06281_),
    .Y(_01206_));
 sky130_fd_sc_hd__nand2_1 _26659_ (.A(_03982_),
    .B(_06233_),
    .Y(_06282_));
 sky130_fd_sc_hd__nand2_1 _26660_ (.A(\gen_regfile_ff.register_file_i.rf_reg[756] ),
    .B(_06237_),
    .Y(_06283_));
 sky130_fd_sc_hd__nand2_1 _26661_ (.A(_06282_),
    .B(_06283_),
    .Y(_01207_));
 sky130_fd_sc_hd__nand2_1 _26662_ (.A(net1584),
    .B(_06233_),
    .Y(_06284_));
 sky130_fd_sc_hd__nand2_1 _26663_ (.A(\gen_regfile_ff.register_file_i.rf_reg[757] ),
    .B(_06237_),
    .Y(_06285_));
 sky130_fd_sc_hd__nand2_1 _26664_ (.A(_06284_),
    .B(_06285_),
    .Y(_01208_));
 sky130_fd_sc_hd__mux2_4 _26665_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[758] ),
    .A1(net1326),
    .S(_06233_),
    .X(_01209_));
 sky130_fd_sc_hd__nand2_2 _26666_ (.A(net1291),
    .B(_06233_),
    .Y(_06286_));
 sky130_fd_sc_hd__nand2_1 _26667_ (.A(\gen_regfile_ff.register_file_i.rf_reg[759] ),
    .B(_06237_),
    .Y(_06287_));
 sky130_fd_sc_hd__nand2_1 _26668_ (.A(_06286_),
    .B(_06287_),
    .Y(_01210_));
 sky130_fd_sc_hd__nand2_1 _26669_ (.A(net1541),
    .B(_06233_),
    .Y(_06288_));
 sky130_fd_sc_hd__nand2_1 _26670_ (.A(\gen_regfile_ff.register_file_i.rf_reg[760] ),
    .B(_06237_),
    .Y(_06289_));
 sky130_fd_sc_hd__nand2_1 _26671_ (.A(_06288_),
    .B(_06289_),
    .Y(_01211_));
 sky130_fd_sc_hd__nand2_1 _26672_ (.A(net1586),
    .B(_06233_),
    .Y(_06290_));
 sky130_fd_sc_hd__nand2_1 _26673_ (.A(\gen_regfile_ff.register_file_i.rf_reg[761] ),
    .B(_06237_),
    .Y(_06291_));
 sky130_fd_sc_hd__nand2_1 _26674_ (.A(_06290_),
    .B(_06291_),
    .Y(_01212_));
 sky130_fd_sc_hd__nand2_1 _26675_ (.A(_02553_),
    .B(_06112_),
    .Y(_06292_));
 sky130_fd_sc_hd__nand2_1 _26676_ (.A(\gen_regfile_ff.register_file_i.rf_reg[104] ),
    .B(_06115_),
    .Y(_06293_));
 sky130_fd_sc_hd__nand2_1 _26677_ (.A(_06292_),
    .B(_06293_),
    .Y(_01213_));
 sky130_fd_sc_hd__nand2_2 _26678_ (.A(net1536),
    .B(_06233_),
    .Y(_06294_));
 sky130_fd_sc_hd__nand2_1 _26679_ (.A(\gen_regfile_ff.register_file_i.rf_reg[762] ),
    .B(_06237_),
    .Y(_06295_));
 sky130_fd_sc_hd__nand2_1 _26680_ (.A(_06295_),
    .B(_06294_),
    .Y(_01214_));
 sky130_fd_sc_hd__nand2_2 _26681_ (.A(net1542),
    .B(_06233_),
    .Y(_06296_));
 sky130_fd_sc_hd__nand2_1 _26682_ (.A(\gen_regfile_ff.register_file_i.rf_reg[763] ),
    .B(_06237_),
    .Y(_06297_));
 sky130_fd_sc_hd__nand2_1 _26683_ (.A(_06296_),
    .B(_06297_),
    .Y(_01215_));
 sky130_fd_sc_hd__mux2_4 _26684_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[764] ),
    .A1(net1294),
    .S(_06233_),
    .X(_01216_));
 sky130_fd_sc_hd__nor2_1 _26685_ (.A(_05084_),
    .B(_06237_),
    .Y(_06298_));
 sky130_fd_sc_hd__a22o_1 _26686_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[765] ),
    .A2(_06237_),
    .B1(net1249),
    .B2(_06298_),
    .X(_01217_));
 sky130_fd_sc_hd__mux2_4 _26687_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[766] ),
    .A1(net1238),
    .S(_06233_),
    .X(_01218_));
 sky130_fd_sc_hd__nor2_1 _26688_ (.A(_05264_),
    .B(_06237_),
    .Y(_06299_));
 sky130_fd_sc_hd__a22o_1 _26689_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[767] ),
    .A2(_06237_),
    .B1(_06299_),
    .B2(net652),
    .X(_01219_));
 sky130_fd_sc_hd__nor2_8 _26690_ (.A(_05572_),
    .B(_06025_),
    .Y(_06300_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_68 ();
 sky130_fd_sc_hd__nand2_1 _26692_ (.A(_01909_),
    .B(_06300_),
    .Y(_06302_));
 sky130_fd_sc_hd__nand3_4 _26693_ (.A(net446),
    .B(_05955_),
    .C(net1253),
    .Y(_06303_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_67 ();
 sky130_fd_sc_hd__nand2_1 _26695_ (.A(\gen_regfile_ff.register_file_i.rf_reg[768] ),
    .B(_06303_),
    .Y(_06305_));
 sky130_fd_sc_hd__nand2_1 _26696_ (.A(_06302_),
    .B(_06305_),
    .Y(_01220_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_66 ();
 sky130_fd_sc_hd__nand2_1 _26698_ (.A(\gen_regfile_ff.register_file_i.rf_reg[769] ),
    .B(_06303_),
    .Y(_06307_));
 sky130_fd_sc_hd__o21ai_0 _26699_ (.A1(_05299_),
    .A2(_06303_),
    .B1(_06307_),
    .Y(_01221_));
 sky130_fd_sc_hd__nand2_1 _26700_ (.A(_05326_),
    .B(_06300_),
    .Y(_06308_));
 sky130_fd_sc_hd__nand2_1 _26701_ (.A(\gen_regfile_ff.register_file_i.rf_reg[770] ),
    .B(_06303_),
    .Y(_06309_));
 sky130_fd_sc_hd__nand2_1 _26702_ (.A(_06308_),
    .B(_06309_),
    .Y(_01222_));
 sky130_fd_sc_hd__nand2_1 _26703_ (.A(\gen_regfile_ff.register_file_i.rf_reg[771] ),
    .B(_06303_),
    .Y(_06310_));
 sky130_fd_sc_hd__o21ai_0 _26704_ (.A1(_05351_),
    .A2(_06303_),
    .B1(_06310_),
    .Y(_01223_));
 sky130_fd_sc_hd__nand2_1 _26705_ (.A(_02653_),
    .B(_06112_),
    .Y(_06311_));
 sky130_fd_sc_hd__nand2_1 _26706_ (.A(\gen_regfile_ff.register_file_i.rf_reg[105] ),
    .B(_06115_),
    .Y(_06312_));
 sky130_fd_sc_hd__nand2_1 _26707_ (.A(_06311_),
    .B(_06312_),
    .Y(_01224_));
 sky130_fd_sc_hd__nand2_1 _26708_ (.A(_02113_),
    .B(_06300_),
    .Y(_06313_));
 sky130_fd_sc_hd__nand2_1 _26709_ (.A(\gen_regfile_ff.register_file_i.rf_reg[772] ),
    .B(_06303_),
    .Y(_06314_));
 sky130_fd_sc_hd__nand2_1 _26710_ (.A(_06313_),
    .B(_06314_),
    .Y(_01225_));
 sky130_fd_sc_hd__nand2_1 _26711_ (.A(_02250_),
    .B(_06300_),
    .Y(_06315_));
 sky130_fd_sc_hd__nand2_1 _26712_ (.A(\gen_regfile_ff.register_file_i.rf_reg[773] ),
    .B(_06303_),
    .Y(_06316_));
 sky130_fd_sc_hd__nand2_1 _26713_ (.A(_06315_),
    .B(_06316_),
    .Y(_01226_));
 sky130_fd_sc_hd__nand2_1 _26714_ (.A(_02360_),
    .B(_06300_),
    .Y(_06317_));
 sky130_fd_sc_hd__nand2_1 _26715_ (.A(\gen_regfile_ff.register_file_i.rf_reg[774] ),
    .B(_06303_),
    .Y(_06318_));
 sky130_fd_sc_hd__nand2_1 _26716_ (.A(_06317_),
    .B(_06318_),
    .Y(_01227_));
 sky130_fd_sc_hd__nand2_1 _26717_ (.A(_02468_),
    .B(_06300_),
    .Y(_06319_));
 sky130_fd_sc_hd__nand2_1 _26718_ (.A(\gen_regfile_ff.register_file_i.rf_reg[775] ),
    .B(_06303_),
    .Y(_06320_));
 sky130_fd_sc_hd__nand2_1 _26719_ (.A(_06319_),
    .B(_06320_),
    .Y(_01228_));
 sky130_fd_sc_hd__nand2_1 _26720_ (.A(_02553_),
    .B(_06300_),
    .Y(_06321_));
 sky130_fd_sc_hd__nand2_1 _26721_ (.A(\gen_regfile_ff.register_file_i.rf_reg[776] ),
    .B(_06303_),
    .Y(_06322_));
 sky130_fd_sc_hd__nand2_1 _26722_ (.A(_06321_),
    .B(_06322_),
    .Y(_01229_));
 sky130_fd_sc_hd__nand2_1 _26723_ (.A(_02653_),
    .B(_06300_),
    .Y(_06323_));
 sky130_fd_sc_hd__nand2_1 _26724_ (.A(\gen_regfile_ff.register_file_i.rf_reg[777] ),
    .B(_06303_),
    .Y(_06324_));
 sky130_fd_sc_hd__nand2_1 _26725_ (.A(_06323_),
    .B(_06324_),
    .Y(_01230_));
 sky130_fd_sc_hd__nand2_1 _26726_ (.A(_02761_),
    .B(_06300_),
    .Y(_06325_));
 sky130_fd_sc_hd__nand2_1 _26727_ (.A(\gen_regfile_ff.register_file_i.rf_reg[778] ),
    .B(_06303_),
    .Y(_06326_));
 sky130_fd_sc_hd__nand2_1 _26728_ (.A(_06325_),
    .B(_06326_),
    .Y(_01231_));
 sky130_fd_sc_hd__nand2_1 _26729_ (.A(_02849_),
    .B(_06300_),
    .Y(_06327_));
 sky130_fd_sc_hd__nand2_1 _26730_ (.A(\gen_regfile_ff.register_file_i.rf_reg[779] ),
    .B(_06303_),
    .Y(_06328_));
 sky130_fd_sc_hd__nand2_1 _26731_ (.A(_06327_),
    .B(_06328_),
    .Y(_01232_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_65 ();
 sky130_fd_sc_hd__nand2_1 _26733_ (.A(_02974_),
    .B(_06300_),
    .Y(_06330_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_64 ();
 sky130_fd_sc_hd__nand2_1 _26735_ (.A(\gen_regfile_ff.register_file_i.rf_reg[780] ),
    .B(_06303_),
    .Y(_06332_));
 sky130_fd_sc_hd__nand2_1 _26736_ (.A(_06330_),
    .B(_06332_),
    .Y(_01233_));
 sky130_fd_sc_hd__nand2_1 _26737_ (.A(_03080_),
    .B(_06300_),
    .Y(_06333_));
 sky130_fd_sc_hd__nand2_1 _26738_ (.A(\gen_regfile_ff.register_file_i.rf_reg[781] ),
    .B(_06303_),
    .Y(_06334_));
 sky130_fd_sc_hd__nand2_1 _26739_ (.A(_06333_),
    .B(_06334_),
    .Y(_01234_));
 sky130_fd_sc_hd__nand2_1 _26740_ (.A(_02761_),
    .B(_06112_),
    .Y(_06335_));
 sky130_fd_sc_hd__nand2_1 _26741_ (.A(\gen_regfile_ff.register_file_i.rf_reg[106] ),
    .B(_06115_),
    .Y(_06336_));
 sky130_fd_sc_hd__nand2_1 _26742_ (.A(_06335_),
    .B(_06336_),
    .Y(_01235_));
 sky130_fd_sc_hd__nand2_1 _26743_ (.A(_03214_),
    .B(_06300_),
    .Y(_06337_));
 sky130_fd_sc_hd__nand2_1 _26744_ (.A(\gen_regfile_ff.register_file_i.rf_reg[782] ),
    .B(_06303_),
    .Y(_06338_));
 sky130_fd_sc_hd__nand2_1 _26745_ (.A(_06337_),
    .B(_06338_),
    .Y(_01236_));
 sky130_fd_sc_hd__nand2_1 _26746_ (.A(_03348_),
    .B(_06300_),
    .Y(_06339_));
 sky130_fd_sc_hd__nand2_1 _26747_ (.A(\gen_regfile_ff.register_file_i.rf_reg[783] ),
    .B(_06303_),
    .Y(_06340_));
 sky130_fd_sc_hd__nand2_1 _26748_ (.A(_06339_),
    .B(_06340_),
    .Y(_01237_));
 sky130_fd_sc_hd__nand2_1 _26749_ (.A(\gen_regfile_ff.register_file_i.rf_reg[784] ),
    .B(_06303_),
    .Y(_06341_));
 sky130_fd_sc_hd__o21ai_0 _26750_ (.A1(_03481_),
    .A2(_06303_),
    .B1(_06341_),
    .Y(_01238_));
 sky130_fd_sc_hd__nand2_1 _26751_ (.A(net1575),
    .B(_06300_),
    .Y(_06342_));
 sky130_fd_sc_hd__nand2_1 _26752_ (.A(\gen_regfile_ff.register_file_i.rf_reg[785] ),
    .B(_06303_),
    .Y(_06343_));
 sky130_fd_sc_hd__nand2_1 _26753_ (.A(_06342_),
    .B(_06343_),
    .Y(_01239_));
 sky130_fd_sc_hd__nand2_1 _26754_ (.A(_03739_),
    .B(_06300_),
    .Y(_06344_));
 sky130_fd_sc_hd__nand2_1 _26755_ (.A(\gen_regfile_ff.register_file_i.rf_reg[786] ),
    .B(_06303_),
    .Y(_06345_));
 sky130_fd_sc_hd__nand2_1 _26756_ (.A(_06344_),
    .B(_06345_),
    .Y(_01240_));
 sky130_fd_sc_hd__nand2_1 _26757_ (.A(net1551),
    .B(_06300_),
    .Y(_06346_));
 sky130_fd_sc_hd__nand2_1 _26758_ (.A(\gen_regfile_ff.register_file_i.rf_reg[787] ),
    .B(_06303_),
    .Y(_06347_));
 sky130_fd_sc_hd__nand2_1 _26759_ (.A(_06346_),
    .B(_06347_),
    .Y(_01241_));
 sky130_fd_sc_hd__nand2_1 _26760_ (.A(_03982_),
    .B(_06300_),
    .Y(_06348_));
 sky130_fd_sc_hd__nand2_1 _26761_ (.A(\gen_regfile_ff.register_file_i.rf_reg[788] ),
    .B(_06303_),
    .Y(_06349_));
 sky130_fd_sc_hd__nand2_1 _26762_ (.A(_06348_),
    .B(_06349_),
    .Y(_01242_));
 sky130_fd_sc_hd__nand2_1 _26763_ (.A(net1584),
    .B(_06300_),
    .Y(_06350_));
 sky130_fd_sc_hd__nand2_1 _26764_ (.A(\gen_regfile_ff.register_file_i.rf_reg[789] ),
    .B(_06303_),
    .Y(_06351_));
 sky130_fd_sc_hd__nand2_1 _26765_ (.A(_06350_),
    .B(_06351_),
    .Y(_01243_));
 sky130_fd_sc_hd__mux2_4 _26766_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[790] ),
    .A1(net1326),
    .S(_06300_),
    .X(_01244_));
 sky130_fd_sc_hd__nand2_2 _26767_ (.A(net1290),
    .B(_06300_),
    .Y(_06352_));
 sky130_fd_sc_hd__nand2_1 _26768_ (.A(\gen_regfile_ff.register_file_i.rf_reg[791] ),
    .B(_06303_),
    .Y(_06353_));
 sky130_fd_sc_hd__nand2_1 _26769_ (.A(_06352_),
    .B(_06353_),
    .Y(_01245_));
 sky130_fd_sc_hd__nand2_1 _26770_ (.A(_02849_),
    .B(_06112_),
    .Y(_06354_));
 sky130_fd_sc_hd__nand2_1 _26771_ (.A(\gen_regfile_ff.register_file_i.rf_reg[107] ),
    .B(_06115_),
    .Y(_06355_));
 sky130_fd_sc_hd__nand2_1 _26772_ (.A(_06354_),
    .B(_06355_),
    .Y(_01246_));
 sky130_fd_sc_hd__nand2_2 _26773_ (.A(net1271),
    .B(_06300_),
    .Y(_06356_));
 sky130_fd_sc_hd__nand2_1 _26774_ (.A(\gen_regfile_ff.register_file_i.rf_reg[792] ),
    .B(_06303_),
    .Y(_06357_));
 sky130_fd_sc_hd__nand2_1 _26775_ (.A(_06356_),
    .B(_06357_),
    .Y(_01247_));
 sky130_fd_sc_hd__nand2_1 _26776_ (.A(net252),
    .B(_06300_),
    .Y(_06358_));
 sky130_fd_sc_hd__nand2_1 _26777_ (.A(\gen_regfile_ff.register_file_i.rf_reg[793] ),
    .B(_06303_),
    .Y(_06359_));
 sky130_fd_sc_hd__nand2_1 _26778_ (.A(_06358_),
    .B(_06359_),
    .Y(_01248_));
 sky130_fd_sc_hd__nand2_4 _26779_ (.A(net1514),
    .B(_06300_),
    .Y(_06360_));
 sky130_fd_sc_hd__nand2_1 _26780_ (.A(\gen_regfile_ff.register_file_i.rf_reg[794] ),
    .B(_06303_),
    .Y(_06361_));
 sky130_fd_sc_hd__nand2_1 _26781_ (.A(_06360_),
    .B(_06361_),
    .Y(_01249_));
 sky130_fd_sc_hd__nand2_1 _26782_ (.A(net1539),
    .B(_06300_),
    .Y(_06362_));
 sky130_fd_sc_hd__nand2_1 _26783_ (.A(\gen_regfile_ff.register_file_i.rf_reg[795] ),
    .B(_06303_),
    .Y(_06363_));
 sky130_fd_sc_hd__nand2_1 _26784_ (.A(_06362_),
    .B(_06363_),
    .Y(_01250_));
 sky130_fd_sc_hd__mux2_4 _26785_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[796] ),
    .A1(net885),
    .S(_06300_),
    .X(_01251_));
 sky130_fd_sc_hd__nor2_1 _26786_ (.A(_05084_),
    .B(_06303_),
    .Y(_06364_));
 sky130_fd_sc_hd__a22o_1 _26787_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[797] ),
    .A2(_06303_),
    .B1(net1254),
    .B2(_06364_),
    .X(_01252_));
 sky130_fd_sc_hd__mux2_4 _26788_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[798] ),
    .A1(net1238),
    .S(_06300_),
    .X(_01253_));
 sky130_fd_sc_hd__nor2_1 _26789_ (.A(_05264_),
    .B(_06303_),
    .Y(_06365_));
 sky130_fd_sc_hd__a22o_1 _26790_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[799] ),
    .A2(_06303_),
    .B1(_06365_),
    .B2(net500),
    .X(_01254_));
 sky130_fd_sc_hd__nor2_8 _26791_ (.A(_05572_),
    .B(_06088_),
    .Y(_06366_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_63 ();
 sky130_fd_sc_hd__nand2_1 _26793_ (.A(_01909_),
    .B(_06366_),
    .Y(_06368_));
 sky130_fd_sc_hd__nand3_4 _26794_ (.A(net446),
    .B(_01919_),
    .C(net1253),
    .Y(_06369_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_62 ();
 sky130_fd_sc_hd__nand2_1 _26796_ (.A(\gen_regfile_ff.register_file_i.rf_reg[800] ),
    .B(_06369_),
    .Y(_06371_));
 sky130_fd_sc_hd__nand2_1 _26797_ (.A(_06368_),
    .B(_06371_),
    .Y(_01255_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_61 ();
 sky130_fd_sc_hd__nand2_1 _26799_ (.A(\gen_regfile_ff.register_file_i.rf_reg[801] ),
    .B(_06369_),
    .Y(_06373_));
 sky130_fd_sc_hd__o21ai_0 _26800_ (.A1(_05299_),
    .A2(_06369_),
    .B1(_06373_),
    .Y(_01256_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_60 ();
 sky130_fd_sc_hd__nand2_1 _26802_ (.A(_02974_),
    .B(_06112_),
    .Y(_06375_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_59 ();
 sky130_fd_sc_hd__nand2_1 _26804_ (.A(\gen_regfile_ff.register_file_i.rf_reg[108] ),
    .B(_06115_),
    .Y(_06377_));
 sky130_fd_sc_hd__nand2_1 _26805_ (.A(_06375_),
    .B(_06377_),
    .Y(_01257_));
 sky130_fd_sc_hd__nand2_1 _26806_ (.A(_05326_),
    .B(_06366_),
    .Y(_06378_));
 sky130_fd_sc_hd__nand2_1 _26807_ (.A(\gen_regfile_ff.register_file_i.rf_reg[802] ),
    .B(_06369_),
    .Y(_06379_));
 sky130_fd_sc_hd__nand2_1 _26808_ (.A(_06378_),
    .B(_06379_),
    .Y(_01258_));
 sky130_fd_sc_hd__nand2_1 _26809_ (.A(\gen_regfile_ff.register_file_i.rf_reg[803] ),
    .B(_06369_),
    .Y(_06380_));
 sky130_fd_sc_hd__o21ai_0 _26810_ (.A1(_05351_),
    .A2(_06369_),
    .B1(_06380_),
    .Y(_01259_));
 sky130_fd_sc_hd__nand2_1 _26811_ (.A(_02113_),
    .B(_06366_),
    .Y(_06381_));
 sky130_fd_sc_hd__nand2_1 _26812_ (.A(\gen_regfile_ff.register_file_i.rf_reg[804] ),
    .B(_06369_),
    .Y(_06382_));
 sky130_fd_sc_hd__nand2_1 _26813_ (.A(_06381_),
    .B(_06382_),
    .Y(_01260_));
 sky130_fd_sc_hd__nand2_1 _26814_ (.A(_02250_),
    .B(_06366_),
    .Y(_06383_));
 sky130_fd_sc_hd__nand2_1 _26815_ (.A(\gen_regfile_ff.register_file_i.rf_reg[805] ),
    .B(_06369_),
    .Y(_06384_));
 sky130_fd_sc_hd__nand2_1 _26816_ (.A(_06383_),
    .B(_06384_),
    .Y(_01261_));
 sky130_fd_sc_hd__nand2_1 _26817_ (.A(_02360_),
    .B(_06366_),
    .Y(_06385_));
 sky130_fd_sc_hd__nand2_1 _26818_ (.A(\gen_regfile_ff.register_file_i.rf_reg[806] ),
    .B(_06369_),
    .Y(_06386_));
 sky130_fd_sc_hd__nand2_1 _26819_ (.A(_06385_),
    .B(_06386_),
    .Y(_01262_));
 sky130_fd_sc_hd__nand2_1 _26820_ (.A(_02468_),
    .B(_06366_),
    .Y(_06387_));
 sky130_fd_sc_hd__nand2_1 _26821_ (.A(\gen_regfile_ff.register_file_i.rf_reg[807] ),
    .B(_06369_),
    .Y(_06388_));
 sky130_fd_sc_hd__nand2_1 _26822_ (.A(_06387_),
    .B(_06388_),
    .Y(_01263_));
 sky130_fd_sc_hd__nand2_1 _26823_ (.A(_02553_),
    .B(_06366_),
    .Y(_06389_));
 sky130_fd_sc_hd__nand2_1 _26824_ (.A(\gen_regfile_ff.register_file_i.rf_reg[808] ),
    .B(_06369_),
    .Y(_06390_));
 sky130_fd_sc_hd__nand2_1 _26825_ (.A(_06389_),
    .B(_06390_),
    .Y(_01264_));
 sky130_fd_sc_hd__nand2_1 _26826_ (.A(_02653_),
    .B(_06366_),
    .Y(_06391_));
 sky130_fd_sc_hd__nand2_1 _26827_ (.A(\gen_regfile_ff.register_file_i.rf_reg[809] ),
    .B(_06369_),
    .Y(_06392_));
 sky130_fd_sc_hd__nand2_1 _26828_ (.A(_06391_),
    .B(_06392_),
    .Y(_01265_));
 sky130_fd_sc_hd__nand2_1 _26829_ (.A(_02761_),
    .B(_06366_),
    .Y(_06393_));
 sky130_fd_sc_hd__nand2_1 _26830_ (.A(\gen_regfile_ff.register_file_i.rf_reg[810] ),
    .B(_06369_),
    .Y(_06394_));
 sky130_fd_sc_hd__nand2_1 _26831_ (.A(_06393_),
    .B(_06394_),
    .Y(_01266_));
 sky130_fd_sc_hd__nand2_1 _26832_ (.A(_02849_),
    .B(_06366_),
    .Y(_06395_));
 sky130_fd_sc_hd__nand2_1 _26833_ (.A(\gen_regfile_ff.register_file_i.rf_reg[811] ),
    .B(_06369_),
    .Y(_06396_));
 sky130_fd_sc_hd__nand2_1 _26834_ (.A(_06395_),
    .B(_06396_),
    .Y(_01267_));
 sky130_fd_sc_hd__nand2_1 _26835_ (.A(_03080_),
    .B(_06112_),
    .Y(_06397_));
 sky130_fd_sc_hd__nand2_1 _26836_ (.A(\gen_regfile_ff.register_file_i.rf_reg[109] ),
    .B(_06115_),
    .Y(_06398_));
 sky130_fd_sc_hd__nand2_1 _26837_ (.A(_06397_),
    .B(_06398_),
    .Y(_01268_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_58 ();
 sky130_fd_sc_hd__nand2_1 _26839_ (.A(_02974_),
    .B(_06366_),
    .Y(_06400_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_57 ();
 sky130_fd_sc_hd__nand2_1 _26841_ (.A(\gen_regfile_ff.register_file_i.rf_reg[812] ),
    .B(_06369_),
    .Y(_06402_));
 sky130_fd_sc_hd__nand2_1 _26842_ (.A(_06400_),
    .B(_06402_),
    .Y(_01269_));
 sky130_fd_sc_hd__nand2_1 _26843_ (.A(_03080_),
    .B(_06366_),
    .Y(_06403_));
 sky130_fd_sc_hd__nand2_1 _26844_ (.A(\gen_regfile_ff.register_file_i.rf_reg[813] ),
    .B(_06369_),
    .Y(_06404_));
 sky130_fd_sc_hd__nand2_1 _26845_ (.A(_06403_),
    .B(_06404_),
    .Y(_01270_));
 sky130_fd_sc_hd__nand2_1 _26846_ (.A(_03214_),
    .B(_06366_),
    .Y(_06405_));
 sky130_fd_sc_hd__nand2_1 _26847_ (.A(\gen_regfile_ff.register_file_i.rf_reg[814] ),
    .B(_06369_),
    .Y(_06406_));
 sky130_fd_sc_hd__nand2_1 _26848_ (.A(_06405_),
    .B(_06406_),
    .Y(_01271_));
 sky130_fd_sc_hd__nand2_1 _26849_ (.A(_03348_),
    .B(_06366_),
    .Y(_06407_));
 sky130_fd_sc_hd__nand2_1 _26850_ (.A(\gen_regfile_ff.register_file_i.rf_reg[815] ),
    .B(_06369_),
    .Y(_06408_));
 sky130_fd_sc_hd__nand2_1 _26851_ (.A(_06407_),
    .B(_06408_),
    .Y(_01272_));
 sky130_fd_sc_hd__nand2_1 _26852_ (.A(\gen_regfile_ff.register_file_i.rf_reg[816] ),
    .B(_06369_),
    .Y(_06409_));
 sky130_fd_sc_hd__o21ai_0 _26853_ (.A1(_03481_),
    .A2(_06369_),
    .B1(_06409_),
    .Y(_01273_));
 sky130_fd_sc_hd__nand2_1 _26854_ (.A(net1575),
    .B(_06366_),
    .Y(_06410_));
 sky130_fd_sc_hd__nand2_1 _26855_ (.A(\gen_regfile_ff.register_file_i.rf_reg[817] ),
    .B(_06369_),
    .Y(_06411_));
 sky130_fd_sc_hd__nand2_1 _26856_ (.A(_06410_),
    .B(_06411_),
    .Y(_01274_));
 sky130_fd_sc_hd__nand2_1 _26857_ (.A(_03739_),
    .B(_06366_),
    .Y(_06412_));
 sky130_fd_sc_hd__nand2_1 _26858_ (.A(\gen_regfile_ff.register_file_i.rf_reg[818] ),
    .B(_06369_),
    .Y(_06413_));
 sky130_fd_sc_hd__nand2_1 _26859_ (.A(_06412_),
    .B(_06413_),
    .Y(_01275_));
 sky130_fd_sc_hd__nand2_1 _26860_ (.A(_03866_),
    .B(_06366_),
    .Y(_06414_));
 sky130_fd_sc_hd__nand2_1 _26861_ (.A(\gen_regfile_ff.register_file_i.rf_reg[819] ),
    .B(_06369_),
    .Y(_06415_));
 sky130_fd_sc_hd__nand2_1 _26862_ (.A(_06414_),
    .B(_06415_),
    .Y(_01276_));
 sky130_fd_sc_hd__nand2_1 _26863_ (.A(net1544),
    .B(_06366_),
    .Y(_06416_));
 sky130_fd_sc_hd__nand2_1 _26864_ (.A(\gen_regfile_ff.register_file_i.rf_reg[820] ),
    .B(_06369_),
    .Y(_06417_));
 sky130_fd_sc_hd__nand2_1 _26865_ (.A(_06416_),
    .B(_06417_),
    .Y(_01277_));
 sky130_fd_sc_hd__nand2_1 _26866_ (.A(net1584),
    .B(_06366_),
    .Y(_06418_));
 sky130_fd_sc_hd__nand2_1 _26867_ (.A(\gen_regfile_ff.register_file_i.rf_reg[821] ),
    .B(_06369_),
    .Y(_06419_));
 sky130_fd_sc_hd__nand2_1 _26868_ (.A(_06418_),
    .B(_06419_),
    .Y(_01278_));
 sky130_fd_sc_hd__nand2_1 _26869_ (.A(_03214_),
    .B(_06112_),
    .Y(_06420_));
 sky130_fd_sc_hd__nand2_1 _26870_ (.A(\gen_regfile_ff.register_file_i.rf_reg[110] ),
    .B(_06115_),
    .Y(_06421_));
 sky130_fd_sc_hd__nand2_1 _26871_ (.A(_06420_),
    .B(_06421_),
    .Y(_01279_));
 sky130_fd_sc_hd__mux2_4 _26872_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[822] ),
    .A1(net1517),
    .S(_06366_),
    .X(_01280_));
 sky130_fd_sc_hd__nand2_2 _26873_ (.A(net1290),
    .B(_06366_),
    .Y(_06422_));
 sky130_fd_sc_hd__nand2_1 _26874_ (.A(\gen_regfile_ff.register_file_i.rf_reg[823] ),
    .B(_06369_),
    .Y(_06423_));
 sky130_fd_sc_hd__nand2_2 _26875_ (.A(_06423_),
    .B(_06422_),
    .Y(_01281_));
 sky130_fd_sc_hd__nand2_2 _26876_ (.A(net1271),
    .B(_06366_),
    .Y(_06424_));
 sky130_fd_sc_hd__nand2_1 _26877_ (.A(\gen_regfile_ff.register_file_i.rf_reg[824] ),
    .B(_06369_),
    .Y(_06425_));
 sky130_fd_sc_hd__nand2_1 _26878_ (.A(_06424_),
    .B(_06425_),
    .Y(_01282_));
 sky130_fd_sc_hd__nand2_1 _26879_ (.A(net1564),
    .B(_06366_),
    .Y(_06426_));
 sky130_fd_sc_hd__nand2_1 _26880_ (.A(\gen_regfile_ff.register_file_i.rf_reg[825] ),
    .B(_06369_),
    .Y(_06427_));
 sky130_fd_sc_hd__nand2_1 _26881_ (.A(_06426_),
    .B(_06427_),
    .Y(_01283_));
 sky130_fd_sc_hd__nand2_4 _26882_ (.A(net1514),
    .B(_06366_),
    .Y(_06428_));
 sky130_fd_sc_hd__nand2_1 _26883_ (.A(\gen_regfile_ff.register_file_i.rf_reg[826] ),
    .B(_06369_),
    .Y(_06429_));
 sky130_fd_sc_hd__nand2_2 _26884_ (.A(_06428_),
    .B(_06429_),
    .Y(_01284_));
 sky130_fd_sc_hd__nand2_1 _26885_ (.A(net1542),
    .B(_06366_),
    .Y(_06430_));
 sky130_fd_sc_hd__nand2_1 _26886_ (.A(\gen_regfile_ff.register_file_i.rf_reg[827] ),
    .B(_06369_),
    .Y(_06431_));
 sky130_fd_sc_hd__nand2_1 _26887_ (.A(_06430_),
    .B(_06431_),
    .Y(_01285_));
 sky130_fd_sc_hd__mux2_4 _26888_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[828] ),
    .A1(net885),
    .S(_06366_),
    .X(_01286_));
 sky130_fd_sc_hd__nor2_1 _26889_ (.A(_05084_),
    .B(_06369_),
    .Y(_06432_));
 sky130_fd_sc_hd__a22o_1 _26890_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[829] ),
    .A2(_06369_),
    .B1(_05079_),
    .B2(_06432_),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_4 _26891_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[830] ),
    .A1(net685),
    .S(_06366_),
    .X(_01288_));
 sky130_fd_sc_hd__nor2_1 _26892_ (.A(_05264_),
    .B(_06369_),
    .Y(_06433_));
 sky130_fd_sc_hd__a22o_1 _26893_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[831] ),
    .A2(_06369_),
    .B1(_06433_),
    .B2(net740),
    .X(_01289_));
 sky130_fd_sc_hd__nand2_1 _26894_ (.A(_03348_),
    .B(_06112_),
    .Y(_06434_));
 sky130_fd_sc_hd__nand2_1 _26895_ (.A(\gen_regfile_ff.register_file_i.rf_reg[111] ),
    .B(_06115_),
    .Y(_06435_));
 sky130_fd_sc_hd__nand2_1 _26896_ (.A(_06434_),
    .B(_06435_),
    .Y(_01290_));
 sky130_fd_sc_hd__nand2_1 _26897_ (.A(_01916_),
    .B(_02468_),
    .Y(_06436_));
 sky130_fd_sc_hd__nand2_1 _26898_ (.A(\gen_regfile_ff.register_file_i.rf_reg[39] ),
    .B(_01921_),
    .Y(_06437_));
 sky130_fd_sc_hd__nand2_1 _26899_ (.A(_06436_),
    .B(_06437_),
    .Y(_01291_));
 sky130_fd_sc_hd__nor2_8 _26900_ (.A(_05572_),
    .B(_06160_),
    .Y(_06438_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_56 ();
 sky130_fd_sc_hd__nand2_1 _26902_ (.A(_01909_),
    .B(_06438_),
    .Y(_06440_));
 sky130_fd_sc_hd__nand3_4 _26903_ (.A(net446),
    .B(_05796_),
    .C(net1253),
    .Y(_06441_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_55 ();
 sky130_fd_sc_hd__nand2_1 _26905_ (.A(\gen_regfile_ff.register_file_i.rf_reg[832] ),
    .B(_06441_),
    .Y(_06443_));
 sky130_fd_sc_hd__nand2_1 _26906_ (.A(_06440_),
    .B(_06443_),
    .Y(_01292_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_54 ();
 sky130_fd_sc_hd__nand2_1 _26908_ (.A(\gen_regfile_ff.register_file_i.rf_reg[833] ),
    .B(_06441_),
    .Y(_06445_));
 sky130_fd_sc_hd__o21ai_0 _26909_ (.A1(_05299_),
    .A2(_06441_),
    .B1(_06445_),
    .Y(_01293_));
 sky130_fd_sc_hd__nand2_1 _26910_ (.A(_05326_),
    .B(_06438_),
    .Y(_06446_));
 sky130_fd_sc_hd__nand2_1 _26911_ (.A(\gen_regfile_ff.register_file_i.rf_reg[834] ),
    .B(_06441_),
    .Y(_06447_));
 sky130_fd_sc_hd__nand2_1 _26912_ (.A(_06446_),
    .B(_06447_),
    .Y(_01294_));
 sky130_fd_sc_hd__nand2_1 _26913_ (.A(\gen_regfile_ff.register_file_i.rf_reg[835] ),
    .B(_06441_),
    .Y(_06448_));
 sky130_fd_sc_hd__o21ai_0 _26914_ (.A1(_05351_),
    .A2(_06441_),
    .B1(_06448_),
    .Y(_01295_));
 sky130_fd_sc_hd__nand2_1 _26915_ (.A(_02113_),
    .B(_06438_),
    .Y(_06449_));
 sky130_fd_sc_hd__nand2_1 _26916_ (.A(\gen_regfile_ff.register_file_i.rf_reg[836] ),
    .B(_06441_),
    .Y(_06450_));
 sky130_fd_sc_hd__nand2_1 _26917_ (.A(_06449_),
    .B(_06450_),
    .Y(_01296_));
 sky130_fd_sc_hd__nand2_1 _26918_ (.A(_02250_),
    .B(_06438_),
    .Y(_06451_));
 sky130_fd_sc_hd__nand2_1 _26919_ (.A(\gen_regfile_ff.register_file_i.rf_reg[837] ),
    .B(_06441_),
    .Y(_06452_));
 sky130_fd_sc_hd__nand2_1 _26920_ (.A(_06451_),
    .B(_06452_),
    .Y(_01297_));
 sky130_fd_sc_hd__nand2_1 _26921_ (.A(_02360_),
    .B(_06438_),
    .Y(_06453_));
 sky130_fd_sc_hd__nand2_1 _26922_ (.A(\gen_regfile_ff.register_file_i.rf_reg[838] ),
    .B(_06441_),
    .Y(_06454_));
 sky130_fd_sc_hd__nand2_1 _26923_ (.A(_06453_),
    .B(_06454_),
    .Y(_01298_));
 sky130_fd_sc_hd__nand2_1 _26924_ (.A(_02468_),
    .B(_06438_),
    .Y(_06455_));
 sky130_fd_sc_hd__nand2_1 _26925_ (.A(\gen_regfile_ff.register_file_i.rf_reg[839] ),
    .B(_06441_),
    .Y(_06456_));
 sky130_fd_sc_hd__nand2_1 _26926_ (.A(_06455_),
    .B(_06456_),
    .Y(_01299_));
 sky130_fd_sc_hd__nand2_1 _26927_ (.A(_02553_),
    .B(_06438_),
    .Y(_06457_));
 sky130_fd_sc_hd__nand2_1 _26928_ (.A(\gen_regfile_ff.register_file_i.rf_reg[840] ),
    .B(_06441_),
    .Y(_06458_));
 sky130_fd_sc_hd__nand2_1 _26929_ (.A(_06457_),
    .B(_06458_),
    .Y(_01300_));
 sky130_fd_sc_hd__nand2_1 _26930_ (.A(_02653_),
    .B(_06438_),
    .Y(_06459_));
 sky130_fd_sc_hd__nand2_1 _26931_ (.A(\gen_regfile_ff.register_file_i.rf_reg[841] ),
    .B(_06441_),
    .Y(_06460_));
 sky130_fd_sc_hd__nand2_1 _26932_ (.A(_06459_),
    .B(_06460_),
    .Y(_01301_));
 sky130_fd_sc_hd__nand2_1 _26933_ (.A(\gen_regfile_ff.register_file_i.rf_reg[112] ),
    .B(_06115_),
    .Y(_06461_));
 sky130_fd_sc_hd__o21ai_0 _26934_ (.A1(_03481_),
    .A2(_06115_),
    .B1(_06461_),
    .Y(_01302_));
 sky130_fd_sc_hd__nand2_1 _26935_ (.A(_02761_),
    .B(_06438_),
    .Y(_06462_));
 sky130_fd_sc_hd__nand2_1 _26936_ (.A(\gen_regfile_ff.register_file_i.rf_reg[842] ),
    .B(_06441_),
    .Y(_06463_));
 sky130_fd_sc_hd__nand2_1 _26937_ (.A(_06462_),
    .B(_06463_),
    .Y(_01303_));
 sky130_fd_sc_hd__nand2_1 _26938_ (.A(_02849_),
    .B(_06438_),
    .Y(_06464_));
 sky130_fd_sc_hd__nand2_1 _26939_ (.A(\gen_regfile_ff.register_file_i.rf_reg[843] ),
    .B(_06441_),
    .Y(_06465_));
 sky130_fd_sc_hd__nand2_1 _26940_ (.A(_06464_),
    .B(_06465_),
    .Y(_01304_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_53 ();
 sky130_fd_sc_hd__nand2_1 _26942_ (.A(_02974_),
    .B(_06438_),
    .Y(_06467_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_52 ();
 sky130_fd_sc_hd__nand2_1 _26944_ (.A(\gen_regfile_ff.register_file_i.rf_reg[844] ),
    .B(_06441_),
    .Y(_06469_));
 sky130_fd_sc_hd__nand2_1 _26945_ (.A(_06467_),
    .B(_06469_),
    .Y(_01305_));
 sky130_fd_sc_hd__nand2_1 _26946_ (.A(_03080_),
    .B(_06438_),
    .Y(_06470_));
 sky130_fd_sc_hd__nand2_1 _26947_ (.A(\gen_regfile_ff.register_file_i.rf_reg[845] ),
    .B(_06441_),
    .Y(_06471_));
 sky130_fd_sc_hd__nand2_1 _26948_ (.A(_06470_),
    .B(_06471_),
    .Y(_01306_));
 sky130_fd_sc_hd__nand2_1 _26949_ (.A(_03214_),
    .B(_06438_),
    .Y(_06472_));
 sky130_fd_sc_hd__nand2_1 _26950_ (.A(\gen_regfile_ff.register_file_i.rf_reg[846] ),
    .B(_06441_),
    .Y(_06473_));
 sky130_fd_sc_hd__nand2_1 _26951_ (.A(_06472_),
    .B(_06473_),
    .Y(_01307_));
 sky130_fd_sc_hd__nand2_1 _26952_ (.A(_03348_),
    .B(_06438_),
    .Y(_06474_));
 sky130_fd_sc_hd__nand2_1 _26953_ (.A(\gen_regfile_ff.register_file_i.rf_reg[847] ),
    .B(_06441_),
    .Y(_06475_));
 sky130_fd_sc_hd__nand2_1 _26954_ (.A(_06474_),
    .B(_06475_),
    .Y(_01308_));
 sky130_fd_sc_hd__nand2_1 _26955_ (.A(\gen_regfile_ff.register_file_i.rf_reg[848] ),
    .B(_06441_),
    .Y(_06476_));
 sky130_fd_sc_hd__o21ai_0 _26956_ (.A1(_03481_),
    .A2(_06441_),
    .B1(_06476_),
    .Y(_01309_));
 sky130_fd_sc_hd__nand2_1 _26957_ (.A(net1575),
    .B(_06438_),
    .Y(_06477_));
 sky130_fd_sc_hd__nand2_1 _26958_ (.A(\gen_regfile_ff.register_file_i.rf_reg[849] ),
    .B(_06441_),
    .Y(_06478_));
 sky130_fd_sc_hd__nand2_1 _26959_ (.A(_06477_),
    .B(_06478_),
    .Y(_01310_));
 sky130_fd_sc_hd__nand2_1 _26960_ (.A(net1576),
    .B(_06438_),
    .Y(_06479_));
 sky130_fd_sc_hd__nand2_1 _26961_ (.A(\gen_regfile_ff.register_file_i.rf_reg[850] ),
    .B(_06441_),
    .Y(_06480_));
 sky130_fd_sc_hd__nand2_1 _26962_ (.A(_06479_),
    .B(_06480_),
    .Y(_01311_));
 sky130_fd_sc_hd__nand2_1 _26963_ (.A(net1551),
    .B(_06438_),
    .Y(_06481_));
 sky130_fd_sc_hd__nand2_1 _26964_ (.A(\gen_regfile_ff.register_file_i.rf_reg[851] ),
    .B(_06441_),
    .Y(_06482_));
 sky130_fd_sc_hd__nand2_1 _26965_ (.A(_06481_),
    .B(_06482_),
    .Y(_01312_));
 sky130_fd_sc_hd__nand2_1 _26966_ (.A(_03614_),
    .B(_06112_),
    .Y(_06483_));
 sky130_fd_sc_hd__nand2_1 _26967_ (.A(\gen_regfile_ff.register_file_i.rf_reg[113] ),
    .B(_06115_),
    .Y(_06484_));
 sky130_fd_sc_hd__nand2_1 _26968_ (.A(_06483_),
    .B(_06484_),
    .Y(_01313_));
 sky130_fd_sc_hd__nand2_1 _26969_ (.A(_03982_),
    .B(_06438_),
    .Y(_06485_));
 sky130_fd_sc_hd__nand2_1 _26970_ (.A(\gen_regfile_ff.register_file_i.rf_reg[852] ),
    .B(_06441_),
    .Y(_06486_));
 sky130_fd_sc_hd__nand2_1 _26971_ (.A(_06485_),
    .B(_06486_),
    .Y(_01314_));
 sky130_fd_sc_hd__nand2_1 _26972_ (.A(net1584),
    .B(_06438_),
    .Y(_06487_));
 sky130_fd_sc_hd__nand2_1 _26973_ (.A(\gen_regfile_ff.register_file_i.rf_reg[853] ),
    .B(_06441_),
    .Y(_06488_));
 sky130_fd_sc_hd__nand2_1 _26974_ (.A(_06487_),
    .B(_06488_),
    .Y(_01315_));
 sky130_fd_sc_hd__mux2_4 _26975_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[854] ),
    .A1(net1517),
    .S(_06438_),
    .X(_01316_));
 sky130_fd_sc_hd__nand2_4 _26976_ (.A(net1290),
    .B(_06438_),
    .Y(_06489_));
 sky130_fd_sc_hd__nand2_1 _26977_ (.A(\gen_regfile_ff.register_file_i.rf_reg[855] ),
    .B(_06441_),
    .Y(_06490_));
 sky130_fd_sc_hd__nand2_2 _26978_ (.A(_06490_),
    .B(_06489_),
    .Y(_01317_));
 sky130_fd_sc_hd__nand2_1 _26979_ (.A(net1315),
    .B(_06438_),
    .Y(_06491_));
 sky130_fd_sc_hd__nand2_1 _26980_ (.A(\gen_regfile_ff.register_file_i.rf_reg[856] ),
    .B(_06441_),
    .Y(_06492_));
 sky130_fd_sc_hd__nand2_1 _26981_ (.A(_06492_),
    .B(_06491_),
    .Y(_01318_));
 sky130_fd_sc_hd__nand2_1 _26982_ (.A(net1564),
    .B(_06438_),
    .Y(_06493_));
 sky130_fd_sc_hd__nand2_1 _26983_ (.A(\gen_regfile_ff.register_file_i.rf_reg[857] ),
    .B(_06441_),
    .Y(_06494_));
 sky130_fd_sc_hd__nand2_1 _26984_ (.A(_06493_),
    .B(_06494_),
    .Y(_01319_));
 sky130_fd_sc_hd__nand2_4 _26985_ (.A(net1514),
    .B(_06438_),
    .Y(_06495_));
 sky130_fd_sc_hd__nand2_1 _26986_ (.A(\gen_regfile_ff.register_file_i.rf_reg[858] ),
    .B(_06441_),
    .Y(_06496_));
 sky130_fd_sc_hd__nand2_2 _26987_ (.A(_06495_),
    .B(_06496_),
    .Y(_01320_));
 sky130_fd_sc_hd__nand2_1 _26988_ (.A(net1529),
    .B(_06438_),
    .Y(_06497_));
 sky130_fd_sc_hd__nand2_1 _26989_ (.A(\gen_regfile_ff.register_file_i.rf_reg[859] ),
    .B(_06441_),
    .Y(_06498_));
 sky130_fd_sc_hd__nand2_1 _26990_ (.A(_06497_),
    .B(_06498_),
    .Y(_01321_));
 sky130_fd_sc_hd__mux2_4 _26991_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[860] ),
    .A1(net1294),
    .S(_06438_),
    .X(_01322_));
 sky130_fd_sc_hd__nor2_1 _26992_ (.A(_05084_),
    .B(_06441_),
    .Y(_06499_));
 sky130_fd_sc_hd__a22o_1 _26993_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[861] ),
    .A2(_06441_),
    .B1(net1246),
    .B2(_06499_),
    .X(_01323_));
 sky130_fd_sc_hd__nand2_1 _26994_ (.A(_03739_),
    .B(_06112_),
    .Y(_06500_));
 sky130_fd_sc_hd__nand2_1 _26995_ (.A(\gen_regfile_ff.register_file_i.rf_reg[114] ),
    .B(_06115_),
    .Y(_06501_));
 sky130_fd_sc_hd__nand2_1 _26996_ (.A(_06500_),
    .B(_06501_),
    .Y(_01324_));
 sky130_fd_sc_hd__mux2_4 _26997_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[862] ),
    .A1(net859),
    .S(_06438_),
    .X(_01325_));
 sky130_fd_sc_hd__nor2_1 _26998_ (.A(_05264_),
    .B(_06441_),
    .Y(_06502_));
 sky130_fd_sc_hd__a22o_1 _26999_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[863] ),
    .A2(_06441_),
    .B1(net740),
    .B2(_06502_),
    .X(_01326_));
 sky130_fd_sc_hd__nor2_8 _27000_ (.A(_05572_),
    .B(_06232_),
    .Y(_06503_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_51 ();
 sky130_fd_sc_hd__nand2_1 _27002_ (.A(_01909_),
    .B(_06503_),
    .Y(_06505_));
 sky130_fd_sc_hd__nand2_8 _27003_ (.A(net1253),
    .B(_06236_),
    .Y(_06506_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_50 ();
 sky130_fd_sc_hd__nand2_1 _27005_ (.A(\gen_regfile_ff.register_file_i.rf_reg[864] ),
    .B(_06506_),
    .Y(_06508_));
 sky130_fd_sc_hd__nand2_1 _27006_ (.A(_06505_),
    .B(_06508_),
    .Y(_01327_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_49 ();
 sky130_fd_sc_hd__nand2_1 _27008_ (.A(\gen_regfile_ff.register_file_i.rf_reg[865] ),
    .B(_06506_),
    .Y(_06510_));
 sky130_fd_sc_hd__o21ai_0 _27009_ (.A1(_05299_),
    .A2(_06506_),
    .B1(_06510_),
    .Y(_01328_));
 sky130_fd_sc_hd__nand2_1 _27010_ (.A(_05326_),
    .B(_06503_),
    .Y(_06511_));
 sky130_fd_sc_hd__nand2_1 _27011_ (.A(\gen_regfile_ff.register_file_i.rf_reg[866] ),
    .B(_06506_),
    .Y(_06512_));
 sky130_fd_sc_hd__nand2_1 _27012_ (.A(_06511_),
    .B(_06512_),
    .Y(_01329_));
 sky130_fd_sc_hd__nand2_1 _27013_ (.A(\gen_regfile_ff.register_file_i.rf_reg[867] ),
    .B(_06506_),
    .Y(_06513_));
 sky130_fd_sc_hd__o21ai_0 _27014_ (.A1(_05351_),
    .A2(_06506_),
    .B1(_06513_),
    .Y(_01330_));
 sky130_fd_sc_hd__nand2_1 _27015_ (.A(_02113_),
    .B(_06503_),
    .Y(_06514_));
 sky130_fd_sc_hd__nand2_1 _27016_ (.A(\gen_regfile_ff.register_file_i.rf_reg[868] ),
    .B(_06506_),
    .Y(_06515_));
 sky130_fd_sc_hd__nand2_1 _27017_ (.A(_06514_),
    .B(_06515_),
    .Y(_01331_));
 sky130_fd_sc_hd__nand2_1 _27018_ (.A(_02250_),
    .B(_06503_),
    .Y(_06516_));
 sky130_fd_sc_hd__nand2_1 _27019_ (.A(\gen_regfile_ff.register_file_i.rf_reg[869] ),
    .B(_06506_),
    .Y(_06517_));
 sky130_fd_sc_hd__nand2_1 _27020_ (.A(_06516_),
    .B(_06517_),
    .Y(_01332_));
 sky130_fd_sc_hd__nand2_1 _27021_ (.A(_02360_),
    .B(_06503_),
    .Y(_06518_));
 sky130_fd_sc_hd__nand2_1 _27022_ (.A(\gen_regfile_ff.register_file_i.rf_reg[870] ),
    .B(_06506_),
    .Y(_06519_));
 sky130_fd_sc_hd__nand2_1 _27023_ (.A(_06518_),
    .B(_06519_),
    .Y(_01333_));
 sky130_fd_sc_hd__nand2_1 _27024_ (.A(_02468_),
    .B(_06503_),
    .Y(_06520_));
 sky130_fd_sc_hd__nand2_1 _27025_ (.A(\gen_regfile_ff.register_file_i.rf_reg[871] ),
    .B(_06506_),
    .Y(_06521_));
 sky130_fd_sc_hd__nand2_1 _27026_ (.A(_06520_),
    .B(_06521_),
    .Y(_01334_));
 sky130_fd_sc_hd__nand2_1 _27027_ (.A(_03866_),
    .B(_06112_),
    .Y(_06522_));
 sky130_fd_sc_hd__nand2_1 _27028_ (.A(\gen_regfile_ff.register_file_i.rf_reg[115] ),
    .B(_06115_),
    .Y(_06523_));
 sky130_fd_sc_hd__nand2_1 _27029_ (.A(_06522_),
    .B(_06523_),
    .Y(_01335_));
 sky130_fd_sc_hd__nand2_1 _27030_ (.A(_02553_),
    .B(_06503_),
    .Y(_06524_));
 sky130_fd_sc_hd__nand2_1 _27031_ (.A(\gen_regfile_ff.register_file_i.rf_reg[872] ),
    .B(_06506_),
    .Y(_06525_));
 sky130_fd_sc_hd__nand2_1 _27032_ (.A(_06524_),
    .B(_06525_),
    .Y(_01336_));
 sky130_fd_sc_hd__nand2_1 _27033_ (.A(_02653_),
    .B(_06503_),
    .Y(_06526_));
 sky130_fd_sc_hd__nand2_1 _27034_ (.A(\gen_regfile_ff.register_file_i.rf_reg[873] ),
    .B(_06506_),
    .Y(_06527_));
 sky130_fd_sc_hd__nand2_1 _27035_ (.A(_06526_),
    .B(_06527_),
    .Y(_01337_));
 sky130_fd_sc_hd__nand2_1 _27036_ (.A(_02761_),
    .B(_06503_),
    .Y(_06528_));
 sky130_fd_sc_hd__nand2_1 _27037_ (.A(\gen_regfile_ff.register_file_i.rf_reg[874] ),
    .B(_06506_),
    .Y(_06529_));
 sky130_fd_sc_hd__nand2_1 _27038_ (.A(_06528_),
    .B(_06529_),
    .Y(_01338_));
 sky130_fd_sc_hd__nand2_1 _27039_ (.A(_02849_),
    .B(_06503_),
    .Y(_06530_));
 sky130_fd_sc_hd__nand2_1 _27040_ (.A(\gen_regfile_ff.register_file_i.rf_reg[875] ),
    .B(_06506_),
    .Y(_06531_));
 sky130_fd_sc_hd__nand2_1 _27041_ (.A(_06530_),
    .B(_06531_),
    .Y(_01339_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_48 ();
 sky130_fd_sc_hd__nand2_1 _27043_ (.A(_02974_),
    .B(_06503_),
    .Y(_06533_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_47 ();
 sky130_fd_sc_hd__nand2_1 _27045_ (.A(\gen_regfile_ff.register_file_i.rf_reg[876] ),
    .B(_06506_),
    .Y(_06535_));
 sky130_fd_sc_hd__nand2_1 _27046_ (.A(_06533_),
    .B(_06535_),
    .Y(_01340_));
 sky130_fd_sc_hd__nand2_1 _27047_ (.A(_03080_),
    .B(_06503_),
    .Y(_06536_));
 sky130_fd_sc_hd__nand2_1 _27048_ (.A(\gen_regfile_ff.register_file_i.rf_reg[877] ),
    .B(_06506_),
    .Y(_06537_));
 sky130_fd_sc_hd__nand2_1 _27049_ (.A(_06536_),
    .B(_06537_),
    .Y(_01341_));
 sky130_fd_sc_hd__nand2_1 _27050_ (.A(_03214_),
    .B(_06503_),
    .Y(_06538_));
 sky130_fd_sc_hd__nand2_1 _27051_ (.A(\gen_regfile_ff.register_file_i.rf_reg[878] ),
    .B(_06506_),
    .Y(_06539_));
 sky130_fd_sc_hd__nand2_1 _27052_ (.A(_06538_),
    .B(_06539_),
    .Y(_01342_));
 sky130_fd_sc_hd__nand2_1 _27053_ (.A(_03348_),
    .B(_06503_),
    .Y(_06540_));
 sky130_fd_sc_hd__nand2_1 _27054_ (.A(\gen_regfile_ff.register_file_i.rf_reg[879] ),
    .B(_06506_),
    .Y(_06541_));
 sky130_fd_sc_hd__nand2_1 _27055_ (.A(_06540_),
    .B(_06541_),
    .Y(_01343_));
 sky130_fd_sc_hd__nand2_1 _27056_ (.A(\gen_regfile_ff.register_file_i.rf_reg[880] ),
    .B(_06506_),
    .Y(_06542_));
 sky130_fd_sc_hd__o21ai_0 _27057_ (.A1(_03481_),
    .A2(_06506_),
    .B1(_06542_),
    .Y(_01344_));
 sky130_fd_sc_hd__nand2_1 _27058_ (.A(net1575),
    .B(_06503_),
    .Y(_06543_));
 sky130_fd_sc_hd__nand2_1 _27059_ (.A(\gen_regfile_ff.register_file_i.rf_reg[881] ),
    .B(_06506_),
    .Y(_06544_));
 sky130_fd_sc_hd__nand2_1 _27060_ (.A(_06543_),
    .B(_06544_),
    .Y(_01345_));
 sky130_fd_sc_hd__nand2_1 _27061_ (.A(_03982_),
    .B(_06112_),
    .Y(_06545_));
 sky130_fd_sc_hd__nand2_1 _27062_ (.A(\gen_regfile_ff.register_file_i.rf_reg[116] ),
    .B(_06115_),
    .Y(_06546_));
 sky130_fd_sc_hd__nand2_1 _27063_ (.A(_06545_),
    .B(_06546_),
    .Y(_01346_));
 sky130_fd_sc_hd__nand2_1 _27064_ (.A(net1576),
    .B(_06503_),
    .Y(_06547_));
 sky130_fd_sc_hd__nand2_1 _27065_ (.A(\gen_regfile_ff.register_file_i.rf_reg[882] ),
    .B(_06506_),
    .Y(_06548_));
 sky130_fd_sc_hd__nand2_1 _27066_ (.A(_06547_),
    .B(_06548_),
    .Y(_01347_));
 sky130_fd_sc_hd__nand2_1 _27067_ (.A(_03866_),
    .B(_06503_),
    .Y(_06549_));
 sky130_fd_sc_hd__nand2_1 _27068_ (.A(\gen_regfile_ff.register_file_i.rf_reg[883] ),
    .B(_06506_),
    .Y(_06550_));
 sky130_fd_sc_hd__nand2_1 _27069_ (.A(_06549_),
    .B(_06550_),
    .Y(_01348_));
 sky130_fd_sc_hd__nand2_1 _27070_ (.A(net1544),
    .B(_06503_),
    .Y(_06551_));
 sky130_fd_sc_hd__nand2_1 _27071_ (.A(\gen_regfile_ff.register_file_i.rf_reg[884] ),
    .B(_06506_),
    .Y(_06552_));
 sky130_fd_sc_hd__nand2_1 _27072_ (.A(_06551_),
    .B(_06552_),
    .Y(_01349_));
 sky130_fd_sc_hd__nand2_1 _27073_ (.A(net1584),
    .B(_06503_),
    .Y(_06553_));
 sky130_fd_sc_hd__nand2_1 _27074_ (.A(\gen_regfile_ff.register_file_i.rf_reg[885] ),
    .B(_06506_),
    .Y(_06554_));
 sky130_fd_sc_hd__nand2_1 _27075_ (.A(_06553_),
    .B(_06554_),
    .Y(_01350_));
 sky130_fd_sc_hd__mux2_4 _27076_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[886] ),
    .A1(_04252_),
    .S(_06503_),
    .X(_01351_));
 sky130_fd_sc_hd__nand2_2 _27077_ (.A(net1523),
    .B(_06503_),
    .Y(_06555_));
 sky130_fd_sc_hd__nand2_1 _27078_ (.A(\gen_regfile_ff.register_file_i.rf_reg[887] ),
    .B(_06506_),
    .Y(_06556_));
 sky130_fd_sc_hd__nand2_1 _27079_ (.A(_06556_),
    .B(_06555_),
    .Y(_01352_));
 sky130_fd_sc_hd__nand2_4 _27080_ (.A(net1271),
    .B(_06503_),
    .Y(_06557_));
 sky130_fd_sc_hd__nand2_1 _27081_ (.A(\gen_regfile_ff.register_file_i.rf_reg[888] ),
    .B(_06506_),
    .Y(_06558_));
 sky130_fd_sc_hd__nand2_2 _27082_ (.A(_06557_),
    .B(_06558_),
    .Y(_01353_));
 sky130_fd_sc_hd__nand2_1 _27083_ (.A(net252),
    .B(_06503_),
    .Y(_06559_));
 sky130_fd_sc_hd__nand2_1 _27084_ (.A(\gen_regfile_ff.register_file_i.rf_reg[889] ),
    .B(_06506_),
    .Y(_06560_));
 sky130_fd_sc_hd__nand2_1 _27085_ (.A(_06559_),
    .B(_06560_),
    .Y(_01354_));
 sky130_fd_sc_hd__nand2_2 _27086_ (.A(net1536),
    .B(_06503_),
    .Y(_06561_));
 sky130_fd_sc_hd__nand2_1 _27087_ (.A(\gen_regfile_ff.register_file_i.rf_reg[890] ),
    .B(_06506_),
    .Y(_06562_));
 sky130_fd_sc_hd__nand2_1 _27088_ (.A(_06561_),
    .B(_06562_),
    .Y(_01355_));
 sky130_fd_sc_hd__nand2_2 _27089_ (.A(net1529),
    .B(_06503_),
    .Y(_06563_));
 sky130_fd_sc_hd__nand2_1 _27090_ (.A(\gen_regfile_ff.register_file_i.rf_reg[891] ),
    .B(_06506_),
    .Y(_06564_));
 sky130_fd_sc_hd__nand2_1 _27091_ (.A(_06563_),
    .B(_06564_),
    .Y(_01356_));
 sky130_fd_sc_hd__nand2_1 _27092_ (.A(net1017),
    .B(_06112_),
    .Y(_06565_));
 sky130_fd_sc_hd__nand2_1 _27093_ (.A(\gen_regfile_ff.register_file_i.rf_reg[117] ),
    .B(_06115_),
    .Y(_06566_));
 sky130_fd_sc_hd__nand2_1 _27094_ (.A(_06565_),
    .B(_06566_),
    .Y(_01357_));
 sky130_fd_sc_hd__mux2_4 _27095_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[892] ),
    .A1(net886),
    .S(_06503_),
    .X(_01358_));
 sky130_fd_sc_hd__nor2_1 _27096_ (.A(_05084_),
    .B(_06506_),
    .Y(_06567_));
 sky130_fd_sc_hd__a22o_1 _27097_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[893] ),
    .A2(_06506_),
    .B1(net1249),
    .B2(_06567_),
    .X(_01359_));
 sky130_fd_sc_hd__mux2_4 _27098_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[894] ),
    .A1(net685),
    .S(_06503_),
    .X(_01360_));
 sky130_fd_sc_hd__nor2_1 _27099_ (.A(_05264_),
    .B(_06506_),
    .Y(_06568_));
 sky130_fd_sc_hd__a22o_1 _27100_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[895] ),
    .A2(_06506_),
    .B1(_06568_),
    .B2(net500),
    .X(_01361_));
 sky130_fd_sc_hd__nand3_4 _27101_ (.A(_05847_),
    .B(_05955_),
    .C(net446),
    .Y(_06569_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_45 ();
 sky130_fd_sc_hd__nand2_1 _27104_ (.A(\gen_regfile_ff.register_file_i.rf_reg[896] ),
    .B(net1482),
    .Y(_06572_));
 sky130_fd_sc_hd__o31ai_1 _27105_ (.A1(_01732_),
    .A2(net258),
    .A3(net1482),
    .B1(_06572_),
    .Y(_01362_));
 sky130_fd_sc_hd__nand2_1 _27106_ (.A(\gen_regfile_ff.register_file_i.rf_reg[897] ),
    .B(net1482),
    .Y(_06573_));
 sky130_fd_sc_hd__o21ai_0 _27107_ (.A1(_05299_),
    .A2(net1482),
    .B1(_06573_),
    .Y(_01363_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_44 ();
 sky130_fd_sc_hd__mux2_1 _27109_ (.A0(_05326_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[898] ),
    .S(_06569_),
    .X(_01364_));
 sky130_fd_sc_hd__nand2_1 _27110_ (.A(\gen_regfile_ff.register_file_i.rf_reg[899] ),
    .B(net1482),
    .Y(_06575_));
 sky130_fd_sc_hd__o21ai_0 _27111_ (.A1(_05351_),
    .A2(net1482),
    .B1(_06575_),
    .Y(_01365_));
 sky130_fd_sc_hd__mux2_1 _27112_ (.A0(_02113_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[900] ),
    .S(net1482),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _27113_ (.A0(_02250_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[901] ),
    .S(_06569_),
    .X(_01367_));
 sky130_fd_sc_hd__mux2_4 _27114_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[118] ),
    .A1(net1326),
    .S(_06112_),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _27115_ (.A0(_02360_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[902] ),
    .S(net1482),
    .X(_01369_));
 sky130_fd_sc_hd__mux2_1 _27116_ (.A0(_02468_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[903] ),
    .S(_06569_),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_1 _27117_ (.A0(_02553_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[904] ),
    .S(_06569_),
    .X(_01371_));
 sky130_fd_sc_hd__mux2_1 _27118_ (.A0(_02653_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[905] ),
    .S(_06569_),
    .X(_01372_));
 sky130_fd_sc_hd__mux2_1 _27119_ (.A0(_02761_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[906] ),
    .S(_06569_),
    .X(_01373_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_43 ();
 sky130_fd_sc_hd__mux2_1 _27121_ (.A0(_02849_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[907] ),
    .S(_06569_),
    .X(_01374_));
 sky130_fd_sc_hd__mux2_1 _27122_ (.A0(_02974_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[908] ),
    .S(_06569_),
    .X(_01375_));
 sky130_fd_sc_hd__mux2_1 _27123_ (.A0(_03080_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[909] ),
    .S(_06569_),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_1 _27124_ (.A0(_03214_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[910] ),
    .S(_06569_),
    .X(_01377_));
 sky130_fd_sc_hd__mux2_1 _27125_ (.A0(_03348_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[911] ),
    .S(_06569_),
    .X(_01378_));
 sky130_fd_sc_hd__nand2_2 _27126_ (.A(net1291),
    .B(_06112_),
    .Y(_06577_));
 sky130_fd_sc_hd__nand2_1 _27127_ (.A(\gen_regfile_ff.register_file_i.rf_reg[119] ),
    .B(_06115_),
    .Y(_06578_));
 sky130_fd_sc_hd__nand2_1 _27128_ (.A(_06577_),
    .B(_06578_),
    .Y(_01379_));
 sky130_fd_sc_hd__nand2_1 _27129_ (.A(\gen_regfile_ff.register_file_i.rf_reg[912] ),
    .B(net1482),
    .Y(_06579_));
 sky130_fd_sc_hd__o21ai_0 _27130_ (.A1(_03481_),
    .A2(net1482),
    .B1(_06579_),
    .Y(_01380_));
 sky130_fd_sc_hd__mux2_1 _27131_ (.A0(net1575),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[913] ),
    .S(net1482),
    .X(_01381_));
 sky130_fd_sc_hd__mux2_1 _27132_ (.A0(net1576),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[914] ),
    .S(net1482),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _27133_ (.A0(net1551),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[915] ),
    .S(_06569_),
    .X(_01383_));
 sky130_fd_sc_hd__mux2_4 _27134_ (.A0(net1537),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[916] ),
    .S(_06569_),
    .X(_01384_));
 sky130_fd_sc_hd__mux2_1 _27135_ (.A0(net1017),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[917] ),
    .S(_06569_),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_4 _27136_ (.A0(net1327),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[918] ),
    .S(_06569_),
    .X(_01386_));
 sky130_fd_sc_hd__mux2_4 _27137_ (.A0(net1504),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[919] ),
    .S(net1482),
    .X(_01387_));
 sky130_fd_sc_hd__mux2_4 _27138_ (.A0(net1317),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[920] ),
    .S(_06569_),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _27139_ (.A0(net252),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[921] ),
    .S(_06569_),
    .X(_01389_));
 sky130_fd_sc_hd__nand2_2 _27140_ (.A(net1270),
    .B(_06112_),
    .Y(_06580_));
 sky130_fd_sc_hd__nand2_1 _27141_ (.A(\gen_regfile_ff.register_file_i.rf_reg[120] ),
    .B(_06115_),
    .Y(_06581_));
 sky130_fd_sc_hd__nand2_1 _27142_ (.A(_06580_),
    .B(_06581_),
    .Y(_01390_));
 sky130_fd_sc_hd__mux2_4 _27143_ (.A0(net251),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[922] ),
    .S(net1482),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_4 _27144_ (.A0(_04865_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[923] ),
    .S(_06569_),
    .X(_01392_));
 sky130_fd_sc_hd__mux2_4 _27145_ (.A0(net1294),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[924] ),
    .S(_06569_),
    .X(_01393_));
 sky130_fd_sc_hd__nor2_1 _27146_ (.A(_05084_),
    .B(net1482),
    .Y(_06582_));
 sky130_fd_sc_hd__a22o_1 _27147_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[925] ),
    .A2(net1482),
    .B1(net1254),
    .B2(_06582_),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_4 _27148_ (.A0(net859),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[926] ),
    .S(net1482),
    .X(_01395_));
 sky130_fd_sc_hd__nor2_1 _27149_ (.A(_05264_),
    .B(net1482),
    .Y(_06583_));
 sky130_fd_sc_hd__a22o_1 _27150_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[927] ),
    .A2(net1482),
    .B1(net500),
    .B2(_06583_),
    .X(_01396_));
 sky130_fd_sc_hd__nand3_4 _27151_ (.A(_05847_),
    .B(_01919_),
    .C(net447),
    .Y(_06584_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_41 ();
 sky130_fd_sc_hd__nand2_1 _27154_ (.A(\gen_regfile_ff.register_file_i.rf_reg[928] ),
    .B(net1481),
    .Y(_06587_));
 sky130_fd_sc_hd__o31ai_1 _27155_ (.A1(_01732_),
    .A2(net258),
    .A3(net1481),
    .B1(_06587_),
    .Y(_01397_));
 sky130_fd_sc_hd__nand2_1 _27156_ (.A(\gen_regfile_ff.register_file_i.rf_reg[929] ),
    .B(net1481),
    .Y(_06588_));
 sky130_fd_sc_hd__o21ai_0 _27157_ (.A1(_05299_),
    .A2(net1481),
    .B1(_06588_),
    .Y(_01398_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_40 ();
 sky130_fd_sc_hd__mux2_1 _27159_ (.A0(_05326_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[930] ),
    .S(_06584_),
    .X(_01399_));
 sky130_fd_sc_hd__nand2_1 _27160_ (.A(\gen_regfile_ff.register_file_i.rf_reg[931] ),
    .B(net1481),
    .Y(_06590_));
 sky130_fd_sc_hd__o21ai_0 _27161_ (.A1(_05351_),
    .A2(net1481),
    .B1(_06590_),
    .Y(_01400_));
 sky130_fd_sc_hd__nand2_4 _27162_ (.A(net1564),
    .B(_06112_),
    .Y(_06591_));
 sky130_fd_sc_hd__nand2_1 _27163_ (.A(\gen_regfile_ff.register_file_i.rf_reg[121] ),
    .B(_06115_),
    .Y(_06592_));
 sky130_fd_sc_hd__nand2_1 _27164_ (.A(_06591_),
    .B(_06592_),
    .Y(_01401_));
 sky130_fd_sc_hd__nand2_1 _27165_ (.A(_01916_),
    .B(_02553_),
    .Y(_06593_));
 sky130_fd_sc_hd__nand2_1 _27166_ (.A(\gen_regfile_ff.register_file_i.rf_reg[40] ),
    .B(_01921_),
    .Y(_06594_));
 sky130_fd_sc_hd__nand2_1 _27167_ (.A(_06593_),
    .B(_06594_),
    .Y(_01402_));
 sky130_fd_sc_hd__mux2_1 _27168_ (.A0(_02113_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[932] ),
    .S(net1481),
    .X(_01403_));
 sky130_fd_sc_hd__mux2_1 _27169_ (.A0(_02250_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[933] ),
    .S(_06584_),
    .X(_01404_));
 sky130_fd_sc_hd__mux2_1 _27170_ (.A0(_02360_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[934] ),
    .S(_06584_),
    .X(_01405_));
 sky130_fd_sc_hd__mux2_1 _27171_ (.A0(_02468_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[935] ),
    .S(_06584_),
    .X(_01406_));
 sky130_fd_sc_hd__mux2_1 _27172_ (.A0(_02553_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[936] ),
    .S(_06584_),
    .X(_01407_));
 sky130_fd_sc_hd__mux2_1 _27173_ (.A0(_02653_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[937] ),
    .S(_06584_),
    .X(_01408_));
 sky130_fd_sc_hd__mux2_1 _27174_ (.A0(_02761_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[938] ),
    .S(_06584_),
    .X(_01409_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_39 ();
 sky130_fd_sc_hd__mux2_1 _27176_ (.A0(_02849_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[939] ),
    .S(_06584_),
    .X(_01410_));
 sky130_fd_sc_hd__mux2_1 _27177_ (.A0(_02974_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[940] ),
    .S(_06584_),
    .X(_01411_));
 sky130_fd_sc_hd__mux2_1 _27178_ (.A0(_03080_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[941] ),
    .S(net1481),
    .X(_01412_));
 sky130_fd_sc_hd__nand2_4 _27179_ (.A(net1515),
    .B(_06112_),
    .Y(_06596_));
 sky130_fd_sc_hd__nand2_1 _27180_ (.A(\gen_regfile_ff.register_file_i.rf_reg[122] ),
    .B(_06115_),
    .Y(_06597_));
 sky130_fd_sc_hd__nand2_2 _27181_ (.A(_06596_),
    .B(_06597_),
    .Y(_01413_));
 sky130_fd_sc_hd__mux2_1 _27182_ (.A0(_03214_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[942] ),
    .S(_06584_),
    .X(_01414_));
 sky130_fd_sc_hd__mux2_1 _27183_ (.A0(_03348_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[943] ),
    .S(_06584_),
    .X(_01415_));
 sky130_fd_sc_hd__nand2_1 _27184_ (.A(\gen_regfile_ff.register_file_i.rf_reg[944] ),
    .B(net1481),
    .Y(_06598_));
 sky130_fd_sc_hd__o21ai_0 _27185_ (.A1(_03481_),
    .A2(net1481),
    .B1(_06598_),
    .Y(_01416_));
 sky130_fd_sc_hd__mux2_1 _27186_ (.A0(net1575),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[945] ),
    .S(net1481),
    .X(_01417_));
 sky130_fd_sc_hd__mux2_1 _27187_ (.A0(_03739_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[946] ),
    .S(_06584_),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_1 _27188_ (.A0(net1551),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[947] ),
    .S(net1481),
    .X(_01419_));
 sky130_fd_sc_hd__mux2_1 _27189_ (.A0(net1537),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[948] ),
    .S(_06584_),
    .X(_01420_));
 sky130_fd_sc_hd__mux2_1 _27190_ (.A0(net1017),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[949] ),
    .S(net1481),
    .X(_01421_));
 sky130_fd_sc_hd__mux2_4 _27191_ (.A0(net1517),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[950] ),
    .S(_06584_),
    .X(_01422_));
 sky130_fd_sc_hd__mux2_4 _27192_ (.A0(net1475),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[951] ),
    .S(_06584_),
    .X(_01423_));
 sky130_fd_sc_hd__nand2_1 _27193_ (.A(net1540),
    .B(_06112_),
    .Y(_06599_));
 sky130_fd_sc_hd__nand2_1 _27194_ (.A(\gen_regfile_ff.register_file_i.rf_reg[123] ),
    .B(_06115_),
    .Y(_06600_));
 sky130_fd_sc_hd__nand2_1 _27195_ (.A(_06599_),
    .B(_06600_),
    .Y(_01424_));
 sky130_fd_sc_hd__mux2_4 _27196_ (.A0(net1316),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[952] ),
    .S(_06584_),
    .X(_01425_));
 sky130_fd_sc_hd__mux2_1 _27197_ (.A0(net252),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[953] ),
    .S(_06584_),
    .X(_01426_));
 sky130_fd_sc_hd__mux2_4 _27198_ (.A0(net251),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[954] ),
    .S(_06584_),
    .X(_01427_));
 sky130_fd_sc_hd__mux2_4 _27199_ (.A0(_04865_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[955] ),
    .S(_06584_),
    .X(_01428_));
 sky130_fd_sc_hd__mux2_4 _27200_ (.A0(net1294),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[956] ),
    .S(net1481),
    .X(_01429_));
 sky130_fd_sc_hd__nor2_1 _27201_ (.A(_05084_),
    .B(net1481),
    .Y(_06601_));
 sky130_fd_sc_hd__a22o_1 _27202_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[957] ),
    .A2(net1481),
    .B1(net1246),
    .B2(_06601_),
    .X(_01430_));
 sky130_fd_sc_hd__mux2_4 _27203_ (.A0(net859),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[958] ),
    .S(net1481),
    .X(_01431_));
 sky130_fd_sc_hd__nor2_1 _27204_ (.A(_05264_),
    .B(net1481),
    .Y(_06602_));
 sky130_fd_sc_hd__a22o_1 _27205_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[959] ),
    .A2(net1481),
    .B1(net957),
    .B2(_06602_),
    .X(_01432_));
 sky130_fd_sc_hd__nand3_4 _27206_ (.A(_05847_),
    .B(_05796_),
    .C(net447),
    .Y(_06603_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_37 ();
 sky130_fd_sc_hd__nand2_1 _27209_ (.A(\gen_regfile_ff.register_file_i.rf_reg[960] ),
    .B(net1480),
    .Y(_06606_));
 sky130_fd_sc_hd__o31ai_1 _27210_ (.A1(_01732_),
    .A2(net258),
    .A3(net1480),
    .B1(_06606_),
    .Y(_01433_));
 sky130_fd_sc_hd__nand2_1 _27211_ (.A(\gen_regfile_ff.register_file_i.rf_reg[961] ),
    .B(net1480),
    .Y(_06607_));
 sky130_fd_sc_hd__o21ai_0 _27212_ (.A1(_05299_),
    .A2(net1480),
    .B1(_06607_),
    .Y(_01434_));
 sky130_fd_sc_hd__mux2_4 _27213_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[124] ),
    .A1(_04975_),
    .S(_06112_),
    .X(_01435_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_36 ();
 sky130_fd_sc_hd__mux2_1 _27215_ (.A0(_05326_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[962] ),
    .S(_06603_),
    .X(_01436_));
 sky130_fd_sc_hd__nand2_1 _27216_ (.A(\gen_regfile_ff.register_file_i.rf_reg[963] ),
    .B(net1480),
    .Y(_06609_));
 sky130_fd_sc_hd__o21ai_0 _27217_ (.A1(_05351_),
    .A2(net1480),
    .B1(_06609_),
    .Y(_01437_));
 sky130_fd_sc_hd__mux2_1 _27218_ (.A0(_02113_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[964] ),
    .S(_06603_),
    .X(_01438_));
 sky130_fd_sc_hd__mux2_1 _27219_ (.A0(_02250_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[965] ),
    .S(_06603_),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _27220_ (.A0(_02360_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[966] ),
    .S(net1480),
    .X(_01440_));
 sky130_fd_sc_hd__mux2_1 _27221_ (.A0(_02468_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[967] ),
    .S(_06603_),
    .X(_01441_));
 sky130_fd_sc_hd__mux2_1 _27222_ (.A0(_02553_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[968] ),
    .S(_06603_),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_1 _27223_ (.A0(_02653_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[969] ),
    .S(net1480),
    .X(_01443_));
 sky130_fd_sc_hd__mux2_1 _27224_ (.A0(_02761_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[970] ),
    .S(_06603_),
    .X(_01444_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_35 ();
 sky130_fd_sc_hd__mux2_1 _27226_ (.A0(_02849_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[971] ),
    .S(_06603_),
    .X(_01445_));
 sky130_fd_sc_hd__nor2_1 _27227_ (.A(_05084_),
    .B(_06115_),
    .Y(_06611_));
 sky130_fd_sc_hd__a22o_1 _27228_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[125] ),
    .A2(_06115_),
    .B1(_05079_),
    .B2(_06611_),
    .X(_01446_));
 sky130_fd_sc_hd__mux2_1 _27229_ (.A0(_02974_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[972] ),
    .S(_06603_),
    .X(_01447_));
 sky130_fd_sc_hd__mux2_1 _27230_ (.A0(_03080_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[973] ),
    .S(net1480),
    .X(_01448_));
 sky130_fd_sc_hd__mux2_1 _27231_ (.A0(_03214_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[974] ),
    .S(_06603_),
    .X(_01449_));
 sky130_fd_sc_hd__mux2_1 _27232_ (.A0(_03348_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[975] ),
    .S(_06603_),
    .X(_01450_));
 sky130_fd_sc_hd__nand2_1 _27233_ (.A(\gen_regfile_ff.register_file_i.rf_reg[976] ),
    .B(net1480),
    .Y(_06612_));
 sky130_fd_sc_hd__o21ai_0 _27234_ (.A1(_03481_),
    .A2(net1480),
    .B1(_06612_),
    .Y(_01451_));
 sky130_fd_sc_hd__mux2_1 _27235_ (.A0(net1575),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[977] ),
    .S(net1480),
    .X(_01452_));
 sky130_fd_sc_hd__mux2_1 _27236_ (.A0(net1576),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[978] ),
    .S(_06603_),
    .X(_01453_));
 sky130_fd_sc_hd__mux2_1 _27237_ (.A0(_03866_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[979] ),
    .S(_06603_),
    .X(_01454_));
 sky130_fd_sc_hd__mux2_4 _27238_ (.A0(net1537),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[980] ),
    .S(_06603_),
    .X(_01455_));
 sky130_fd_sc_hd__mux2_1 _27239_ (.A0(net1017),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[981] ),
    .S(_06603_),
    .X(_01456_));
 sky130_fd_sc_hd__mux2_4 _27240_ (.A0(\gen_regfile_ff.register_file_i.rf_reg[126] ),
    .A1(net1237),
    .S(_06112_),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_4 _27241_ (.A0(net1327),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[982] ),
    .S(_06603_),
    .X(_01458_));
 sky130_fd_sc_hd__mux2_4 _27242_ (.A0(net1475),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[983] ),
    .S(_06603_),
    .X(_01459_));
 sky130_fd_sc_hd__mux2_4 _27243_ (.A0(net1316),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[984] ),
    .S(_06603_),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _27244_ (.A0(net252),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[985] ),
    .S(_06603_),
    .X(_01461_));
 sky130_fd_sc_hd__mux2_4 _27245_ (.A0(net251),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[986] ),
    .S(net1480),
    .X(_01462_));
 sky130_fd_sc_hd__mux2_4 _27246_ (.A0(_04865_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[987] ),
    .S(_06603_),
    .X(_01463_));
 sky130_fd_sc_hd__mux2_4 _27247_ (.A0(net250),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[988] ),
    .S(net1480),
    .X(_01464_));
 sky130_fd_sc_hd__nor2_1 _27248_ (.A(_05084_),
    .B(net1480),
    .Y(_06613_));
 sky130_fd_sc_hd__a22o_1 _27249_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[989] ),
    .A2(net1480),
    .B1(net1249),
    .B2(_06613_),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_4 _27250_ (.A0(net685),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[990] ),
    .S(net1480),
    .X(_01466_));
 sky130_fd_sc_hd__nor2_1 _27251_ (.A(_05264_),
    .B(net1480),
    .Y(_06614_));
 sky130_fd_sc_hd__a22o_1 _27252_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[991] ),
    .A2(net1480),
    .B1(_06614_),
    .B2(net500),
    .X(_01467_));
 sky130_fd_sc_hd__nor2_1 _27253_ (.A(_05264_),
    .B(_06115_),
    .Y(_06615_));
 sky130_fd_sc_hd__a22o_1 _27254_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[127] ),
    .A2(_06115_),
    .B1(_06615_),
    .B2(net740),
    .X(_01468_));
 sky130_fd_sc_hd__nand2_8 _27255_ (.A(_05847_),
    .B(_06236_),
    .Y(_06616_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_33 ();
 sky130_fd_sc_hd__nand2_1 _27258_ (.A(\gen_regfile_ff.register_file_i.rf_reg[992] ),
    .B(_06616_),
    .Y(_06619_));
 sky130_fd_sc_hd__o31ai_1 _27259_ (.A1(_01732_),
    .A2(net258),
    .A3(_06616_),
    .B1(_06619_),
    .Y(_01469_));
 sky130_fd_sc_hd__nand2_1 _27260_ (.A(\gen_regfile_ff.register_file_i.rf_reg[993] ),
    .B(_06616_),
    .Y(_06620_));
 sky130_fd_sc_hd__o21ai_0 _27261_ (.A1(_05299_),
    .A2(_06616_),
    .B1(_06620_),
    .Y(_01470_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_32 ();
 sky130_fd_sc_hd__mux2_1 _27263_ (.A0(_05326_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[994] ),
    .S(_06616_),
    .X(_01471_));
 sky130_fd_sc_hd__nand2_1 _27264_ (.A(\gen_regfile_ff.register_file_i.rf_reg[995] ),
    .B(_06616_),
    .Y(_06622_));
 sky130_fd_sc_hd__o21ai_0 _27265_ (.A1(_05351_),
    .A2(_06616_),
    .B1(_06622_),
    .Y(_01472_));
 sky130_fd_sc_hd__mux2_1 _27266_ (.A0(_02113_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[996] ),
    .S(_06616_),
    .X(_01473_));
 sky130_fd_sc_hd__mux2_1 _27267_ (.A0(_02250_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[997] ),
    .S(_06616_),
    .X(_01474_));
 sky130_fd_sc_hd__mux2_1 _27268_ (.A0(_02360_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[998] ),
    .S(_06616_),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _27269_ (.A0(_02468_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[999] ),
    .S(_06616_),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_1 _27270_ (.A0(_02553_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1000] ),
    .S(_06616_),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_1 _27271_ (.A0(_02653_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1001] ),
    .S(_06616_),
    .X(_01478_));
 sky130_fd_sc_hd__nand2_1 _27272_ (.A(_01909_),
    .B(_02119_),
    .Y(_06623_));
 sky130_fd_sc_hd__nand2_1 _27273_ (.A(\gen_regfile_ff.register_file_i.rf_reg[128] ),
    .B(_02123_),
    .Y(_06624_));
 sky130_fd_sc_hd__nand2_1 _27274_ (.A(_06623_),
    .B(_06624_),
    .Y(_01479_));
 sky130_fd_sc_hd__mux2_1 _27275_ (.A0(_02761_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1002] ),
    .S(_06616_),
    .X(_01480_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_31 ();
 sky130_fd_sc_hd__mux2_1 _27277_ (.A0(_02849_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1003] ),
    .S(_06616_),
    .X(_01481_));
 sky130_fd_sc_hd__mux2_1 _27278_ (.A0(_02974_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1004] ),
    .S(_06616_),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_1 _27279_ (.A0(_03080_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1005] ),
    .S(_06616_),
    .X(_01483_));
 sky130_fd_sc_hd__mux2_1 _27280_ (.A0(_03214_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1006] ),
    .S(_06616_),
    .X(_01484_));
 sky130_fd_sc_hd__mux2_1 _27281_ (.A0(_03348_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1007] ),
    .S(_06616_),
    .X(_01485_));
 sky130_fd_sc_hd__nand2_1 _27282_ (.A(\gen_regfile_ff.register_file_i.rf_reg[1008] ),
    .B(_06616_),
    .Y(_06626_));
 sky130_fd_sc_hd__o21ai_0 _27283_ (.A1(_03481_),
    .A2(_06616_),
    .B1(_06626_),
    .Y(_01486_));
 sky130_fd_sc_hd__mux2_1 _27284_ (.A0(net1575),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1009] ),
    .S(_06616_),
    .X(_01487_));
 sky130_fd_sc_hd__mux2_1 _27285_ (.A0(_03739_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1010] ),
    .S(_06616_),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_1 _27286_ (.A0(_03866_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1011] ),
    .S(_06616_),
    .X(_01489_));
 sky130_fd_sc_hd__nand2_1 _27287_ (.A(\gen_regfile_ff.register_file_i.rf_reg[129] ),
    .B(_02123_),
    .Y(_06627_));
 sky130_fd_sc_hd__o21ai_0 _27288_ (.A1(_02123_),
    .A2(_05299_),
    .B1(_06627_),
    .Y(_01490_));
 sky130_fd_sc_hd__mux2_4 _27289_ (.A0(net1537),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1012] ),
    .S(_06616_),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_1 _27290_ (.A0(net1017),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1013] ),
    .S(_06616_),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_4 _27291_ (.A0(net1327),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1014] ),
    .S(_06616_),
    .X(_01493_));
 sky130_fd_sc_hd__mux2_4 _27292_ (.A0(net1290),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1015] ),
    .S(_06616_),
    .X(_01494_));
 sky130_fd_sc_hd__mux2_4 _27293_ (.A0(net1317),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1016] ),
    .S(_06616_),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _27294_ (.A0(net252),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1017] ),
    .S(_06616_),
    .X(_01496_));
 sky130_fd_sc_hd__mux2_4 _27295_ (.A0(net1515),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1018] ),
    .S(_06616_),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_4 _27296_ (.A0(_04865_),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1019] ),
    .S(_06616_),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_4 _27297_ (.A0(net1294),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1020] ),
    .S(_06616_),
    .X(_01499_));
 sky130_fd_sc_hd__nor2_1 _27298_ (.A(_05084_),
    .B(_06616_),
    .Y(_06628_));
 sky130_fd_sc_hd__a22o_1 _27299_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[1021] ),
    .A2(_06616_),
    .B1(net1246),
    .B2(_06628_),
    .X(_01500_));
 sky130_fd_sc_hd__nand2_1 _27300_ (.A(_02119_),
    .B(_05326_),
    .Y(_06629_));
 sky130_fd_sc_hd__nand2_1 _27301_ (.A(\gen_regfile_ff.register_file_i.rf_reg[130] ),
    .B(_02123_),
    .Y(_06630_));
 sky130_fd_sc_hd__nand2_1 _27302_ (.A(_06629_),
    .B(_06630_),
    .Y(_01501_));
 sky130_fd_sc_hd__mux2_4 _27303_ (.A0(net859),
    .A1(\gen_regfile_ff.register_file_i.rf_reg[1022] ),
    .S(_06616_),
    .X(_01502_));
 sky130_fd_sc_hd__nor2_1 _27304_ (.A(_05264_),
    .B(_06616_),
    .Y(_06631_));
 sky130_fd_sc_hd__a22o_1 _27305_ (.A1(\gen_regfile_ff.register_file_i.rf_reg[1023] ),
    .A2(_06616_),
    .B1(net957),
    .B2(_06631_),
    .X(_01503_));
 sky130_fd_sc_hd__nand2_1 _27306_ (.A(\gen_regfile_ff.register_file_i.rf_reg[131] ),
    .B(_02123_),
    .Y(_06632_));
 sky130_fd_sc_hd__o21ai_0 _27307_ (.A1(_02123_),
    .A2(_05351_),
    .B1(_06632_),
    .Y(_01504_));
 sky130_fd_sc_hd__nand2_1 _27308_ (.A(_01916_),
    .B(_02653_),
    .Y(_06633_));
 sky130_fd_sc_hd__nand2_1 _27309_ (.A(\gen_regfile_ff.register_file_i.rf_reg[41] ),
    .B(_01921_),
    .Y(_06634_));
 sky130_fd_sc_hd__dfrtp_4 _27310_ (.D(_00008_),
    .Q(\load_store_unit_i.data_type_q[2] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfrtp_4 _27311_ (.D(_00009_),
    .Q(\load_store_unit_i.data_type_q[1] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfrtp_2 _27312_ (.D(_00010_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_4 _27313_ (.D(_00011_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_4 _27314_ (.D(_00012_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_4 _27315_ (.D(_00013_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfstp_1 _27316_ (.D(_00014_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .SET_B(net463),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_regs_0_core_clock (.A(clk_i),
    .X(delaynet_0_core_clock));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_30 ();
 sky130_fd_sc_hd__buf_4 _27319_ (.A(net471),
    .X(alert_minor_o));
 sky130_fd_sc_hd__buf_4 _27320_ (.A(net472),
    .X(data_addr_o[0]));
 sky130_fd_sc_hd__buf_4 _27321_ (.A(net473),
    .X(data_addr_o[1]));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__buf_4 _27352_ (.A(net474),
    .X(instr_addr_o[0]));
 sky130_fd_sc_hd__buf_4 _27353_ (.A(net475),
    .X(instr_addr_o[1]));
 sky130_fd_sc_hd__dfrtp_1 \core_busy_q$_DFF_PN0_  (.D(core_busy_d),
    .Q(core_busy_q),
    .RESET_B(net455),
    .CLK(clknet_leaf_21_clk_i_regs));
 sky130_fd_sc_hd__dlxtn_1 \core_clock_gate_i.en_latch$_DLATCH_N_  (.D(_00006_),
    .Q(\core_clock_gate_i.en_latch ),
    .GATE_N(clknet_leaf_21_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcountinhibit_q[0]$_DFFE_PN0P_  (.D(_00015_),
    .Q(\cs_registers_i.mcountinhibit[0] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcountinhibit_q[2]$_DFFE_PN0P_  (.D(_00016_),
    .Q(\cs_registers_i.mcountinhibit[2] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_q[0]$_DFFE_PN0P_  (.D(_00017_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[0] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[10]$_DFFE_PN0P_  (.D(_00018_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[10] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[11]$_DFFE_PN0P_  (.D(_00019_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[11] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[12]$_DFFE_PN0P_  (.D(_00020_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[12] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[13]$_DFFE_PN0P_  (.D(_00021_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[13] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[14]$_DFFE_PN0P_  (.D(_00022_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[14] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[15]$_DFFE_PN0P_  (.D(_00023_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[15] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[16]$_DFFE_PN0P_  (.D(_00024_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[16] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[17]$_DFFE_PN0P_  (.D(_00025_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[17] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[18]$_DFFE_PN0P_  (.D(_00026_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[18] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[19]$_DFFE_PN0P_  (.D(_00027_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[19] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[1]$_DFFE_PN0P_  (.D(_00028_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[1] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[20]$_DFFE_PN0P_  (.D(_00029_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[20] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[21]$_DFFE_PN0P_  (.D(_00030_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[21] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_q[22]$_DFFE_PN0P_  (.D(_00031_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[22] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[23]$_DFFE_PN0P_  (.D(_00032_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[23] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_q[24]$_DFFE_PN0P_  (.D(_00033_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[24] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[25]$_DFFE_PN0P_  (.D(_00034_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[25] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[26]$_DFFE_PN0P_  (.D(_00035_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[26] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_q[27]$_DFFE_PN0P_  (.D(_00036_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[27] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[28]$_DFFE_PN0P_  (.D(_00037_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[28] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[29]$_DFFE_PN0P_  (.D(_00038_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[29] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.mcycle_counter_i.counter_q[2]$_DFFE_PN0P_  (.D(_00039_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[2] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[30]$_DFFE_PN0P_  (.D(_00040_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[30] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[31]$_DFFE_PN0P_  (.D(_00041_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[31] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[32]$_DFFE_PN0P_  (.D(_00042_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[32] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[33]$_DFFE_PN0P_  (.D(_00043_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[33] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[34]$_DFFE_PN0P_  (.D(_00044_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[34] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[35]$_DFFE_PN0P_  (.D(_00045_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[35] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[36]$_DFFE_PN0P_  (.D(_00046_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[36] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[37]$_DFFE_PN0P_  (.D(_00047_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[37] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[38]$_DFFE_PN0P_  (.D(_00048_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[38] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[39]$_DFFE_PN0P_  (.D(_00049_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[39] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[3]$_DFFE_PN0P_  (.D(_00050_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[3] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[40]$_DFFE_PN0P_  (.D(_00051_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[40] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[41]$_DFFE_PN0P_  (.D(_00052_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[41] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[42]$_DFFE_PN0P_  (.D(_00053_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[42] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[43]$_DFFE_PN0P_  (.D(_00054_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[43] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[44]$_DFFE_PN0P_  (.D(_00055_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[44] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[45]$_DFFE_PN0P_  (.D(_00056_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[45] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[46]$_DFFE_PN0P_  (.D(_00057_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[46] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[47]$_DFFE_PN0P_  (.D(_00058_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[47] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[48]$_DFFE_PN0P_  (.D(_00059_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[48] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[49]$_DFFE_PN0P_  (.D(_00060_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[49] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[4]$_DFFE_PN0P_  (.D(_00061_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[4] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[50]$_DFFE_PN0P_  (.D(_00062_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[50] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[51]$_DFFE_PN0P_  (.D(_00063_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[51] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[52]$_DFFE_PN0P_  (.D(_00064_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[52] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[53]$_DFFE_PN0P_  (.D(_00065_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[53] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[54]$_DFFE_PN0P_  (.D(_00066_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[54] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[55]$_DFFE_PN0P_  (.D(_00067_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[55] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[56]$_DFFE_PN0P_  (.D(_00068_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[56] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.mcycle_counter_i.counter_q[57]$_DFFE_PN0P_  (.D(_00069_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[57] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[58]$_DFFE_PN0P_  (.D(_00070_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[58] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[59]$_DFFE_PN0P_  (.D(_00071_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[59] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[5]$_DFFE_PN0P_  (.D(_00072_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[5] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[60]$_DFFE_PN0P_  (.D(_00073_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[60] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[61]$_DFFE_PN0P_  (.D(_00074_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[61] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[62]$_DFFE_PN0P_  (.D(_00075_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[62] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[63]$_DFFE_PN0P_  (.D(_00076_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[63] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[6]$_DFFE_PN0P_  (.D(_00077_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[6] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[7]$_DFFE_PN0P_  (.D(_00078_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[7] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[8]$_DFFE_PN0P_  (.D(_00079_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[8] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.mcycle_counter_i.counter_q[9]$_DFFE_PN0P_  (.D(_00080_),
    .Q(\cs_registers_i.mcycle_counter_i.counter[9] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[0]$_DFFE_PN0P_  (.D(_00081_),
    .Q(\cs_registers_i.mhpmcounter[2][0] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[10]$_DFFE_PN0P_  (.D(_00082_),
    .Q(\cs_registers_i.mhpmcounter[2][10] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[11]$_DFFE_PN0P_  (.D(_00083_),
    .Q(\cs_registers_i.mhpmcounter[2][11] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[12]$_DFFE_PN0P_  (.D(_00084_),
    .Q(\cs_registers_i.mhpmcounter[2][12] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.minstret_counter_i.counter_q[13]$_DFFE_PN0P_  (.D(_00085_),
    .Q(\cs_registers_i.mhpmcounter[2][13] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[14]$_DFFE_PN0P_  (.D(_00086_),
    .Q(\cs_registers_i.mhpmcounter[2][14] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[15]$_DFFE_PN0P_  (.D(_00087_),
    .Q(\cs_registers_i.mhpmcounter[2][15] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[16]$_DFFE_PN0P_  (.D(_00088_),
    .Q(\cs_registers_i.mhpmcounter[2][16] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[17]$_DFFE_PN0P_  (.D(_00089_),
    .Q(\cs_registers_i.mhpmcounter[2][17] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[18]$_DFFE_PN0P_  (.D(_00090_),
    .Q(\cs_registers_i.mhpmcounter[2][18] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[19]$_DFFE_PN0P_  (.D(_00091_),
    .Q(\cs_registers_i.mhpmcounter[2][19] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[1]$_DFFE_PN0P_  (.D(_00092_),
    .Q(\cs_registers_i.mhpmcounter[2][1] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[20]$_DFFE_PN0P_  (.D(_00093_),
    .Q(\cs_registers_i.mhpmcounter[2][20] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[21]$_DFFE_PN0P_  (.D(_00094_),
    .Q(\cs_registers_i.mhpmcounter[2][21] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[22]$_DFFE_PN0P_  (.D(_00095_),
    .Q(\cs_registers_i.mhpmcounter[2][22] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[23]$_DFFE_PN0P_  (.D(_00096_),
    .Q(\cs_registers_i.mhpmcounter[2][23] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.minstret_counter_i.counter_q[24]$_DFFE_PN0P_  (.D(_00097_),
    .Q(\cs_registers_i.mhpmcounter[2][24] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.minstret_counter_i.counter_q[25]$_DFFE_PN0P_  (.D(_00098_),
    .Q(\cs_registers_i.mhpmcounter[2][25] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[26]$_DFFE_PN0P_  (.D(_00099_),
    .Q(\cs_registers_i.mhpmcounter[2][26] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[27]$_DFFE_PN0P_  (.D(_00100_),
    .Q(\cs_registers_i.mhpmcounter[2][27] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[28]$_DFFE_PN0P_  (.D(_00101_),
    .Q(\cs_registers_i.mhpmcounter[2][28] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[29]$_DFFE_PN0P_  (.D(_00102_),
    .Q(\cs_registers_i.mhpmcounter[2][29] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[2]$_DFFE_PN0P_  (.D(_00103_),
    .Q(\cs_registers_i.mhpmcounter[2][2] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[30]$_DFFE_PN0P_  (.D(_00104_),
    .Q(\cs_registers_i.mhpmcounter[2][30] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[31]$_DFFE_PN0P_  (.D(_00105_),
    .Q(\cs_registers_i.mhpmcounter[2][31] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[32]$_DFFE_PN0P_  (.D(_00106_),
    .Q(\cs_registers_i.mhpmcounter[2][32] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[33]$_DFFE_PN0P_  (.D(_00107_),
    .Q(\cs_registers_i.mhpmcounter[2][33] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.minstret_counter_i.counter_q[34]$_DFFE_PN0P_  (.D(_00108_),
    .Q(\cs_registers_i.mhpmcounter[2][34] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[35]$_DFFE_PN0P_  (.D(_00109_),
    .Q(\cs_registers_i.mhpmcounter[2][35] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[36]$_DFFE_PN0P_  (.D(_00110_),
    .Q(\cs_registers_i.mhpmcounter[2][36] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[37]$_DFFE_PN0P_  (.D(_00111_),
    .Q(\cs_registers_i.mhpmcounter[2][37] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[38]$_DFFE_PN0P_  (.D(_00112_),
    .Q(\cs_registers_i.mhpmcounter[2][38] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.minstret_counter_i.counter_q[39]$_DFFE_PN0P_  (.D(_00113_),
    .Q(\cs_registers_i.mhpmcounter[2][39] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[3]$_DFFE_PN0P_  (.D(_00114_),
    .Q(\cs_registers_i.mhpmcounter[2][3] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.minstret_counter_i.counter_q[40]$_DFFE_PN0P_  (.D(_00115_),
    .Q(\cs_registers_i.mhpmcounter[2][40] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[41]$_DFFE_PN0P_  (.D(_00116_),
    .Q(\cs_registers_i.mhpmcounter[2][41] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[42]$_DFFE_PN0P_  (.D(_00117_),
    .Q(\cs_registers_i.mhpmcounter[2][42] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[43]$_DFFE_PN0P_  (.D(_00118_),
    .Q(\cs_registers_i.mhpmcounter[2][43] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.minstret_counter_i.counter_q[44]$_DFFE_PN0P_  (.D(_00119_),
    .Q(\cs_registers_i.mhpmcounter[2][44] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[45]$_DFFE_PN0P_  (.D(_00120_),
    .Q(\cs_registers_i.mhpmcounter[2][45] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.minstret_counter_i.counter_q[46]$_DFFE_PN0P_  (.D(_00121_),
    .Q(\cs_registers_i.mhpmcounter[2][46] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[47]$_DFFE_PN0P_  (.D(_00122_),
    .Q(\cs_registers_i.mhpmcounter[2][47] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[48]$_DFFE_PN0P_  (.D(_00123_),
    .Q(\cs_registers_i.mhpmcounter[2][48] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.minstret_counter_i.counter_q[49]$_DFFE_PN0P_  (.D(_00124_),
    .Q(\cs_registers_i.mhpmcounter[2][49] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.minstret_counter_i.counter_q[4]$_DFFE_PN0P_  (.D(_00125_),
    .Q(\cs_registers_i.mhpmcounter[2][4] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[50]$_DFFE_PN0P_  (.D(_00126_),
    .Q(\cs_registers_i.mhpmcounter[2][50] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[51]$_DFFE_PN0P_  (.D(_00127_),
    .Q(\cs_registers_i.mhpmcounter[2][51] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[52]$_DFFE_PN0P_  (.D(_00128_),
    .Q(\cs_registers_i.mhpmcounter[2][52] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[53]$_DFFE_PN0P_  (.D(_00129_),
    .Q(\cs_registers_i.mhpmcounter[2][53] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[54]$_DFFE_PN0P_  (.D(_00130_),
    .Q(\cs_registers_i.mhpmcounter[2][54] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[55]$_DFFE_PN0P_  (.D(_00131_),
    .Q(\cs_registers_i.mhpmcounter[2][55] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.minstret_counter_i.counter_q[56]$_DFFE_PN0P_  (.D(_00132_),
    .Q(\cs_registers_i.mhpmcounter[2][56] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[57]$_DFFE_PN0P_  (.D(_00133_),
    .Q(\cs_registers_i.mhpmcounter[2][57] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[58]$_DFFE_PN0P_  (.D(_00134_),
    .Q(\cs_registers_i.mhpmcounter[2][58] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[59]$_DFFE_PN0P_  (.D(_00135_),
    .Q(\cs_registers_i.mhpmcounter[2][59] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[5]$_DFFE_PN0P_  (.D(_00136_),
    .Q(\cs_registers_i.mhpmcounter[2][5] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[60]$_DFFE_PN0P_  (.D(_00137_),
    .Q(\cs_registers_i.mhpmcounter[2][60] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[61]$_DFFE_PN0P_  (.D(_00138_),
    .Q(\cs_registers_i.mhpmcounter[2][61] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[62]$_DFFE_PN0P_  (.D(_00139_),
    .Q(\cs_registers_i.mhpmcounter[2][62] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[63]$_DFFE_PN0P_  (.D(_00140_),
    .Q(\cs_registers_i.mhpmcounter[2][63] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[6]$_DFFE_PN0P_  (.D(_00141_),
    .Q(\cs_registers_i.mhpmcounter[2][6] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[7]$_DFFE_PN0P_  (.D(_00142_),
    .Q(\cs_registers_i.mhpmcounter[2][7] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[8]$_DFFE_PN0P_  (.D(_00143_),
    .Q(\cs_registers_i.mhpmcounter[2][8] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.minstret_counter_i.counter_q[9]$_DFFE_PN0P_  (.D(_00144_),
    .Q(\cs_registers_i.mhpmcounter[2][9] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfstp_2 \cs_registers_i.priv_lvl_q[0]$_DFFE_PN1P_  (.D(_00145_),
    .Q(\cs_registers_i.priv_lvl_q[0] ),
    .SET_B(net454),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfstp_1 \cs_registers_i.priv_lvl_q[1]$_DFFE_PN1P_  (.D(_00146_),
    .Q(\cs_registers_i.priv_lvl_q[1] ),
    .SET_B(net454),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfstp_1 \cs_registers_i.u_dcsr_csr.rdata_q[0]$_DFFE_PN1P_  (.D(_00147_),
    .Q(\cs_registers_i.dcsr_q[0] ),
    .SET_B(net454),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dcsr_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_00148_),
    .Q(\cs_registers_i.dcsr_q[11] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_dcsr_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_00149_),
    .Q(\cs_registers_i.dcsr_q[12] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dcsr_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_00150_),
    .Q(\cs_registers_i.dcsr_q[13] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_dcsr_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_00151_),
    .Q(\cs_registers_i.dcsr_q[15] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfstp_1 \cs_registers_i.u_dcsr_csr.rdata_q[1]$_DFFE_PN1P_  (.D(_00152_),
    .Q(\cs_registers_i.dcsr_q[1] ),
    .SET_B(net454),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.u_dcsr_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_00153_),
    .Q(\cs_registers_i.dcsr_q[2] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dcsr_csr.rdata_q[6]$_DFFE_PN0P_  (.D(_00154_),
    .Q(\cs_registers_i.dcsr_q[6] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dcsr_csr.rdata_q[7]$_DFFE_PN0P_  (.D(_00155_),
    .Q(\cs_registers_i.dcsr_q[7] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dcsr_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_00156_),
    .Q(\cs_registers_i.dcsr_q[8] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[10]$_DFFE_PN0P_  (.D(_00157_),
    .Q(\cs_registers_i.csr_depc_o[10] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_00158_),
    .Q(\cs_registers_i.csr_depc_o[11] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_00159_),
    .Q(\cs_registers_i.csr_depc_o[12] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_00160_),
    .Q(\cs_registers_i.csr_depc_o[13] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.u_depc_csr.rdata_q[14]$_DFFE_PN0P_  (.D(_00161_),
    .Q(\cs_registers_i.csr_depc_o[14] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_00162_),
    .Q(\cs_registers_i.csr_depc_o[15] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[16]$_DFFE_PN0P_  (.D(_00163_),
    .Q(\cs_registers_i.csr_depc_o[16] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[17]$_DFFE_PN0P_  (.D(_00164_),
    .Q(\cs_registers_i.csr_depc_o[17] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[18]$_DFFE_PN0P_  (.D(_00165_),
    .Q(\cs_registers_i.csr_depc_o[18] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[19]$_DFFE_PN0P_  (.D(_00166_),
    .Q(\cs_registers_i.csr_depc_o[19] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.u_depc_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_00167_),
    .Q(\cs_registers_i.csr_depc_o[1] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[20]$_DFFE_PN0P_  (.D(_00168_),
    .Q(\cs_registers_i.csr_depc_o[20] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[21]$_DFFE_PN0P_  (.D(_00169_),
    .Q(\cs_registers_i.csr_depc_o[21] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[22]$_DFFE_PN0P_  (.D(_00170_),
    .Q(\cs_registers_i.csr_depc_o[22] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[23]$_DFFE_PN0P_  (.D(_00171_),
    .Q(\cs_registers_i.csr_depc_o[23] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[24]$_DFFE_PN0P_  (.D(_00172_),
    .Q(\cs_registers_i.csr_depc_o[24] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[25]$_DFFE_PN0P_  (.D(_00173_),
    .Q(\cs_registers_i.csr_depc_o[25] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[26]$_DFFE_PN0P_  (.D(_00174_),
    .Q(\cs_registers_i.csr_depc_o[26] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[27]$_DFFE_PN0P_  (.D(_00175_),
    .Q(\cs_registers_i.csr_depc_o[27] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[28]$_DFFE_PN0P_  (.D(_00176_),
    .Q(\cs_registers_i.csr_depc_o[28] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[29]$_DFFE_PN0P_  (.D(_00177_),
    .Q(\cs_registers_i.csr_depc_o[29] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_00178_),
    .Q(\cs_registers_i.csr_depc_o[2] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[30]$_DFFE_PN0P_  (.D(_00179_),
    .Q(\cs_registers_i.csr_depc_o[30] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[31]$_DFFE_PN0P_  (.D(_00180_),
    .Q(\cs_registers_i.csr_depc_o[31] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_00181_),
    .Q(\cs_registers_i.csr_depc_o[3] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_depc_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_00182_),
    .Q(\cs_registers_i.csr_depc_o[4] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_00183_),
    .Q(\cs_registers_i.csr_depc_o[5] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[6]$_DFFE_PN0P_  (.D(_00184_),
    .Q(\cs_registers_i.csr_depc_o[6] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[7]$_DFFE_PN0P_  (.D(_00185_),
    .Q(\cs_registers_i.csr_depc_o[7] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_00186_),
    .Q(\cs_registers_i.csr_depc_o[8] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_depc_csr.rdata_q[9]$_DFFE_PN0P_  (.D(_00187_),
    .Q(\cs_registers_i.csr_depc_o[9] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_00188_),
    .Q(\cs_registers_i.dscratch0_q[0] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[10]$_DFFE_PN0P_  (.D(_00189_),
    .Q(\cs_registers_i.dscratch0_q[10] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_00190_),
    .Q(\cs_registers_i.dscratch0_q[11] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_00191_),
    .Q(\cs_registers_i.dscratch0_q[12] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_00192_),
    .Q(\cs_registers_i.dscratch0_q[13] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[14]$_DFFE_PN0P_  (.D(_00193_),
    .Q(\cs_registers_i.dscratch0_q[14] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_00194_),
    .Q(\cs_registers_i.dscratch0_q[15] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[16]$_DFFE_PN0P_  (.D(_00195_),
    .Q(\cs_registers_i.dscratch0_q[16] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[17]$_DFFE_PN0P_  (.D(_00196_),
    .Q(\cs_registers_i.dscratch0_q[17] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[18]$_DFFE_PN0P_  (.D(_00197_),
    .Q(\cs_registers_i.dscratch0_q[18] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[19]$_DFFE_PN0P_  (.D(_00198_),
    .Q(\cs_registers_i.dscratch0_q[19] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_00199_),
    .Q(\cs_registers_i.dscratch0_q[1] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[20]$_DFFE_PN0P_  (.D(_00200_),
    .Q(\cs_registers_i.dscratch0_q[20] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[21]$_DFFE_PN0P_  (.D(_00201_),
    .Q(\cs_registers_i.dscratch0_q[21] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[22]$_DFFE_PN0P_  (.D(_00202_),
    .Q(\cs_registers_i.dscratch0_q[22] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[23]$_DFFE_PN0P_  (.D(_00203_),
    .Q(\cs_registers_i.dscratch0_q[23] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[24]$_DFFE_PN0P_  (.D(_00204_),
    .Q(\cs_registers_i.dscratch0_q[24] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[25]$_DFFE_PN0P_  (.D(_00205_),
    .Q(\cs_registers_i.dscratch0_q[25] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[26]$_DFFE_PN0P_  (.D(_00206_),
    .Q(\cs_registers_i.dscratch0_q[26] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[27]$_DFFE_PN0P_  (.D(_00207_),
    .Q(\cs_registers_i.dscratch0_q[27] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[28]$_DFFE_PN0P_  (.D(_00208_),
    .Q(\cs_registers_i.dscratch0_q[28] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[29]$_DFFE_PN0P_  (.D(_00209_),
    .Q(\cs_registers_i.dscratch0_q[29] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_00210_),
    .Q(\cs_registers_i.dscratch0_q[2] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[30]$_DFFE_PN0P_  (.D(_00211_),
    .Q(\cs_registers_i.dscratch0_q[30] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[31]$_DFFE_PN0P_  (.D(_00212_),
    .Q(\cs_registers_i.dscratch0_q[31] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_00213_),
    .Q(\cs_registers_i.dscratch0_q[3] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_00214_),
    .Q(\cs_registers_i.dscratch0_q[4] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_00215_),
    .Q(\cs_registers_i.dscratch0_q[5] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[6]$_DFFE_PN0P_  (.D(_00216_),
    .Q(\cs_registers_i.dscratch0_q[6] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[7]$_DFFE_PN0P_  (.D(_00217_),
    .Q(\cs_registers_i.dscratch0_q[7] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_00218_),
    .Q(\cs_registers_i.dscratch0_q[8] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch0_csr.rdata_q[9]$_DFFE_PN0P_  (.D(_00219_),
    .Q(\cs_registers_i.dscratch0_q[9] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_00220_),
    .Q(\cs_registers_i.dscratch1_q[0] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[10]$_DFFE_PN0P_  (.D(_00221_),
    .Q(\cs_registers_i.dscratch1_q[10] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_00222_),
    .Q(\cs_registers_i.dscratch1_q[11] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_00223_),
    .Q(\cs_registers_i.dscratch1_q[12] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_00224_),
    .Q(\cs_registers_i.dscratch1_q[13] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[14]$_DFFE_PN0P_  (.D(_00225_),
    .Q(\cs_registers_i.dscratch1_q[14] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_00226_),
    .Q(\cs_registers_i.dscratch1_q[15] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[16]$_DFFE_PN0P_  (.D(_00227_),
    .Q(\cs_registers_i.dscratch1_q[16] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[17]$_DFFE_PN0P_  (.D(_00228_),
    .Q(\cs_registers_i.dscratch1_q[17] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[18]$_DFFE_PN0P_  (.D(_00229_),
    .Q(\cs_registers_i.dscratch1_q[18] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[19]$_DFFE_PN0P_  (.D(_00230_),
    .Q(\cs_registers_i.dscratch1_q[19] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_00231_),
    .Q(\cs_registers_i.dscratch1_q[1] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[20]$_DFFE_PN0P_  (.D(_00232_),
    .Q(\cs_registers_i.dscratch1_q[20] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[21]$_DFFE_PN0P_  (.D(_00233_),
    .Q(\cs_registers_i.dscratch1_q[21] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[22]$_DFFE_PN0P_  (.D(_00234_),
    .Q(\cs_registers_i.dscratch1_q[22] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[23]$_DFFE_PN0P_  (.D(_00235_),
    .Q(\cs_registers_i.dscratch1_q[23] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[24]$_DFFE_PN0P_  (.D(_00236_),
    .Q(\cs_registers_i.dscratch1_q[24] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[25]$_DFFE_PN0P_  (.D(_00237_),
    .Q(\cs_registers_i.dscratch1_q[25] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[26]$_DFFE_PN0P_  (.D(_00238_),
    .Q(\cs_registers_i.dscratch1_q[26] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[27]$_DFFE_PN0P_  (.D(_00239_),
    .Q(\cs_registers_i.dscratch1_q[27] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[28]$_DFFE_PN0P_  (.D(_00240_),
    .Q(\cs_registers_i.dscratch1_q[28] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[29]$_DFFE_PN0P_  (.D(_00241_),
    .Q(\cs_registers_i.dscratch1_q[29] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_00242_),
    .Q(\cs_registers_i.dscratch1_q[2] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[30]$_DFFE_PN0P_  (.D(_00243_),
    .Q(\cs_registers_i.dscratch1_q[30] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[31]$_DFFE_PN0P_  (.D(_00244_),
    .Q(\cs_registers_i.dscratch1_q[31] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_00245_),
    .Q(\cs_registers_i.dscratch1_q[3] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_00246_),
    .Q(\cs_registers_i.dscratch1_q[4] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_00247_),
    .Q(\cs_registers_i.dscratch1_q[5] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[6]$_DFFE_PN0P_  (.D(_00248_),
    .Q(\cs_registers_i.dscratch1_q[6] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[7]$_DFFE_PN0P_  (.D(_00249_),
    .Q(\cs_registers_i.dscratch1_q[7] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_00250_),
    .Q(\cs_registers_i.dscratch1_q[8] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_dscratch1_csr.rdata_q[9]$_DFFE_PN0P_  (.D(_00251_),
    .Q(\cs_registers_i.dscratch1_q[9] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mcause_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_00252_),
    .Q(\cs_registers_i.mcause_q[0] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mcause_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_00253_),
    .Q(\cs_registers_i.mcause_q[1] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mcause_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_00254_),
    .Q(\cs_registers_i.mcause_q[2] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mcause_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_00255_),
    .Q(\cs_registers_i.mcause_q[3] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mcause_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_00256_),
    .Q(\cs_registers_i.mcause_q[4] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mcause_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_00257_),
    .Q(\cs_registers_i.mcause_q[5] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mepc_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_00258_),
    .Q(\cs_registers_i.csr_mepc_o[0] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mepc_csr.rdata_q[10]$_DFFE_PN0P_  (.D(_00259_),
    .Q(\cs_registers_i.csr_mepc_o[10] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mepc_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_00260_),
    .Q(\cs_registers_i.csr_mepc_o[11] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.u_mepc_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_00261_),
    .Q(\cs_registers_i.csr_mepc_o[12] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mepc_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_00262_),
    .Q(\cs_registers_i.csr_mepc_o[13] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mepc_csr.rdata_q[14]$_DFFE_PN0P_  (.D(_00263_),
    .Q(\cs_registers_i.csr_mepc_o[14] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mepc_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_00264_),
    .Q(\cs_registers_i.csr_mepc_o[15] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mepc_csr.rdata_q[16]$_DFFE_PN0P_  (.D(_00265_),
    .Q(\cs_registers_i.csr_mepc_o[16] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mepc_csr.rdata_q[17]$_DFFE_PN0P_  (.D(_00266_),
    .Q(\cs_registers_i.csr_mepc_o[17] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.u_mepc_csr.rdata_q[18]$_DFFE_PN0P_  (.D(_00267_),
    .Q(\cs_registers_i.csr_mepc_o[18] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.u_mepc_csr.rdata_q[19]$_DFFE_PN0P_  (.D(_00268_),
    .Q(\cs_registers_i.csr_mepc_o[19] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.u_mepc_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_00269_),
    .Q(\cs_registers_i.csr_mepc_o[1] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mepc_csr.rdata_q[20]$_DFFE_PN0P_  (.D(_00270_),
    .Q(\cs_registers_i.csr_mepc_o[20] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mepc_csr.rdata_q[21]$_DFFE_PN0P_  (.D(_00271_),
    .Q(\cs_registers_i.csr_mepc_o[21] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.u_mepc_csr.rdata_q[22]$_DFFE_PN0P_  (.D(_00272_),
    .Q(\cs_registers_i.csr_mepc_o[22] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.u_mepc_csr.rdata_q[23]$_DFFE_PN0P_  (.D(_00273_),
    .Q(\cs_registers_i.csr_mepc_o[23] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mepc_csr.rdata_q[24]$_DFFE_PN0P_  (.D(_00274_),
    .Q(\cs_registers_i.csr_mepc_o[24] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mepc_csr.rdata_q[25]$_DFFE_PN0P_  (.D(_00275_),
    .Q(\cs_registers_i.csr_mepc_o[25] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mepc_csr.rdata_q[26]$_DFFE_PN0P_  (.D(_00276_),
    .Q(\cs_registers_i.csr_mepc_o[26] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mepc_csr.rdata_q[27]$_DFFE_PN0P_  (.D(_00277_),
    .Q(\cs_registers_i.csr_mepc_o[27] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mepc_csr.rdata_q[28]$_DFFE_PN0P_  (.D(_00278_),
    .Q(\cs_registers_i.csr_mepc_o[28] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mepc_csr.rdata_q[29]$_DFFE_PN0P_  (.D(_00279_),
    .Q(\cs_registers_i.csr_mepc_o[29] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mepc_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_00280_),
    .Q(\cs_registers_i.csr_mepc_o[2] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mepc_csr.rdata_q[30]$_DFFE_PN0P_  (.D(_00281_),
    .Q(\cs_registers_i.csr_mepc_o[30] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mepc_csr.rdata_q[31]$_DFFE_PN0P_  (.D(_00282_),
    .Q(\cs_registers_i.csr_mepc_o[31] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mepc_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_00283_),
    .Q(\cs_registers_i.csr_mepc_o[3] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mepc_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_00284_),
    .Q(\cs_registers_i.csr_mepc_o[4] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mepc_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_00285_),
    .Q(\cs_registers_i.csr_mepc_o[5] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mepc_csr.rdata_q[6]$_DFFE_PN0P_  (.D(_00286_),
    .Q(\cs_registers_i.csr_mepc_o[6] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.u_mepc_csr.rdata_q[7]$_DFFE_PN0P_  (.D(_00287_),
    .Q(\cs_registers_i.csr_mepc_o[7] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mepc_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_00288_),
    .Q(\cs_registers_i.csr_mepc_o[8] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mepc_csr.rdata_q[9]$_DFFE_PN0P_  (.D(_00289_),
    .Q(\cs_registers_i.csr_mepc_o[9] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mie_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_00290_),
    .Q(\cs_registers_i.mie_q[0] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mie_csr.rdata_q[10]$_DFFE_PN0P_  (.D(_00291_),
    .Q(\cs_registers_i.mie_q[10] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mie_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_00292_),
    .Q(\cs_registers_i.mie_q[11] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mie_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_00293_),
    .Q(\cs_registers_i.mie_q[12] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mie_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_00294_),
    .Q(\cs_registers_i.mie_q[13] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mie_csr.rdata_q[14]$_DFFE_PN0P_  (.D(_00295_),
    .Q(\cs_registers_i.mie_q[14] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mie_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_00296_),
    .Q(\cs_registers_i.mie_q[15] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mie_csr.rdata_q[16]$_DFFE_PN0P_  (.D(_00297_),
    .Q(\cs_registers_i.mie_q[16] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mie_csr.rdata_q[17]$_DFFE_PN0P_  (.D(_00298_),
    .Q(\cs_registers_i.mie_q[17] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mie_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_00299_),
    .Q(\cs_registers_i.mie_q[1] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.u_mie_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_00300_),
    .Q(\cs_registers_i.mie_q[2] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.u_mie_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_00301_),
    .Q(\cs_registers_i.mie_q[3] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mie_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_00302_),
    .Q(\cs_registers_i.mie_q[4] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.u_mie_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_00303_),
    .Q(\cs_registers_i.mie_q[5] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mie_csr.rdata_q[6]$_DFFE_PN0P_  (.D(_00304_),
    .Q(\cs_registers_i.mie_q[6] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mie_csr.rdata_q[7]$_DFFE_PN0P_  (.D(_00305_),
    .Q(\cs_registers_i.mie_q[7] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.u_mie_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_00306_),
    .Q(\cs_registers_i.mie_q[8] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mie_csr.rdata_q[9]$_DFFE_PN0P_  (.D(_00307_),
    .Q(\cs_registers_i.mie_q[9] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_00308_),
    .Q(\cs_registers_i.mscratch_q[0] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[10]$_DFFE_PN0P_  (.D(_00309_),
    .Q(\cs_registers_i.mscratch_q[10] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_00310_),
    .Q(\cs_registers_i.mscratch_q[11] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_00311_),
    .Q(\cs_registers_i.mscratch_q[12] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_00312_),
    .Q(\cs_registers_i.mscratch_q[13] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[14]$_DFFE_PN0P_  (.D(_00313_),
    .Q(\cs_registers_i.mscratch_q[14] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_00314_),
    .Q(\cs_registers_i.mscratch_q[15] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[16]$_DFFE_PN0P_  (.D(_00315_),
    .Q(\cs_registers_i.mscratch_q[16] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[17]$_DFFE_PN0P_  (.D(_00316_),
    .Q(\cs_registers_i.mscratch_q[17] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[18]$_DFFE_PN0P_  (.D(_00317_),
    .Q(\cs_registers_i.mscratch_q[18] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[19]$_DFFE_PN0P_  (.D(_00318_),
    .Q(\cs_registers_i.mscratch_q[19] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_00319_),
    .Q(\cs_registers_i.mscratch_q[1] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[20]$_DFFE_PN0P_  (.D(_00320_),
    .Q(\cs_registers_i.mscratch_q[20] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[21]$_DFFE_PN0P_  (.D(_00321_),
    .Q(\cs_registers_i.mscratch_q[21] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[22]$_DFFE_PN0P_  (.D(_00322_),
    .Q(\cs_registers_i.mscratch_q[22] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[23]$_DFFE_PN0P_  (.D(_00323_),
    .Q(\cs_registers_i.mscratch_q[23] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[24]$_DFFE_PN0P_  (.D(_00324_),
    .Q(\cs_registers_i.mscratch_q[24] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[25]$_DFFE_PN0P_  (.D(_00325_),
    .Q(\cs_registers_i.mscratch_q[25] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[26]$_DFFE_PN0P_  (.D(_00326_),
    .Q(\cs_registers_i.mscratch_q[26] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[27]$_DFFE_PN0P_  (.D(_00327_),
    .Q(\cs_registers_i.mscratch_q[27] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[28]$_DFFE_PN0P_  (.D(_00328_),
    .Q(\cs_registers_i.mscratch_q[28] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[29]$_DFFE_PN0P_  (.D(_00329_),
    .Q(\cs_registers_i.mscratch_q[29] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_00330_),
    .Q(\cs_registers_i.mscratch_q[2] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[30]$_DFFE_PN0P_  (.D(_00331_),
    .Q(\cs_registers_i.mscratch_q[30] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[31]$_DFFE_PN0P_  (.D(_00332_),
    .Q(\cs_registers_i.mscratch_q[31] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_00333_),
    .Q(\cs_registers_i.mscratch_q[3] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_00334_),
    .Q(\cs_registers_i.mscratch_q[4] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_00335_),
    .Q(\cs_registers_i.mscratch_q[5] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[6]$_DFFE_PN0P_  (.D(_00336_),
    .Q(\cs_registers_i.mscratch_q[6] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[7]$_DFFE_PN0P_  (.D(_00337_),
    .Q(\cs_registers_i.mscratch_q[7] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_00338_),
    .Q(\cs_registers_i.mscratch_q[8] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mscratch_csr.rdata_q[9]$_DFFE_PN0P_  (.D(_00339_),
    .Q(\cs_registers_i.mscratch_q[9] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_cause_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_00340_),
    .Q(\cs_registers_i.mstack_cause_q[0] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_cause_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_00341_),
    .Q(\cs_registers_i.mstack_cause_q[1] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_cause_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_00342_),
    .Q(\cs_registers_i.mstack_cause_q[2] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_cause_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_00343_),
    .Q(\cs_registers_i.mstack_cause_q[3] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_cause_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_00344_),
    .Q(\cs_registers_i.mstack_cause_q[4] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_cause_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_00345_),
    .Q(\cs_registers_i.mstack_cause_q[5] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_00346_),
    .Q(\cs_registers_i.mstack_q[0] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_00347_),
    .Q(\cs_registers_i.mstack_q[1] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfstp_1 \cs_registers_i.u_mstack_csr.rdata_q[2]$_DFFE_PN1P_  (.D(_00348_),
    .Q(\cs_registers_i.mstack_q[2] ),
    .SET_B(net452),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_00349_),
    .Q(\cs_registers_i.mstack_epc_q[0] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[10]$_DFFE_PN0P_  (.D(_00350_),
    .Q(\cs_registers_i.mstack_epc_q[10] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_00351_),
    .Q(\cs_registers_i.mstack_epc_q[11] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_00352_),
    .Q(\cs_registers_i.mstack_epc_q[12] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_00353_),
    .Q(\cs_registers_i.mstack_epc_q[13] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[14]$_DFFE_PN0P_  (.D(_00354_),
    .Q(\cs_registers_i.mstack_epc_q[14] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_00355_),
    .Q(\cs_registers_i.mstack_epc_q[15] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[16]$_DFFE_PN0P_  (.D(_00356_),
    .Q(\cs_registers_i.mstack_epc_q[16] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[17]$_DFFE_PN0P_  (.D(_00357_),
    .Q(\cs_registers_i.mstack_epc_q[17] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[18]$_DFFE_PN0P_  (.D(_00358_),
    .Q(\cs_registers_i.mstack_epc_q[18] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[19]$_DFFE_PN0P_  (.D(_00359_),
    .Q(\cs_registers_i.mstack_epc_q[19] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_00360_),
    .Q(\cs_registers_i.mstack_epc_q[1] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[20]$_DFFE_PN0P_  (.D(_00361_),
    .Q(\cs_registers_i.mstack_epc_q[20] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[21]$_DFFE_PN0P_  (.D(_00362_),
    .Q(\cs_registers_i.mstack_epc_q[21] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[22]$_DFFE_PN0P_  (.D(_00363_),
    .Q(\cs_registers_i.mstack_epc_q[22] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[23]$_DFFE_PN0P_  (.D(_00364_),
    .Q(\cs_registers_i.mstack_epc_q[23] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[24]$_DFFE_PN0P_  (.D(_00365_),
    .Q(\cs_registers_i.mstack_epc_q[24] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[25]$_DFFE_PN0P_  (.D(_00366_),
    .Q(\cs_registers_i.mstack_epc_q[25] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[26]$_DFFE_PN0P_  (.D(_00367_),
    .Q(\cs_registers_i.mstack_epc_q[26] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[27]$_DFFE_PN0P_  (.D(_00368_),
    .Q(\cs_registers_i.mstack_epc_q[27] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[28]$_DFFE_PN0P_  (.D(_00369_),
    .Q(\cs_registers_i.mstack_epc_q[28] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[29]$_DFFE_PN0P_  (.D(_00370_),
    .Q(\cs_registers_i.mstack_epc_q[29] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_00371_),
    .Q(\cs_registers_i.mstack_epc_q[2] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[30]$_DFFE_PN0P_  (.D(_00372_),
    .Q(\cs_registers_i.mstack_epc_q[30] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[31]$_DFFE_PN0P_  (.D(_00373_),
    .Q(\cs_registers_i.mstack_epc_q[31] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_00374_),
    .Q(\cs_registers_i.mstack_epc_q[3] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_00375_),
    .Q(\cs_registers_i.mstack_epc_q[4] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_00376_),
    .Q(\cs_registers_i.mstack_epc_q[5] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[6]$_DFFE_PN0P_  (.D(_00377_),
    .Q(\cs_registers_i.mstack_epc_q[6] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[7]$_DFFE_PN0P_  (.D(_00378_),
    .Q(\cs_registers_i.mstack_epc_q[7] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_00379_),
    .Q(\cs_registers_i.mstack_epc_q[8] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstack_epc_csr.rdata_q[9]$_DFFE_PN0P_  (.D(_00380_),
    .Q(\cs_registers_i.mstack_epc_q[9] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mstatus_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_00381_),
    .Q(\cs_registers_i.csr_mstatus_tw_o ),
    .RESET_B(net454),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstatus_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_00382_),
    .Q(\cs_registers_i.mstatus_q[1] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mstatus_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_00383_),
    .Q(\cs_registers_i.mstack_d[0] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mstatus_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_00384_),
    .Q(\cs_registers_i.mstack_d[1] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfstp_1 \cs_registers_i.u_mstatus_csr.rdata_q[4]$_DFFE_PN1P_  (.D(_00385_),
    .Q(\cs_registers_i.mstack_d[2] ),
    .SET_B(net452),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.u_mstatus_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_00386_),
    .Q(\cs_registers_i.csr_mstatus_mie_o ),
    .RESET_B(net452),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rdata_q[0]$_DFFE_PN0P_  (.D(_00387_),
    .Q(\cs_registers_i.mtval_q[0] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rdata_q[10]$_DFFE_PN0P_  (.D(_00388_),
    .Q(\cs_registers_i.mtval_q[10] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_00389_),
    .Q(\cs_registers_i.mtval_q[11] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.u_mtval_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_00390_),
    .Q(\cs_registers_i.mtval_q[12] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.u_mtval_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_00391_),
    .Q(\cs_registers_i.mtval_q[13] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.u_mtval_csr.rdata_q[14]$_DFFE_PN0P_  (.D(_00392_),
    .Q(\cs_registers_i.mtval_q[14] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.u_mtval_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_00393_),
    .Q(\cs_registers_i.mtval_q[15] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rdata_q[16]$_DFFE_PN0P_  (.D(_00394_),
    .Q(\cs_registers_i.mtval_q[16] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.u_mtval_csr.rdata_q[17]$_DFFE_PN0P_  (.D(_00395_),
    .Q(\cs_registers_i.mtval_q[17] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rdata_q[18]$_DFFE_PN0P_  (.D(_00396_),
    .Q(\cs_registers_i.mtval_q[18] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rdata_q[19]$_DFFE_PN0P_  (.D(_00397_),
    .Q(\cs_registers_i.mtval_q[19] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rdata_q[1]$_DFFE_PN0P_  (.D(_00398_),
    .Q(\cs_registers_i.mtval_q[1] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rdata_q[20]$_DFFE_PN0P_  (.D(_00399_),
    .Q(\cs_registers_i.mtval_q[20] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rdata_q[21]$_DFFE_PN0P_  (.D(_00400_),
    .Q(\cs_registers_i.mtval_q[21] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rdata_q[22]$_DFFE_PN0P_  (.D(_00401_),
    .Q(\cs_registers_i.mtval_q[22] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rdata_q[23]$_DFFE_PN0P_  (.D(_00402_),
    .Q(\cs_registers_i.mtval_q[23] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rdata_q[24]$_DFFE_PN0P_  (.D(_00403_),
    .Q(\cs_registers_i.mtval_q[24] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rdata_q[25]$_DFFE_PN0P_  (.D(_00404_),
    .Q(\cs_registers_i.mtval_q[25] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rdata_q[26]$_DFFE_PN0P_  (.D(_00405_),
    .Q(\cs_registers_i.mtval_q[26] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rdata_q[27]$_DFFE_PN0P_  (.D(_00406_),
    .Q(\cs_registers_i.mtval_q[27] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rdata_q[28]$_DFFE_PN0P_  (.D(_00407_),
    .Q(\cs_registers_i.mtval_q[28] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rdata_q[29]$_DFFE_PN0P_  (.D(_00408_),
    .Q(\cs_registers_i.mtval_q[29] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rdata_q[2]$_DFFE_PN0P_  (.D(_00409_),
    .Q(\cs_registers_i.mtval_q[2] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rdata_q[30]$_DFFE_PN0P_  (.D(_00410_),
    .Q(\cs_registers_i.mtval_q[30] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rdata_q[31]$_DFFE_PN0P_  (.D(_00411_),
    .Q(\cs_registers_i.mtval_q[31] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rdata_q[3]$_DFFE_PN0P_  (.D(_00412_),
    .Q(\cs_registers_i.mtval_q[3] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rdata_q[4]$_DFFE_PN0P_  (.D(_00413_),
    .Q(\cs_registers_i.mtval_q[4] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rdata_q[5]$_DFFE_PN0P_  (.D(_00414_),
    .Q(\cs_registers_i.mtval_q[5] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rdata_q[6]$_DFFE_PN0P_  (.D(_00415_),
    .Q(\cs_registers_i.mtval_q[6] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.u_mtval_csr.rdata_q[7]$_DFFE_PN0P_  (.D(_00416_),
    .Q(\cs_registers_i.mtval_q[7] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_00417_),
    .Q(\cs_registers_i.mtval_q[8] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtval_csr.rdata_q[9]$_DFFE_PN0P_  (.D(_00418_),
    .Q(\cs_registers_i.mtval_q[9] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtvec_csr.rdata_q[10]$_DFFE_PN0P_  (.D(_00419_),
    .Q(\cs_registers_i.csr_mtvec_o[10] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtvec_csr.rdata_q[11]$_DFFE_PN0P_  (.D(_00420_),
    .Q(\cs_registers_i.csr_mtvec_o[11] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtvec_csr.rdata_q[12]$_DFFE_PN0P_  (.D(_00421_),
    .Q(\cs_registers_i.csr_mtvec_o[12] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtvec_csr.rdata_q[13]$_DFFE_PN0P_  (.D(_00422_),
    .Q(\cs_registers_i.csr_mtvec_o[13] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtvec_csr.rdata_q[14]$_DFFE_PN0P_  (.D(_00423_),
    .Q(\cs_registers_i.csr_mtvec_o[14] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtvec_csr.rdata_q[15]$_DFFE_PN0P_  (.D(_00424_),
    .Q(\cs_registers_i.csr_mtvec_o[15] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtvec_csr.rdata_q[16]$_DFFE_PN0P_  (.D(_00425_),
    .Q(\cs_registers_i.csr_mtvec_o[16] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtvec_csr.rdata_q[17]$_DFFE_PN0P_  (.D(_00426_),
    .Q(\cs_registers_i.csr_mtvec_o[17] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtvec_csr.rdata_q[18]$_DFFE_PN0P_  (.D(_00427_),
    .Q(\cs_registers_i.csr_mtvec_o[18] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtvec_csr.rdata_q[19]$_DFFE_PN0P_  (.D(_00428_),
    .Q(\cs_registers_i.csr_mtvec_o[19] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtvec_csr.rdata_q[20]$_DFFE_PN0P_  (.D(_00429_),
    .Q(\cs_registers_i.csr_mtvec_o[20] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtvec_csr.rdata_q[21]$_DFFE_PN0P_  (.D(_00430_),
    .Q(\cs_registers_i.csr_mtvec_o[21] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtvec_csr.rdata_q[22]$_DFFE_PN0P_  (.D(_00431_),
    .Q(\cs_registers_i.csr_mtvec_o[22] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtvec_csr.rdata_q[23]$_DFFE_PN0P_  (.D(_00432_),
    .Q(\cs_registers_i.csr_mtvec_o[23] ),
    .RESET_B(net452),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtvec_csr.rdata_q[24]$_DFFE_PN0P_  (.D(_00433_),
    .Q(\cs_registers_i.csr_mtvec_o[24] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtvec_csr.rdata_q[25]$_DFFE_PN0P_  (.D(_00434_),
    .Q(\cs_registers_i.csr_mtvec_o[25] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtvec_csr.rdata_q[26]$_DFFE_PN0P_  (.D(_00435_),
    .Q(\cs_registers_i.csr_mtvec_o[26] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtvec_csr.rdata_q[27]$_DFFE_PN0P_  (.D(_00436_),
    .Q(\cs_registers_i.csr_mtvec_o[27] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtvec_csr.rdata_q[28]$_DFFE_PN0P_  (.D(_00437_),
    .Q(\cs_registers_i.csr_mtvec_o[28] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtvec_csr.rdata_q[29]$_DFFE_PN0P_  (.D(_00438_),
    .Q(\cs_registers_i.csr_mtvec_o[29] ),
    .RESET_B(net453),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtvec_csr.rdata_q[30]$_DFFE_PN0P_  (.D(_00439_),
    .Q(\cs_registers_i.csr_mtvec_o[30] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfrtp_2 \cs_registers_i.u_mtvec_csr.rdata_q[31]$_DFFE_PN0P_  (.D(_00440_),
    .Q(\cs_registers_i.csr_mtvec_o[31] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfrtp_1 \cs_registers_i.u_mtvec_csr.rdata_q[8]$_DFFE_PN0P_  (.D(_00441_),
    .Q(\cs_registers_i.csr_mtvec_o[8] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_4 \cs_registers_i.u_mtvec_csr.rdata_q[9]$_DFFE_PN0P_  (.D(_00442_),
    .Q(\cs_registers_i.csr_mtvec_o[9] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_by_zero_q$_DFFE_PN0P_  (.D(_00443_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_by_zero_q ),
    .RESET_B(net463),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_4 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0]$_DFFE_PN0P_  (.D(_00444_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_4 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1]$_DFFE_PN0P_  (.D(_00445_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_4 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2]$_DFFE_PN0P_  (.D(_00446_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_4 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[3]$_DFFE_PN0P_  (.D(_00447_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_4 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[4]$_DFFE_PN0P_  (.D(_00448_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfstp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0]$_DFF_PN1_  (.D(_00000_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .SET_B(net462),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_4 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3]$_DFF_PN0_  (.D(_00001_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_4 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1]$_DFF_PN0_  (.D(_00002_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[3]$_DFF_PN0_  (.D(_00003_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_valid ),
    .RESET_B(net463),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_4 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4]$_DFF_PN0_  (.D(_00004_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_4 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6]$_DFF_PN0_  (.D(_00005_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[0]$_DFFE_PN0P_  (.D(_00449_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[0] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[10]$_DFFE_PN0P_  (.D(_00450_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[10] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[11]$_DFFE_PN0P_  (.D(_00451_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[11] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[12]$_DFFE_PN0P_  (.D(_00452_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[12] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[13]$_DFFE_PN0P_  (.D(_00453_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[13] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[14]$_DFFE_PN0P_  (.D(_00454_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[14] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[15]$_DFFE_PN0P_  (.D(_00455_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[15] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[16]$_DFFE_PN0P_  (.D(_00456_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[16] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[17]$_DFFE_PN0P_  (.D(_00457_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[17] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[18]$_DFFE_PN0P_  (.D(_00458_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[18] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[19]$_DFFE_PN0P_  (.D(_00459_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[19] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[1]$_DFFE_PN0P_  (.D(_00460_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[1] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[20]$_DFFE_PN0P_  (.D(_00461_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[20] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[21]$_DFFE_PN0P_  (.D(_00462_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[21] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[22]$_DFFE_PN0P_  (.D(_00463_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[22] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[23]$_DFFE_PN0P_  (.D(_00464_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[23] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[24]$_DFFE_PN0P_  (.D(_00465_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[24] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[25]$_DFFE_PN0P_  (.D(_00466_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[25] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[26]$_DFFE_PN0P_  (.D(_00467_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[26] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[27]$_DFFE_PN0P_  (.D(_00468_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[27] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[28]$_DFFE_PN0P_  (.D(_00469_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[28] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[29]$_DFFE_PN0P_  (.D(_00470_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[29] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[2]$_DFFE_PN0P_  (.D(_00471_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[2] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[30]$_DFFE_PN0P_  (.D(_00472_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[30] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[31]$_DFFE_PN0P_  (.D(_00473_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[3]$_DFFE_PN0P_  (.D(_00474_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[3] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[4]$_DFFE_PN0P_  (.D(_00475_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[4] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[5]$_DFFE_PN0P_  (.D(_00476_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[5] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[6]$_DFFE_PN0P_  (.D(_00477_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[6] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[7]$_DFFE_PN0P_  (.D(_00478_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[7] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[8]$_DFFE_PN0P_  (.D(_00479_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[8] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[9]$_DFFE_PN0P_  (.D(_00480_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[9] ),
    .RESET_B(net461),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[0]$_DFFE_PN0P_  (.D(_00481_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[0] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[10]$_DFFE_PN0P_  (.D(_00482_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[10] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[11]$_DFFE_PN0P_  (.D(_00483_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[11] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[12]$_DFFE_PN0P_  (.D(_00484_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[12] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[13]$_DFFE_PN0P_  (.D(_00485_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[13] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[14]$_DFFE_PN0P_  (.D(_00486_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[14] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[15]$_DFFE_PN0P_  (.D(_00487_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[15] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[16]$_DFFE_PN0P_  (.D(_00488_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[16] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[17]$_DFFE_PN0P_  (.D(_00489_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[17] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[18]$_DFFE_PN0P_  (.D(_00490_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[18] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[19]$_DFFE_PN0P_  (.D(_00491_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[19] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[1]$_DFFE_PN0P_  (.D(_00492_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[1] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[20]$_DFFE_PN0P_  (.D(_00493_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[20] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[21]$_DFFE_PN0P_  (.D(_00494_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[21] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[22]$_DFFE_PN0P_  (.D(_00495_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[22] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[23]$_DFFE_PN0P_  (.D(_00496_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[23] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[24]$_DFFE_PN0P_  (.D(_00497_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[24] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[25]$_DFFE_PN0P_  (.D(_00498_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[25] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[26]$_DFFE_PN0P_  (.D(_00499_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[26] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[27]$_DFFE_PN0P_  (.D(_00500_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[27] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[28]$_DFFE_PN0P_  (.D(_00501_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[28] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[29]$_DFFE_PN0P_  (.D(_00502_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[29] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[2]$_DFFE_PN0P_  (.D(_00503_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[2] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[30]$_DFFE_PN0P_  (.D(_00504_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[30] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[31]$_DFFE_PN0P_  (.D(_00505_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[31] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[3]$_DFFE_PN0P_  (.D(_00506_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[3] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[4]$_DFFE_PN0P_  (.D(_00507_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[4] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[5]$_DFFE_PN0P_  (.D(_00508_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[5] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[6]$_DFFE_PN0P_  (.D(_00509_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[6] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[7]$_DFFE_PN0P_  (.D(_00510_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[7] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[8]$_DFFE_PN0P_  (.D(_00511_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[8] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfrtp_1 \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[9]$_DFFE_PN0P_  (.D(_00512_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfrtp_1 \fetch_enable_q$_DFFE_PN0P_  (.D(_00513_),
    .Q(fetch_enable_q),
    .RESET_B(net466),
    .CLK(clknet_leaf_21_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[0]$_DFFE_PN0P_  (.D(_00514_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[32] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_32_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[100]$_DFFE_PN0P_  (.D(_00515_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[132] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_16_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[101]$_DFFE_PN0P_  (.D(_00516_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[133] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_16_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[102]$_DFFE_PN0P_  (.D(_00517_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[134] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_22_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[103]$_DFFE_PN0P_  (.D(_00518_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[135] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_25_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[104]$_DFFE_PN0P_  (.D(_00519_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[136] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_41_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[105]$_DFFE_PN0P_  (.D(_00520_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[137] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_34_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[106]$_DFFE_PN0P_  (.D(_00521_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[138] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_14_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[107]$_DFFE_PN0P_  (.D(_00522_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[139] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_16_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[108]$_DFFE_PN0P_  (.D(_00523_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[140] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_29_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[109]$_DFFE_PN0P_  (.D(_00524_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[141] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_34_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[10]$_DFFE_PN0P_  (.D(_00525_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[42] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_13_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[110]$_DFFE_PN0P_  (.D(_00526_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[142] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_27_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[111]$_DFFE_PN0P_  (.D(_00527_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[143] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_33_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[112]$_DFFE_PN0P_  (.D(_00528_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[144] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_30_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[113]$_DFFE_PN0P_  (.D(_00529_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[145] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_33_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[114]$_DFFE_PN0P_  (.D(_00530_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[146] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_12_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[115]$_DFFE_PN0P_  (.D(_00531_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[147] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_41_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[116]$_DFFE_PN0P_  (.D(_00532_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[148] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_15_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[117]$_DFFE_PN0P_  (.D(_00533_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[149] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_24_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[118]$_DFFE_PN0P_  (.D(_00534_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[150] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_16_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[119]$_DFFE_PN0P_  (.D(_00535_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[151] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_23_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[11]$_DFFE_PN0P_  (.D(_00536_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[43] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_14_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[120]$_DFFE_PN0P_  (.D(_00537_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[152] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_26_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[121]$_DFFE_PN0P_  (.D(_00538_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[153] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_28_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[122]$_DFFE_PN0P_  (.D(_00539_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[154] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_23_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[123]$_DFFE_PN0P_  (.D(_00540_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[155] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_24_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[124]$_DFFE_PN0P_  (.D(_00541_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[156] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_24_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[125]$_DFFE_PN0P_  (.D(_00542_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[157] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_34_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[126]$_DFFE_PN0P_  (.D(_00543_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[158] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_28_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[127]$_DFFE_PN0P_  (.D(_00544_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[159] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_30_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[128]$_DFFE_PN0P_  (.D(_00545_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[160] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_32_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[129]$_DFFE_PN0P_  (.D(_00546_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[161] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_30_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[12]$_DFFE_PN0P_  (.D(_00547_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[44] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_28_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[130]$_DFFE_PN0P_  (.D(_00548_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[162] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_32_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[131]$_DFFE_PN0P_  (.D(_00549_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[163] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_39_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[132]$_DFFE_PN0P_  (.D(_00550_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[164] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_17_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[133]$_DFFE_PN0P_  (.D(_00551_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[165] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_17_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[134]$_DFFE_PN0P_  (.D(_00552_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[166] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_22_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[135]$_DFFE_PN0P_  (.D(_00553_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[167] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_23_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[136]$_DFFE_PN0P_  (.D(_00554_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[168] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_36_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[137]$_DFFE_PN0P_  (.D(_00555_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[169] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_29_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[138]$_DFFE_PN0P_  (.D(_00556_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[170] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_14_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[139]$_DFFE_PN0P_  (.D(_00557_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[171] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_18_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[13]$_DFFE_PN0P_  (.D(_00558_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[45] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_35_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[140]$_DFFE_PN0P_  (.D(_00559_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[172] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_24_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[141]$_DFFE_PN0P_  (.D(_00560_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[173] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_34_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[142]$_DFFE_PN0P_  (.D(_00561_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[174] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_26_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[143]$_DFFE_PN0P_  (.D(_00562_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[175] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_34_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[144]$_DFFE_PN0P_  (.D(_00563_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[176] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_30_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[145]$_DFFE_PN0P_  (.D(_00564_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[177] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_34_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[146]$_DFFE_PN0P_  (.D(_00565_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[178] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_38_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[147]$_DFFE_PN0P_  (.D(_00566_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[179] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_41_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[148]$_DFFE_PN0P_  (.D(_00567_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[180] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_18_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[149]$_DFFE_PN0P_  (.D(_00568_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[181] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_24_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[14]$_DFFE_PN0P_  (.D(_00569_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[46] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_26_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[150]$_DFFE_PN0P_  (.D(_00570_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[182] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_16_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[151]$_DFFE_PN0P_  (.D(_00571_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[183] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_22_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[152]$_DFFE_PN0P_  (.D(_00572_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[184] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_26_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[153]$_DFFE_PN0P_  (.D(_00573_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[185] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_28_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[154]$_DFFE_PN0P_  (.D(_00574_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[186] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_22_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[155]$_DFFE_PN0P_  (.D(_00575_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[187] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_23_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[156]$_DFFE_PN0P_  (.D(_00576_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[188] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_24_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[157]$_DFFE_PN0P_  (.D(_00577_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[189] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_34_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[158]$_DFFE_PN0P_  (.D(_00578_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[190] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_28_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[159]$_DFFE_PN0P_  (.D(_00579_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[191] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_30_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[15]$_DFFE_PN0P_  (.D(_00580_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[47] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_33_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[160]$_DFFE_PN0P_  (.D(_00581_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[192] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_35_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[161]$_DFFE_PN0P_  (.D(_00582_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[193] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_31_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[162]$_DFFE_PN0P_  (.D(_00583_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[194] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_36_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[163]$_DFFE_PN0P_  (.D(_00584_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[195] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_38_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[164]$_DFFE_PN0P_  (.D(_00585_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[196] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_17_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[165]$_DFFE_PN0P_  (.D(_00586_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[197] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_17_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[166]$_DFFE_PN0P_  (.D(_00587_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[198] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_16_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[167]$_DFFE_PN0P_  (.D(_00588_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[199] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_23_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[168]$_DFFE_PN0P_  (.D(_00589_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[200] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_37_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[169]$_DFFE_PN0P_  (.D(_00590_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[201] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_28_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[16]$_DFFE_PN0P_  (.D(_00591_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[48] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_31_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[170]$_DFFE_PN0P_  (.D(_00592_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[202] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_18_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[171]$_DFFE_PN0P_  (.D(_00593_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[203] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_18_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[172]$_DFFE_PN0P_  (.D(_00594_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[204] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_24_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[173]$_DFFE_PN0P_  (.D(_00595_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[205] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_34_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[174]$_DFFE_PN0P_  (.D(_00596_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[206] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_27_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[175]$_DFFE_PN0P_  (.D(_00597_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[207] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_34_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[176]$_DFFE_PN0P_  (.D(_00598_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[208] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_31_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[177]$_DFFE_PN0P_  (.D(_00599_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[209] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_35_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[178]$_DFFE_PN0P_  (.D(_00600_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[210] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_39_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[179]$_DFFE_PN0P_  (.D(_00601_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[211] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_36_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[17]$_DFFE_PN0P_  (.D(_00602_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[49] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_35_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[180]$_DFFE_PN0P_  (.D(_00603_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[212] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_18_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[181]$_DFFE_PN0P_  (.D(_00604_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[213] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_23_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[182]$_DFFE_PN0P_  (.D(_00605_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[214] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_17_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[183]$_DFFE_PN0P_  (.D(_00606_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[215] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_22_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[184]$_DFFE_PN0P_  (.D(_00607_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[216] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_26_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[185]$_DFFE_PN0P_  (.D(_00608_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[217] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_28_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[186]$_DFFE_PN0P_  (.D(_00609_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[218] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_22_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[187]$_DFFE_PN0P_  (.D(_00610_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[219] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_23_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[188]$_DFFE_PN0P_  (.D(_00611_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[220] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_25_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[189]$_DFFE_PN0P_  (.D(_00612_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[221] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_37_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[18]$_DFFE_PN0P_  (.D(_00613_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[50] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_38_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[190]$_DFFE_PN0P_  (.D(_00614_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[222] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_27_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[191]$_DFFE_PN0P_  (.D(_00615_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[223] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_31_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[192]$_DFFE_PN0P_  (.D(_00616_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[224] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_32_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[193]$_DFFE_PN0P_  (.D(_00617_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[225] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_30_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[194]$_DFFE_PN0P_  (.D(_00618_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[226] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_36_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[195]$_DFFE_PN0P_  (.D(_00619_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[227] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_38_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[196]$_DFFE_PN0P_  (.D(_00620_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[228] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_17_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[197]$_DFFE_PN0P_  (.D(_00621_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[229] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_17_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[198]$_DFFE_PN0P_  (.D(_00622_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[230] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_22_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[199]$_DFFE_PN0P_  (.D(_00623_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[231] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_23_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[19]$_DFFE_PN0P_  (.D(_00624_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[51] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_36_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[1]$_DFFE_PN0P_  (.D(_00625_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[33] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_31_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[200]$_DFFE_PN0P_  (.D(_00626_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[232] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_37_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[201]$_DFFE_PN0P_  (.D(_00627_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[233] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_28_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[202]$_DFFE_PN0P_  (.D(_00628_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[234] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_18_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[203]$_DFFE_PN0P_  (.D(_00629_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[235] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_18_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[204]$_DFFE_PN0P_  (.D(_00630_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[236] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_24_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[205]$_DFFE_PN0P_  (.D(_00631_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[237] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_34_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[206]$_DFFE_PN0P_  (.D(_00632_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[238] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_27_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[207]$_DFFE_PN0P_  (.D(_00633_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[239] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_34_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[208]$_DFFE_PN0P_  (.D(_00634_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[240] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_30_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[209]$_DFFE_PN0P_  (.D(_00635_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[241] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_35_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[20]$_DFFE_PN0P_  (.D(_00636_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[52] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_13_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[210]$_DFFE_PN0P_  (.D(_00637_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[242] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_27_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[211]$_DFFE_PN0P_  (.D(_00638_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[243] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_36_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[212]$_DFFE_PN0P_  (.D(_00639_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[244] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_18_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[213]$_DFFE_PN0P_  (.D(_00640_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[245] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_24_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[214]$_DFFE_PN0P_  (.D(_00641_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[246] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_16_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[215]$_DFFE_PN0P_  (.D(_00642_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[247] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_22_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[216]$_DFFE_PN0P_  (.D(_00643_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[248] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_26_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[217]$_DFFE_PN0P_  (.D(_00644_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[249] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_29_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[218]$_DFFE_PN0P_  (.D(_00645_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[250] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_22_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[219]$_DFFE_PN0P_  (.D(_00646_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[251] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_23_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[21]$_DFFE_PN0P_  (.D(_00647_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[53] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_25_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[220]$_DFFE_PN0P_  (.D(_00648_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[252] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_24_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[221]$_DFFE_PN0P_  (.D(_00649_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[253] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_35_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[222]$_DFFE_PN0P_  (.D(_00650_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[254] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_27_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[223]$_DFFE_PN0P_  (.D(_00651_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[255] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_30_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[224]$_DFFE_PN0P_  (.D(_00652_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[256] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[225]$_DFFE_PN0P_  (.D(_00653_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[257] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_51_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[226]$_DFFE_PN0P_  (.D(_00654_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[258] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_60_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[227]$_DFFE_PN0P_  (.D(_00655_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[259] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_52_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[228]$_DFFE_PN0P_  (.D(_00656_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[260] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_94_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[229]$_DFFE_PN0P_  (.D(_00657_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[261] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_4_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[22]$_DFFE_PN0P_  (.D(_00658_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[54] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_16_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[230]$_DFFE_PN0P_  (.D(_00659_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[262] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_95_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[231]$_DFFE_PN0P_  (.D(_00660_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[263] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_19_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[232]$_DFFE_PN0P_  (.D(_00661_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[264] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[233]$_DFFE_PN0P_  (.D(_00662_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[265] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_75_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[234]$_DFFE_PN0P_  (.D(_00663_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[266] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_98_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[235]$_DFFE_PN0P_  (.D(_00664_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[267] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_92_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[236]$_DFFE_PN0P_  (.D(_00665_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[268] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_80_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[237]$_DFFE_PN0P_  (.D(_00666_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[269] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_54_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[238]$_DFFE_PN0P_  (.D(_00667_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[270] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[239]$_DFFE_PN0P_  (.D(_00668_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[271] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_60_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[23]$_DFFE_PN0P_  (.D(_00669_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[55] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_25_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[240]$_DFFE_PN0P_  (.D(_00670_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[272] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[241]$_DFFE_PN0P_  (.D(_00671_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[273] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[242]$_DFFE_PN0P_  (.D(_00672_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[274] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[243]$_DFFE_PN0P_  (.D(_00673_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[275] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_63_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[244]$_DFFE_PN0P_  (.D(_00674_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[276] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_19_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[245]$_DFFE_PN0P_  (.D(_00675_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[277] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_88_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[246]$_DFFE_PN0P_  (.D(_00676_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[278] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_5_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[247]$_DFFE_PN0P_  (.D(_00677_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[279] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_95_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[248]$_DFFE_PN0P_  (.D(_00678_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[280] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_11_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[249]$_DFFE_PN0P_  (.D(_00679_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[281] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_69_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[24]$_DFFE_PN0P_  (.D(_00680_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[56] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_26_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[250]$_DFFE_PN0P_  (.D(_00681_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[282] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_90_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[251]$_DFFE_PN0P_  (.D(_00682_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[283] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[252]$_DFFE_PN0P_  (.D(_00683_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[284] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_12_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[253]$_DFFE_PN0P_  (.D(_00684_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[285] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_43_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[254]$_DFFE_PN0P_  (.D(_00685_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[286] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_63_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[255]$_DFFE_PN0P_  (.D(_00686_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[287] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_46_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[256]$_DFFE_PN0P_  (.D(_00687_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[288] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[257]$_DFFE_PN0P_  (.D(_00688_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[289] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_51_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[258]$_DFFE_PN0P_  (.D(_00689_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[290] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_60_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[259]$_DFFE_PN0P_  (.D(_00690_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[291] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[25]$_DFFE_PN0P_  (.D(_00691_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[57] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_27_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[260]$_DFFE_PN0P_  (.D(_00692_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[292] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_94_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[261]$_DFFE_PN0P_  (.D(_00693_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[293] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_4_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[262]$_DFFE_PN0P_  (.D(_00694_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[294] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_97_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[263]$_DFFE_PN0P_  (.D(_00695_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[295] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_19_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[264]$_DFFE_PN0P_  (.D(_00696_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[296] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_63_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[265]$_DFFE_PN0P_  (.D(_00697_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[297] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_74_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[266]$_DFFE_PN0P_  (.D(_00698_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[298] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_99_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[267]$_DFFE_PN0P_  (.D(_00699_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[299] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_96_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[268]$_DFFE_PN0P_  (.D(_00700_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[300] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_80_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[269]$_DFFE_PN0P_  (.D(_00701_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[301] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_61_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[26]$_DFFE_PN0P_  (.D(_00702_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[58] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_13_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[270]$_DFFE_PN0P_  (.D(_00703_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[302] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_14_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[271]$_DFFE_PN0P_  (.D(_00704_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[303] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_61_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[272]$_DFFE_PN0P_  (.D(_00705_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[304] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[273]$_DFFE_PN0P_  (.D(_00706_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[305] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_52_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[274]$_DFFE_PN0P_  (.D(_00707_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[306] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_69_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[275]$_DFFE_PN0P_  (.D(_00708_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[307] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_64_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[276]$_DFFE_PN0P_  (.D(_00709_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[308] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_18_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[277]$_DFFE_PN0P_  (.D(_00710_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[309] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[278]$_DFFE_PN0P_  (.D(_00711_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[310] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_5_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[279]$_DFFE_PN0P_  (.D(_00712_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[311] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_95_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[27]$_DFFE_PN0P_  (.D(_00713_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[59] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_13_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[280]$_DFFE_PN0P_  (.D(_00714_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[312] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_11_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[281]$_DFFE_PN0P_  (.D(_00715_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[313] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[282]$_DFFE_PN0P_  (.D(_00716_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[314] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_92_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[283]$_DFFE_PN0P_  (.D(_00717_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[315] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_80_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[284]$_DFFE_PN0P_  (.D(_00718_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[316] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_12_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[285]$_DFFE_PN0P_  (.D(_00719_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[317] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_73_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[286]$_DFFE_PN0P_  (.D(_00720_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[318] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[287]$_DFFE_PN0P_  (.D(_00721_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[319] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_45_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[288]$_DFFE_PN0P_  (.D(_00722_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[320] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[289]$_DFFE_PN0P_  (.D(_00723_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[321] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_51_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[28]$_DFFE_PN0P_  (.D(_00724_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[60] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_25_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[290]$_DFFE_PN0P_  (.D(_00725_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[322] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_60_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[291]$_DFFE_PN0P_  (.D(_00726_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[323] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_72_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[292]$_DFFE_PN0P_  (.D(_00727_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[324] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_98_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[293]$_DFFE_PN0P_  (.D(_00728_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[325] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_4_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[294]$_DFFE_PN0P_  (.D(_00729_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[326] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_97_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[295]$_DFFE_PN0P_  (.D(_00730_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[327] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_19_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[296]$_DFFE_PN0P_  (.D(_00731_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[328] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_63_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[297]$_DFFE_PN0P_  (.D(_00732_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[329] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_75_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[298]$_DFFE_PN0P_  (.D(_00733_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[330] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_99_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[299]$_DFFE_PN0P_  (.D(_00734_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[331] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_96_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[29]$_DFFE_PN0P_  (.D(_00735_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[61] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_35_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[2]$_DFFE_PN0P_  (.D(_00736_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[34] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_31_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[300]$_DFFE_PN0P_  (.D(_00737_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[332] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_79_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[301]$_DFFE_PN0P_  (.D(_00738_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[333] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_60_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[302]$_DFFE_PN0P_  (.D(_00739_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[334] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[303]$_DFFE_PN0P_  (.D(_00740_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[335] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_61_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[304]$_DFFE_PN0P_  (.D(_00741_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[336] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[305]$_DFFE_PN0P_  (.D(_00742_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[337] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_52_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[306]$_DFFE_PN0P_  (.D(_00743_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[338] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[307]$_DFFE_PN0P_  (.D(_00744_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[339] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_64_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[308]$_DFFE_PN0P_  (.D(_00745_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[340] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_19_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[309]$_DFFE_PN0P_  (.D(_00746_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[341] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_69_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[30]$_DFFE_PN0P_  (.D(_00747_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[62] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_38_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[310]$_DFFE_PN0P_  (.D(_00748_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[342] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_5_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[311]$_DFFE_PN0P_  (.D(_00749_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[343] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_95_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[312]$_DFFE_PN0P_  (.D(_00750_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[344] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_10_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[313]$_DFFE_PN0P_  (.D(_00751_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[345] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_69_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[314]$_DFFE_PN0P_  (.D(_00752_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[346] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_92_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[315]$_DFFE_PN0P_  (.D(_00753_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[347] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[316]$_DFFE_PN0P_  (.D(_00754_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[348] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_11_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[317]$_DFFE_PN0P_  (.D(_00755_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[349] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_43_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[318]$_DFFE_PN0P_  (.D(_00756_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[350] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[319]$_DFFE_PN0P_  (.D(_00757_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[351] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_48_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[31]$_DFFE_PN0P_  (.D(_00758_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[63] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_31_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[320]$_DFFE_PN0P_  (.D(_00759_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[352] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_54_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[321]$_DFFE_PN0P_  (.D(_00760_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[353] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_51_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[322]$_DFFE_PN0P_  (.D(_00761_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[354] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_60_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[323]$_DFFE_PN0P_  (.D(_00762_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[355] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_72_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[324]$_DFFE_PN0P_  (.D(_00763_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[356] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_98_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[325]$_DFFE_PN0P_  (.D(_00764_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[357] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_4_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[326]$_DFFE_PN0P_  (.D(_00765_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[358] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_97_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[327]$_DFFE_PN0P_  (.D(_00766_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[359] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_19_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[328]$_DFFE_PN0P_  (.D(_00767_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[360] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_63_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[329]$_DFFE_PN0P_  (.D(_00768_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[361] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_74_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[32]$_DFFE_PN0P_  (.D(_00769_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[64] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_33_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[330]$_DFFE_PN0P_  (.D(_00770_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[362] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_99_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[331]$_DFFE_PN0P_  (.D(_00771_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[363] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_93_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[332]$_DFFE_PN0P_  (.D(_00772_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[364] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_79_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[333]$_DFFE_PN0P_  (.D(_00773_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[365] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_60_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[334]$_DFFE_PN0P_  (.D(_00774_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[366] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_14_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[335]$_DFFE_PN0P_  (.D(_00775_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[367] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_60_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[336]$_DFFE_PN0P_  (.D(_00776_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[368] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[337]$_DFFE_PN0P_  (.D(_00777_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[369] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_51_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[338]$_DFFE_PN0P_  (.D(_00778_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[370] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[339]$_DFFE_PN0P_  (.D(_00779_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[371] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_61_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[33]$_DFFE_PN0P_  (.D(_00780_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[65] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_31_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[340]$_DFFE_PN0P_  (.D(_00781_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[372] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_19_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[341]$_DFFE_PN0P_  (.D(_00782_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[373] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[342]$_DFFE_PN0P_  (.D(_00783_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[374] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[343]$_DFFE_PN0P_  (.D(_00784_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[375] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_95_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[344]$_DFFE_PN0P_  (.D(_00785_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[376] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_10_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[345]$_DFFE_PN0P_  (.D(_00786_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[377] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_69_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[346]$_DFFE_PN0P_  (.D(_00787_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[378] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_92_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[347]$_DFFE_PN0P_  (.D(_00788_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[379] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_85_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[348]$_DFFE_PN0P_  (.D(_00789_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[380] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_78_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[349]$_DFFE_PN0P_  (.D(_00790_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[381] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_43_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[34]$_DFFE_PN0P_  (.D(_00791_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[66] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_32_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[350]$_DFFE_PN0P_  (.D(_00792_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[382] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[351]$_DFFE_PN0P_  (.D(_00793_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[383] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_48_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[352]$_DFFE_PN0P_  (.D(_00794_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[384] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_55_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[353]$_DFFE_PN0P_  (.D(_00795_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[385] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_51_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[354]$_DFFE_PN0P_  (.D(_00796_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[386] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[355]$_DFFE_PN0P_  (.D(_00797_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[387] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_72_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[356]$_DFFE_PN0P_  (.D(_00798_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[388] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_98_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[357]$_DFFE_PN0P_  (.D(_00799_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[389] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_20_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[358]$_DFFE_PN0P_  (.D(_00800_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[390] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_97_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[359]$_DFFE_PN0P_  (.D(_00801_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[391] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_3_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[35]$_DFFE_PN0P_  (.D(_00802_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[67] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_38_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[360]$_DFFE_PN0P_  (.D(_00803_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[392] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[361]$_DFFE_PN0P_  (.D(_00804_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[393] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_72_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[362]$_DFFE_PN0P_  (.D(_00805_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[394] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_1_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[363]$_DFFE_PN0P_  (.D(_00806_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[395] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_96_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[364]$_DFFE_PN0P_  (.D(_00807_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[396] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_80_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[365]$_DFFE_PN0P_  (.D(_00808_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[397] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_57_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[366]$_DFFE_PN0P_  (.D(_00809_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[398] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_19_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[367]$_DFFE_PN0P_  (.D(_00810_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[399] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_59_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_2 \gen_regfile_ff.register_file_i.rf_reg_q[368]$_DFFE_PN0P_  (.D(_00811_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[400] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[369]$_DFFE_PN0P_  (.D(_00812_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[401] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_52_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[36]$_DFFE_PN0P_  (.D(_00813_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[68] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_16_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[370]$_DFFE_PN0P_  (.D(_00814_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[402] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[371]$_DFFE_PN0P_  (.D(_00815_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[403] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_64_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[372]$_DFFE_PN0P_  (.D(_00816_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[404] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_18_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[373]$_DFFE_PN0P_  (.D(_00817_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[405] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_88_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[374]$_DFFE_PN0P_  (.D(_00818_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[406] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[375]$_DFFE_PN0P_  (.D(_00819_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[407] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_96_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[376]$_DFFE_PN0P_  (.D(_00820_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[408] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_14_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[377]$_DFFE_PN0P_  (.D(_00821_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[409] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[378]$_DFFE_PN0P_  (.D(_00822_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[410] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[379]$_DFFE_PN0P_  (.D(_00823_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[411] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_85_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[37]$_DFFE_PN0P_  (.D(_00824_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[69] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_15_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[380]$_DFFE_PN0P_  (.D(_00825_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[412] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_11_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[381]$_DFFE_PN0P_  (.D(_00826_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[413] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_73_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[382]$_DFFE_PN0P_  (.D(_00827_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[414] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[383]$_DFFE_PN0P_  (.D(_00828_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[415] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_45_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[384]$_DFFE_PN0P_  (.D(_00829_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[416] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_55_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[385]$_DFFE_PN0P_  (.D(_00830_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[417] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_50_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[386]$_DFFE_PN0P_  (.D(_00831_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[418] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_58_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[387]$_DFFE_PN0P_  (.D(_00832_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[419] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_72_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[388]$_DFFE_PN0P_  (.D(_00833_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[420] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_98_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[389]$_DFFE_PN0P_  (.D(_00834_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[421] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_20_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[38]$_DFFE_PN0P_  (.D(_00835_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[70] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_15_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[390]$_DFFE_PN0P_  (.D(_00836_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[422] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_97_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[391]$_DFFE_PN0P_  (.D(_00837_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[423] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_3_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[392]$_DFFE_PN0P_  (.D(_00838_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[424] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[393]$_DFFE_PN0P_  (.D(_00839_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[425] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_73_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[394]$_DFFE_PN0P_  (.D(_00840_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[426] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_1_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[395]$_DFFE_PN0P_  (.D(_00841_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[427] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_96_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[396]$_DFFE_PN0P_  (.D(_00842_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[428] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_80_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[397]$_DFFE_PN0P_  (.D(_00843_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[429] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_57_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[398]$_DFFE_PN0P_  (.D(_00844_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[430] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_20_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[399]$_DFFE_PN0P_  (.D(_00845_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[431] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_60_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[39]$_DFFE_PN0P_  (.D(_00846_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[71] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_12_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[3]$_DFFE_PN0P_  (.D(_00847_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[35] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_38_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[400]$_DFFE_PN0P_  (.D(_00848_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[432] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_54_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[401]$_DFFE_PN0P_  (.D(_00849_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[433] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_50_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[402]$_DFFE_PN0P_  (.D(_00850_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[434] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[403]$_DFFE_PN0P_  (.D(_00851_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[435] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_64_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[404]$_DFFE_PN0P_  (.D(_00852_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[436] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_18_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[405]$_DFFE_PN0P_  (.D(_00853_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[437] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[406]$_DFFE_PN0P_  (.D(_00854_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[438] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_1_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[407]$_DFFE_PN0P_  (.D(_00855_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[439] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_95_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[408]$_DFFE_PN0P_  (.D(_00856_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[440] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_14_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[409]$_DFFE_PN0P_  (.D(_00857_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[441] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_88_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[40]$_DFFE_PN0P_  (.D(_00858_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[72] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_37_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[410]$_DFFE_PN0P_  (.D(_00859_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[442] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[411]$_DFFE_PN0P_  (.D(_00860_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[443] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_83_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[412]$_DFFE_PN0P_  (.D(_00861_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[444] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_12_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[413]$_DFFE_PN0P_  (.D(_00862_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[445] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_74_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[414]$_DFFE_PN0P_  (.D(_00863_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[446] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[415]$_DFFE_PN0P_  (.D(_00864_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[447] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_45_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[416]$_DFFE_PN0P_  (.D(_00865_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[448] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_54_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[417]$_DFFE_PN0P_  (.D(_00866_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[449] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_50_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[418]$_DFFE_PN0P_  (.D(_00867_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[450] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_57_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[419]$_DFFE_PN0P_  (.D(_00868_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[451] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_72_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[41]$_DFFE_PN0P_  (.D(_00869_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[73] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_28_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[420]$_DFFE_PN0P_  (.D(_00870_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[452] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_98_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[421]$_DFFE_PN0P_  (.D(_00871_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[453] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_20_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[422]$_DFFE_PN0P_  (.D(_00872_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[454] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_97_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[423]$_DFFE_PN0P_  (.D(_00873_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[455] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[424]$_DFFE_PN0P_  (.D(_00874_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[456] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[425]$_DFFE_PN0P_  (.D(_00875_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[457] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_73_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[426]$_DFFE_PN0P_  (.D(_00876_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[458] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_1_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[427]$_DFFE_PN0P_  (.D(_00877_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[459] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_96_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[428]$_DFFE_PN0P_  (.D(_00878_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[460] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[429]$_DFFE_PN0P_  (.D(_00879_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[461] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[42]$_DFFE_PN0P_  (.D(_00880_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[74] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_13_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[430]$_DFFE_PN0P_  (.D(_00881_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[462] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_20_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[431]$_DFFE_PN0P_  (.D(_00882_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[463] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_59_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_2 \gen_regfile_ff.register_file_i.rf_reg_q[432]$_DFFE_PN0P_  (.D(_00883_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[464] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[433]$_DFFE_PN0P_  (.D(_00884_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[465] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_50_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[434]$_DFFE_PN0P_  (.D(_00885_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[466] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[435]$_DFFE_PN0P_  (.D(_00886_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[467] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_64_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[436]$_DFFE_PN0P_  (.D(_00887_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[468] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_19_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[437]$_DFFE_PN0P_  (.D(_00888_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[469] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[438]$_DFFE_PN0P_  (.D(_00889_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[470] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[439]$_DFFE_PN0P_  (.D(_00890_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[471] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_95_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[43]$_DFFE_PN0P_  (.D(_00891_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[75] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_14_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[440]$_DFFE_PN0P_  (.D(_00892_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[472] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_10_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[441]$_DFFE_PN0P_  (.D(_00893_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[473] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_69_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[442]$_DFFE_PN0P_  (.D(_00894_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[474] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_92_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[443]$_DFFE_PN0P_  (.D(_00895_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[475] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_82_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[444]$_DFFE_PN0P_  (.D(_00896_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[476] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_11_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[445]$_DFFE_PN0P_  (.D(_00897_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[477] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_43_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[446]$_DFFE_PN0P_  (.D(_00898_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[478] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[447]$_DFFE_PN0P_  (.D(_00899_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[479] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_49_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[448]$_DFFE_PN0P_  (.D(_00900_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[480] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_55_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[449]$_DFFE_PN0P_  (.D(_00901_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[481] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_50_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[44]$_DFFE_PN0P_  (.D(_00902_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[76] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_25_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[450]$_DFFE_PN0P_  (.D(_00903_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[482] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[451]$_DFFE_PN0P_  (.D(_00904_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[483] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[452]$_DFFE_PN0P_  (.D(_00905_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[484] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_98_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[453]$_DFFE_PN0P_  (.D(_00906_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[485] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_20_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[454]$_DFFE_PN0P_  (.D(_00907_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[486] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_97_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[455]$_DFFE_PN0P_  (.D(_00908_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[487] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[456]$_DFFE_PN0P_  (.D(_00909_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[488] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[457]$_DFFE_PN0P_  (.D(_00910_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[489] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_73_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[458]$_DFFE_PN0P_  (.D(_00911_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[490] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_1_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[459]$_DFFE_PN0P_  (.D(_00912_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[491] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_96_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[45]$_DFFE_PN0P_  (.D(_00913_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[77] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_35_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[460]$_DFFE_PN0P_  (.D(_00914_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[492] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[461]$_DFFE_PN0P_  (.D(_00915_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[493] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_57_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[462]$_DFFE_PN0P_  (.D(_00916_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[494] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_20_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[463]$_DFFE_PN0P_  (.D(_00917_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[495] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_60_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[464]$_DFFE_PN0P_  (.D(_00918_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[496] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[465]$_DFFE_PN0P_  (.D(_00919_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[497] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_52_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[466]$_DFFE_PN0P_  (.D(_00920_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[498] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[467]$_DFFE_PN0P_  (.D(_00921_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[499] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_64_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[468]$_DFFE_PN0P_  (.D(_00922_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[500] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_19_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[469]$_DFFE_PN0P_  (.D(_00923_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[501] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[46]$_DFFE_PN0P_  (.D(_00924_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[78] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_26_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[470]$_DFFE_PN0P_  (.D(_00925_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[502] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_1_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[471]$_DFFE_PN0P_  (.D(_00926_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[503] ),
    .RESET_B(net148),
    .CLK(clknet_leaf_95_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[472]$_DFFE_PN0P_  (.D(_00927_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[504] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_10_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[473]$_DFFE_PN0P_  (.D(_00928_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[505] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_69_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[474]$_DFFE_PN0P_  (.D(_00929_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[506] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_90_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[475]$_DFFE_PN0P_  (.D(_00930_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[507] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_82_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[476]$_DFFE_PN0P_  (.D(_00931_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[508] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_11_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[477]$_DFFE_PN0P_  (.D(_00932_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[509] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_43_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[478]$_DFFE_PN0P_  (.D(_00933_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[510] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[479]$_DFFE_PN0P_  (.D(_00934_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[511] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_49_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[47]$_DFFE_PN0P_  (.D(_00935_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[79] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_33_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[480]$_DFFE_PN0P_  (.D(_00936_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[512] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_55_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[481]$_DFFE_PN0P_  (.D(_00937_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[513] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_51_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[482]$_DFFE_PN0P_  (.D(_00938_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[514] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_58_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[483]$_DFFE_PN0P_  (.D(_00939_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[515] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_61_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[484]$_DFFE_PN0P_  (.D(_00940_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[516] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_7_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[485]$_DFFE_PN0P_  (.D(_00941_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[517] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[486]$_DFFE_PN0P_  (.D(_00942_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[518] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_93_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[487]$_DFFE_PN0P_  (.D(_00943_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[519] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_79_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[488]$_DFFE_PN0P_  (.D(_00944_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[520] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[489]$_DFFE_PN0P_  (.D(_00945_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[521] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_71_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[48]$_DFFE_PN0P_  (.D(_00946_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[80] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_32_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[490]$_DFFE_PN0P_  (.D(_00947_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[522] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_91_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[491]$_DFFE_PN0P_  (.D(_00948_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[523] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_91_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[492]$_DFFE_PN0P_  (.D(_00949_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[524] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_80_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[493]$_DFFE_PN0P_  (.D(_00950_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[525] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_57_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[494]$_DFFE_PN0P_  (.D(_00951_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[526] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_78_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[495]$_DFFE_PN0P_  (.D(_00952_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[527] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_59_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[496]$_DFFE_PN0P_  (.D(_00953_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[528] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_57_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[497]$_DFFE_PN0P_  (.D(_00954_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[529] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_55_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[498]$_DFFE_PN0P_  (.D(_00955_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[530] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_76_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[499]$_DFFE_PN0P_  (.D(_00956_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[531] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_64_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[49]$_DFFE_PN0P_  (.D(_00957_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[81] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_35_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[4]$_DFFE_PN0P_  (.D(_00958_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[36] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_15_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[500]$_DFFE_PN0P_  (.D(_00959_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[532] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_8_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[501]$_DFFE_PN0P_  (.D(_00960_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[533] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_88_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[502]$_DFFE_PN0P_  (.D(_00961_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[534] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_7_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[503]$_DFFE_PN0P_  (.D(_00962_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[535] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[504]$_DFFE_PN0P_  (.D(_00963_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[536] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_76_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[505]$_DFFE_PN0P_  (.D(_00964_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[537] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[506]$_DFFE_PN0P_  (.D(_00965_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[538] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[507]$_DFFE_PN0P_  (.D(_00966_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[539] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_88_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[508]$_DFFE_PN0P_  (.D(_00967_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[540] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_76_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[509]$_DFFE_PN0P_  (.D(_00968_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[541] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_41_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[50]$_DFFE_PN0P_  (.D(_00969_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[82] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_27_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[510]$_DFFE_PN0P_  (.D(_00970_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[542] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_77_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[511]$_DFFE_PN0P_  (.D(_00971_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[543] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_48_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[512]$_DFFE_PN0P_  (.D(_00972_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[544] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_55_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[513]$_DFFE_PN0P_  (.D(_00973_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[545] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_50_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[514]$_DFFE_PN0P_  (.D(_00974_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[546] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_58_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[515]$_DFFE_PN0P_  (.D(_00975_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[547] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[516]$_DFFE_PN0P_  (.D(_00976_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[548] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_82_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[517]$_DFFE_PN0P_  (.D(_00977_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[549] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[518]$_DFFE_PN0P_  (.D(_00978_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[550] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_94_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[519]$_DFFE_PN0P_  (.D(_00979_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[551] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[51]$_DFFE_PN0P_  (.D(_00980_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[83] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_36_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[520]$_DFFE_PN0P_  (.D(_00981_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[552] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[521]$_DFFE_PN0P_  (.D(_00982_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[553] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_70_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[522]$_DFFE_PN0P_  (.D(_00983_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[554] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_91_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[523]$_DFFE_PN0P_  (.D(_00984_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[555] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_92_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[524]$_DFFE_PN0P_  (.D(_00985_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[556] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_80_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[525]$_DFFE_PN0P_  (.D(_00986_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[557] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_57_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[526]$_DFFE_PN0P_  (.D(_00987_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[558] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_39_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[527]$_DFFE_PN0P_  (.D(_00988_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[559] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_59_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[528]$_DFFE_PN0P_  (.D(_00989_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[560] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[529]$_DFFE_PN0P_  (.D(_00990_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[561] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_55_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[52]$_DFFE_PN0P_  (.D(_00991_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[84] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_13_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[530]$_DFFE_PN0P_  (.D(_00992_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[562] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_75_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[531]$_DFFE_PN0P_  (.D(_00993_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[563] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_64_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[532]$_DFFE_PN0P_  (.D(_00994_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[564] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[533]$_DFFE_PN0P_  (.D(_00995_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[565] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_88_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[534]$_DFFE_PN0P_  (.D(_00996_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[566] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_7_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[535]$_DFFE_PN0P_  (.D(_00997_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[567] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_91_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[536]$_DFFE_PN0P_  (.D(_00998_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[568] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_76_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[537]$_DFFE_PN0P_  (.D(_00999_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[569] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[538]$_DFFE_PN0P_  (.D(_01000_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[570] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[539]$_DFFE_PN0P_  (.D(_01001_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[571] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[53]$_DFFE_PN0P_  (.D(_01002_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[85] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_25_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[540]$_DFFE_PN0P_  (.D(_01003_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[572] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_77_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[541]$_DFFE_PN0P_  (.D(_01004_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[573] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_41_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[542]$_DFFE_PN0P_  (.D(_01005_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[574] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_40_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[543]$_DFFE_PN0P_  (.D(_01006_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[575] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_49_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[544]$_DFFE_PN0P_  (.D(_01007_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[576] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_55_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[545]$_DFFE_PN0P_  (.D(_01008_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[577] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_49_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[546]$_DFFE_PN0P_  (.D(_01009_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[578] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_58_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[547]$_DFFE_PN0P_  (.D(_01010_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[579] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_63_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[548]$_DFFE_PN0P_  (.D(_01011_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[580] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_82_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[549]$_DFFE_PN0P_  (.D(_01012_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[581] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_4_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[54]$_DFFE_PN0P_  (.D(_01013_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[86] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_16_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[550]$_DFFE_PN0P_  (.D(_01014_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[582] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_93_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[551]$_DFFE_PN0P_  (.D(_01015_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[583] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_8_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[552]$_DFFE_PN0P_  (.D(_01016_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[584] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[553]$_DFFE_PN0P_  (.D(_01017_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[585] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_70_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[554]$_DFFE_PN0P_  (.D(_01018_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[586] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_96_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[555]$_DFFE_PN0P_  (.D(_01019_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[587] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_92_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[556]$_DFFE_PN0P_  (.D(_01020_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[588] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_80_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[557]$_DFFE_PN0P_  (.D(_01021_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[589] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_57_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[558]$_DFFE_PN0P_  (.D(_01022_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[590] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_39_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[559]$_DFFE_PN0P_  (.D(_01023_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[591] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_59_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[55]$_DFFE_PN0P_  (.D(_01024_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[87] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_15_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[560]$_DFFE_PN0P_  (.D(_01025_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[592] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[561]$_DFFE_PN0P_  (.D(_01026_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[593] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_50_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[562]$_DFFE_PN0P_  (.D(_01027_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[594] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_74_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[563]$_DFFE_PN0P_  (.D(_01028_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[595] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_64_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[564]$_DFFE_PN0P_  (.D(_01029_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[596] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_8_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[565]$_DFFE_PN0P_  (.D(_01030_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[597] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_88_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[566]$_DFFE_PN0P_  (.D(_01031_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[598] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_6_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[567]$_DFFE_PN0P_  (.D(_01032_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[599] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_91_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[568]$_DFFE_PN0P_  (.D(_01033_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[600] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_79_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[569]$_DFFE_PN0P_  (.D(_01034_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[601] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[56]$_DFFE_PN0P_  (.D(_01035_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[88] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_26_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[570]$_DFFE_PN0P_  (.D(_01036_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[602] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[571]$_DFFE_PN0P_  (.D(_01037_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[603] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[572]$_DFFE_PN0P_  (.D(_01038_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[604] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_76_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[573]$_DFFE_PN0P_  (.D(_01039_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[605] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_41_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[574]$_DFFE_PN0P_  (.D(_01040_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[606] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_39_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[575]$_DFFE_PN0P_  (.D(_01041_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[607] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_48_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[576]$_DFFE_PN0P_  (.D(_01042_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[608] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_55_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[577]$_DFFE_PN0P_  (.D(_01043_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[609] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_49_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[578]$_DFFE_PN0P_  (.D(_01044_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[610] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_58_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[579]$_DFFE_PN0P_  (.D(_01045_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[611] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[57]$_DFFE_PN0P_  (.D(_01046_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[89] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_27_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[580]$_DFFE_PN0P_  (.D(_01047_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[612] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_7_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[581]$_DFFE_PN0P_  (.D(_01048_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[613] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[582]$_DFFE_PN0P_  (.D(_01049_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[614] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_94_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[583]$_DFFE_PN0P_  (.D(_01050_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[615] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[584]$_DFFE_PN0P_  (.D(_01051_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[616] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[585]$_DFFE_PN0P_  (.D(_01052_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[617] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_70_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[586]$_DFFE_PN0P_  (.D(_01053_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[618] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_91_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[587]$_DFFE_PN0P_  (.D(_01054_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[619] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_92_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[588]$_DFFE_PN0P_  (.D(_01055_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[620] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_80_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[589]$_DFFE_PN0P_  (.D(_01056_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[621] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_57_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[58]$_DFFE_PN0P_  (.D(_01057_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[90] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_13_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[590]$_DFFE_PN0P_  (.D(_01058_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[622] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_39_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[591]$_DFFE_PN0P_  (.D(_01059_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[623] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_59_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[592]$_DFFE_PN0P_  (.D(_01060_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[624] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_55_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[593]$_DFFE_PN0P_  (.D(_01061_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[625] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_50_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[594]$_DFFE_PN0P_  (.D(_01062_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[626] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_76_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[595]$_DFFE_PN0P_  (.D(_01063_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[627] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_64_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[596]$_DFFE_PN0P_  (.D(_01064_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[628] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[597]$_DFFE_PN0P_  (.D(_01065_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[629] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_88_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[598]$_DFFE_PN0P_  (.D(_01066_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[630] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_6_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[599]$_DFFE_PN0P_  (.D(_01067_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[631] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_90_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[59]$_DFFE_PN0P_  (.D(_01068_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[91] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_26_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[5]$_DFFE_PN0P_  (.D(_01069_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[37] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_14_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[600]$_DFFE_PN0P_  (.D(_01070_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[632] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_76_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[601]$_DFFE_PN0P_  (.D(_01071_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[633] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[602]$_DFFE_PN0P_  (.D(_01072_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[634] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[603]$_DFFE_PN0P_  (.D(_01073_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[635] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[604]$_DFFE_PN0P_  (.D(_01074_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[636] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_77_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[605]$_DFFE_PN0P_  (.D(_01075_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[637] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_41_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[606]$_DFFE_PN0P_  (.D(_01076_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[638] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_40_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[607]$_DFFE_PN0P_  (.D(_01077_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[639] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_48_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[608]$_DFFE_PN0P_  (.D(_01078_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[640] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_54_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[609]$_DFFE_PN0P_  (.D(_01079_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[641] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_51_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[60]$_DFFE_PN0P_  (.D(_01080_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[92] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_25_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[610]$_DFFE_PN0P_  (.D(_01081_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[642] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_59_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[611]$_DFFE_PN0P_  (.D(_01082_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[643] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_63_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[612]$_DFFE_PN0P_  (.D(_01083_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[644] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_83_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[613]$_DFFE_PN0P_  (.D(_01084_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[645] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_10_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[614]$_DFFE_PN0P_  (.D(_01085_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[646] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[615]$_DFFE_PN0P_  (.D(_01086_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[647] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_10_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[616]$_DFFE_PN0P_  (.D(_01087_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[648] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[617]$_DFFE_PN0P_  (.D(_01088_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[649] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_72_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[618]$_DFFE_PN0P_  (.D(_01089_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[650] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_91_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[619]$_DFFE_PN0P_  (.D(_01090_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[651] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_93_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[61]$_DFFE_PN0P_  (.D(_01091_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[93] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_37_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[620]$_DFFE_PN0P_  (.D(_01092_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[652] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_75_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[621]$_DFFE_PN0P_  (.D(_01093_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[653] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_58_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[622]$_DFFE_PN0P_  (.D(_01094_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[654] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_78_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[623]$_DFFE_PN0P_  (.D(_01095_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[655] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_59_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[624]$_DFFE_PN0P_  (.D(_01096_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[656] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[625]$_DFFE_PN0P_  (.D(_01097_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[657] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_54_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[626]$_DFFE_PN0P_  (.D(_01098_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[658] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_75_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[627]$_DFFE_PN0P_  (.D(_01099_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[659] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[628]$_DFFE_PN0P_  (.D(_01100_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[660] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_10_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[629]$_DFFE_PN0P_  (.D(_01101_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[661] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[62]$_DFFE_PN0P_  (.D(_01102_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[94] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_28_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[630]$_DFFE_PN0P_  (.D(_01103_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[662] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_8_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[631]$_DFFE_PN0P_  (.D(_01104_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[663] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_90_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[632]$_DFFE_PN0P_  (.D(_01105_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[664] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_79_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[633]$_DFFE_PN0P_  (.D(_01106_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[665] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[634]$_DFFE_PN0P_  (.D(_01107_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[666] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[635]$_DFFE_PN0P_  (.D(_01108_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[667] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_88_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[636]$_DFFE_PN0P_  (.D(_01109_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[668] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_79_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[637]$_DFFE_PN0P_  (.D(_01110_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[669] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_40_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[638]$_DFFE_PN0P_  (.D(_01111_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[670] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_39_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[639]$_DFFE_PN0P_  (.D(_01112_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[671] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_48_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[63]$_DFFE_PN0P_  (.D(_01113_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[95] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_33_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[640]$_DFFE_PN0P_  (.D(_01114_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[672] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[641]$_DFFE_PN0P_  (.D(_01115_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[673] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_51_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[642]$_DFFE_PN0P_  (.D(_01116_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[674] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_58_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[643]$_DFFE_PN0P_  (.D(_01117_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[675] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_63_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[644]$_DFFE_PN0P_  (.D(_01118_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[676] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_93_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[645]$_DFFE_PN0P_  (.D(_01119_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[677] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_10_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[646]$_DFFE_PN0P_  (.D(_01120_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[678] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_93_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[647]$_DFFE_PN0P_  (.D(_01121_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[679] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_8_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[648]$_DFFE_PN0P_  (.D(_01122_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[680] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[649]$_DFFE_PN0P_  (.D(_01123_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[681] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_72_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[64]$_DFFE_PN0P_  (.D(_01124_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[96] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_33_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[650]$_DFFE_PN0P_  (.D(_01125_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[682] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_91_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[651]$_DFFE_PN0P_  (.D(_01126_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[683] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_90_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[652]$_DFFE_PN0P_  (.D(_01127_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[684] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_75_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[653]$_DFFE_PN0P_  (.D(_01128_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[685] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_58_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[654]$_DFFE_PN0P_  (.D(_01129_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[686] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_77_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[655]$_DFFE_PN0P_  (.D(_01130_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[687] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_59_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[656]$_DFFE_PN0P_  (.D(_01131_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[688] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[657]$_DFFE_PN0P_  (.D(_01132_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[689] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_54_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[658]$_DFFE_PN0P_  (.D(_01133_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[690] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_75_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[659]$_DFFE_PN0P_  (.D(_01134_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[691] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[65]$_DFFE_PN0P_  (.D(_01135_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[97] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_31_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[660]$_DFFE_PN0P_  (.D(_01136_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[692] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_8_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[661]$_DFFE_PN0P_  (.D(_01137_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[693] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[662]$_DFFE_PN0P_  (.D(_01138_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[694] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_7_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[663]$_DFFE_PN0P_  (.D(_01139_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[695] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_90_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[664]$_DFFE_PN0P_  (.D(_01140_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[696] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_79_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[665]$_DFFE_PN0P_  (.D(_01141_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[697] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[666]$_DFFE_PN0P_  (.D(_01142_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[698] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_90_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[667]$_DFFE_PN0P_  (.D(_01143_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[699] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[668]$_DFFE_PN0P_  (.D(_01144_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[700] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_79_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[669]$_DFFE_PN0P_  (.D(_01145_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[701] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_42_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[66]$_DFFE_PN0P_  (.D(_01146_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[98] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_32_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[670]$_DFFE_PN0P_  (.D(_01147_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[702] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_40_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[671]$_DFFE_PN0P_  (.D(_01148_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[703] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_48_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[672]$_DFFE_PN0P_  (.D(_01149_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[704] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_54_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[673]$_DFFE_PN0P_  (.D(_01150_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[705] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_51_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[674]$_DFFE_PN0P_  (.D(_01151_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[706] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_58_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[675]$_DFFE_PN0P_  (.D(_01152_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[707] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_63_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[676]$_DFFE_PN0P_  (.D(_01153_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[708] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_83_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[677]$_DFFE_PN0P_  (.D(_01154_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[709] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[678]$_DFFE_PN0P_  (.D(_01155_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[710] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_93_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[679]$_DFFE_PN0P_  (.D(_01156_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[711] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_8_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[67]$_DFFE_PN0P_  (.D(_01157_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[99] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_38_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[680]$_DFFE_PN0P_  (.D(_01158_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[712] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[681]$_DFFE_PN0P_  (.D(_01159_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[713] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_72_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[682]$_DFFE_PN0P_  (.D(_01160_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[714] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_91_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[683]$_DFFE_PN0P_  (.D(_01161_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[715] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_93_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[684]$_DFFE_PN0P_  (.D(_01162_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[716] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_76_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[685]$_DFFE_PN0P_  (.D(_01163_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[717] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_58_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[686]$_DFFE_PN0P_  (.D(_01164_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[718] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_77_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[687]$_DFFE_PN0P_  (.D(_01165_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[719] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_59_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[688]$_DFFE_PN0P_  (.D(_01166_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[720] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[689]$_DFFE_PN0P_  (.D(_01167_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[721] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_54_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[68]$_DFFE_PN0P_  (.D(_01168_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[100] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_15_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[690]$_DFFE_PN0P_  (.D(_01169_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[722] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_75_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[691]$_DFFE_PN0P_  (.D(_01170_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[723] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[692]$_DFFE_PN0P_  (.D(_01171_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[724] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[693]$_DFFE_PN0P_  (.D(_01172_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[725] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_88_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[694]$_DFFE_PN0P_  (.D(_01173_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[726] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_7_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[695]$_DFFE_PN0P_  (.D(_01174_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[727] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_90_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[696]$_DFFE_PN0P_  (.D(_01175_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[728] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_79_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[697]$_DFFE_PN0P_  (.D(_01176_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[729] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[698]$_DFFE_PN0P_  (.D(_01177_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[730] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_90_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[699]$_DFFE_PN0P_  (.D(_01178_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[731] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[69]$_DFFE_PN0P_  (.D(_01179_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[101] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_13_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[6]$_DFFE_PN0P_  (.D(_01180_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[38] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_15_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[700]$_DFFE_PN0P_  (.D(_01181_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[732] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_78_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[701]$_DFFE_PN0P_  (.D(_01182_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[733] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_40_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[702]$_DFFE_PN0P_  (.D(_01183_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[734] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_39_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[703]$_DFFE_PN0P_  (.D(_01184_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[735] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_49_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[704]$_DFFE_PN0P_  (.D(_01185_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[736] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_55_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[705]$_DFFE_PN0P_  (.D(_01186_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[737] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_49_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[706]$_DFFE_PN0P_  (.D(_01187_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[738] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_60_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[707]$_DFFE_PN0P_  (.D(_01188_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[739] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_63_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[708]$_DFFE_PN0P_  (.D(_01189_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[740] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_83_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[709]$_DFFE_PN0P_  (.D(_01190_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[741] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[70]$_DFFE_PN0P_  (.D(_01191_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[102] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_15_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[710]$_DFFE_PN0P_  (.D(_01192_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[742] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_93_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[711]$_DFFE_PN0P_  (.D(_01193_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[743] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_8_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[712]$_DFFE_PN0P_  (.D(_01194_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[744] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[713]$_DFFE_PN0P_  (.D(_01195_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[745] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_71_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[714]$_DFFE_PN0P_  (.D(_01196_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[746] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_91_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[715]$_DFFE_PN0P_  (.D(_01197_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[747] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_92_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[716]$_DFFE_PN0P_  (.D(_01198_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[748] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_75_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[717]$_DFFE_PN0P_  (.D(_01199_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[749] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_58_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[718]$_DFFE_PN0P_  (.D(_01200_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[750] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_77_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[719]$_DFFE_PN0P_  (.D(_01201_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[751] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_59_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[71]$_DFFE_PN0P_  (.D(_01202_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[103] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_12_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[720]$_DFFE_PN0P_  (.D(_01203_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[752] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[721]$_DFFE_PN0P_  (.D(_01204_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[753] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_55_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[722]$_DFFE_PN0P_  (.D(_01205_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[754] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_74_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[723]$_DFFE_PN0P_  (.D(_01206_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[755] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[724]$_DFFE_PN0P_  (.D(_01207_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[756] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_8_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[725]$_DFFE_PN0P_  (.D(_01208_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[757] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[726]$_DFFE_PN0P_  (.D(_01209_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[758] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_7_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[727]$_DFFE_PN0P_  (.D(_01210_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[759] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_90_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[728]$_DFFE_PN0P_  (.D(_01211_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[760] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_79_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[729]$_DFFE_PN0P_  (.D(_01212_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[761] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[72]$_DFFE_PN0P_  (.D(_01213_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[104] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_37_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[730]$_DFFE_PN0P_  (.D(_01214_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[762] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_90_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[731]$_DFFE_PN0P_  (.D(_01215_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[763] ),
    .RESET_B(net469),
    .CLK(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[732]$_DFFE_PN0P_  (.D(_01216_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[764] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_78_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[733]$_DFFE_PN0P_  (.D(_01217_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[765] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_42_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[734]$_DFFE_PN0P_  (.D(_01218_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[766] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_41_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[735]$_DFFE_PN0P_  (.D(_01219_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[767] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_48_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[736]$_DFFE_PN0P_  (.D(_01220_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[768] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[737]$_DFFE_PN0P_  (.D(_01221_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[769] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_45_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[738]$_DFFE_PN0P_  (.D(_01222_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[770] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_44_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[739]$_DFFE_PN0P_  (.D(_01223_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[771] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_74_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[73]$_DFFE_PN0P_  (.D(_01224_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[105] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_28_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[740]$_DFFE_PN0P_  (.D(_01225_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[772] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_94_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[741]$_DFFE_PN0P_  (.D(_01226_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[773] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_3_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[742]$_DFFE_PN0P_  (.D(_01227_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[774] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_98_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[743]$_DFFE_PN0P_  (.D(_01228_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[775] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_5_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[744]$_DFFE_PN0P_  (.D(_01229_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[776] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_71_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[745]$_DFFE_PN0P_  (.D(_01230_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[777] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_74_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[746]$_DFFE_PN0P_  (.D(_01231_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[778] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_99_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[747]$_DFFE_PN0P_  (.D(_01232_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[779] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_6_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[748]$_DFFE_PN0P_  (.D(_01233_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[780] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[749]$_DFFE_PN0P_  (.D(_01234_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[781] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_45_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[74]$_DFFE_PN0P_  (.D(_01235_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[106] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_13_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[750]$_DFFE_PN0P_  (.D(_01236_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[782] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_4_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[751]$_DFFE_PN0P_  (.D(_01237_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[783] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_61_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[752]$_DFFE_PN0P_  (.D(_01238_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[784] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_46_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[753]$_DFFE_PN0P_  (.D(_01239_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[785] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_52_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[754]$_DFFE_PN0P_  (.D(_01240_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[786] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_70_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[755]$_DFFE_PN0P_  (.D(_01241_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[787] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_44_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[756]$_DFFE_PN0P_  (.D(_01242_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[788] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_4_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[757]$_DFFE_PN0P_  (.D(_01243_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[789] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[758]$_DFFE_PN0P_  (.D(_01244_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[790] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_6_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[759]$_DFFE_PN0P_  (.D(_01245_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[791] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_94_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[75]$_DFFE_PN0P_  (.D(_01246_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[107] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_14_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[760]$_DFFE_PN0P_  (.D(_01247_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[792] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_11_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[761]$_DFFE_PN0P_  (.D(_01248_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[793] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[762]$_DFFE_PN0P_  (.D(_01249_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[794] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[763]$_DFFE_PN0P_  (.D(_01250_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[795] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[764]$_DFFE_PN0P_  (.D(_01251_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[796] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_77_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[765]$_DFFE_PN0P_  (.D(_01252_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[797] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_40_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[766]$_DFFE_PN0P_  (.D(_01253_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[798] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_71_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[767]$_DFFE_PN0P_  (.D(_01254_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[799] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_46_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[768]$_DFFE_PN0P_  (.D(_01255_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[800] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_41_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[769]$_DFFE_PN0P_  (.D(_01256_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[801] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_45_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[76]$_DFFE_PN0P_  (.D(_01257_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[108] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_29_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[770]$_DFFE_PN0P_  (.D(_01258_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[802] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_44_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[771]$_DFFE_PN0P_  (.D(_01259_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[803] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_74_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[772]$_DFFE_PN0P_  (.D(_01260_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[804] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_7_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[773]$_DFFE_PN0P_  (.D(_01261_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[805] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_3_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[774]$_DFFE_PN0P_  (.D(_01262_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[806] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_98_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[775]$_DFFE_PN0P_  (.D(_01263_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[807] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_3_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[776]$_DFFE_PN0P_  (.D(_01264_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[808] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_71_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[777]$_DFFE_PN0P_  (.D(_01265_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[809] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_73_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[778]$_DFFE_PN0P_  (.D(_01266_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[810] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[779]$_DFFE_PN0P_  (.D(_01267_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[811] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_5_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[77]$_DFFE_PN0P_  (.D(_01268_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[109] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_35_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[780]$_DFFE_PN0P_  (.D(_01269_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[812] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[781]$_DFFE_PN0P_  (.D(_01270_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[813] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_43_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[782]$_DFFE_PN0P_  (.D(_01271_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[814] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_4_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[783]$_DFFE_PN0P_  (.D(_01272_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[815] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[784]$_DFFE_PN0P_  (.D(_01273_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[816] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[785]$_DFFE_PN0P_  (.D(_01274_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[817] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[786]$_DFFE_PN0P_  (.D(_01275_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[818] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_75_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[787]$_DFFE_PN0P_  (.D(_01276_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[819] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_73_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[788]$_DFFE_PN0P_  (.D(_01277_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[820] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_5_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[789]$_DFFE_PN0P_  (.D(_01278_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[821] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_85_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[78]$_DFFE_PN0P_  (.D(_01279_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[110] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_12_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[790]$_DFFE_PN0P_  (.D(_01280_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[822] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[791]$_DFFE_PN0P_  (.D(_01281_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[823] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_98_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[792]$_DFFE_PN0P_  (.D(_01282_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[824] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_11_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[793]$_DFFE_PN0P_  (.D(_01283_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[825] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_85_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[794]$_DFFE_PN0P_  (.D(_01284_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[826] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[795]$_DFFE_PN0P_  (.D(_01285_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[827] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_85_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[796]$_DFFE_PN0P_  (.D(_01286_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[828] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_78_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[797]$_DFFE_PN0P_  (.D(_01287_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[829] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_39_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[798]$_DFFE_PN0P_  (.D(_01288_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[830] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_71_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[799]$_DFFE_PN0P_  (.D(_01289_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[831] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_46_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[79]$_DFFE_PN0P_  (.D(_01290_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[111] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_33_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[7]$_DFFE_PN0P_  (.D(_01291_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[39] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_13_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[800]$_DFFE_PN0P_  (.D(_01292_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[832] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_42_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[801]$_DFFE_PN0P_  (.D(_01293_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[833] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_44_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[802]$_DFFE_PN0P_  (.D(_01294_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[834] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_43_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[803]$_DFFE_PN0P_  (.D(_01295_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[835] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_76_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[804]$_DFFE_PN0P_  (.D(_01296_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[836] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_83_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[805]$_DFFE_PN0P_  (.D(_01297_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[837] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_3_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[806]$_DFFE_PN0P_  (.D(_01298_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[838] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_97_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[807]$_DFFE_PN0P_  (.D(_01299_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[839] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_3_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[808]$_DFFE_PN0P_  (.D(_01300_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[840] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_71_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[809]$_DFFE_PN0P_  (.D(_01301_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[841] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_74_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[80]$_DFFE_PN0P_  (.D(_01302_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[112] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_31_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[810]$_DFFE_PN0P_  (.D(_01303_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[842] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[811]$_DFFE_PN0P_  (.D(_01304_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[843] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_6_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[812]$_DFFE_PN0P_  (.D(_01305_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[844] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_82_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[813]$_DFFE_PN0P_  (.D(_01306_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[845] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_43_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[814]$_DFFE_PN0P_  (.D(_01307_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[846] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_4_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[815]$_DFFE_PN0P_  (.D(_01308_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[847] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[816]$_DFFE_PN0P_  (.D(_01309_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[848] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[817]$_DFFE_PN0P_  (.D(_01310_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[849] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_44_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[818]$_DFFE_PN0P_  (.D(_01311_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[850] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_70_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[819]$_DFFE_PN0P_  (.D(_01312_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[851] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_44_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[81]$_DFFE_PN0P_  (.D(_01313_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[113] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_35_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[820]$_DFFE_PN0P_  (.D(_01314_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[852] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_5_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[821]$_DFFE_PN0P_  (.D(_01315_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[853] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[822]$_DFFE_PN0P_  (.D(_01316_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[854] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[823]$_DFFE_PN0P_  (.D(_01317_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[855] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_94_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[824]$_DFFE_PN0P_  (.D(_01318_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[856] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_11_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[825]$_DFFE_PN0P_  (.D(_01319_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[857] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_80_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[826]$_DFFE_PN0P_  (.D(_01320_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[858] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[827]$_DFFE_PN0P_  (.D(_01321_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[859] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_85_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[828]$_DFFE_PN0P_  (.D(_01322_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[860] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_78_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[829]$_DFFE_PN0P_  (.D(_01323_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[861] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_40_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[82]$_DFFE_PN0P_  (.D(_01324_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[114] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_27_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[830]$_DFFE_PN0P_  (.D(_01325_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[862] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_69_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[831]$_DFFE_PN0P_  (.D(_01326_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[863] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_46_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[832]$_DFFE_PN0P_  (.D(_01327_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[864] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_41_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[833]$_DFFE_PN0P_  (.D(_01328_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[865] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_46_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[834]$_DFFE_PN0P_  (.D(_01329_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[866] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_44_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[835]$_DFFE_PN0P_  (.D(_01330_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[867] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_76_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[836]$_DFFE_PN0P_  (.D(_01331_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[868] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_7_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[837]$_DFFE_PN0P_  (.D(_01332_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[869] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_3_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[838]$_DFFE_PN0P_  (.D(_01333_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[870] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_98_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[839]$_DFFE_PN0P_  (.D(_01334_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[871] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_3_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[83]$_DFFE_PN0P_  (.D(_01335_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[115] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_36_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[840]$_DFFE_PN0P_  (.D(_01336_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[872] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_71_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[841]$_DFFE_PN0P_  (.D(_01337_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[873] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_74_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[842]$_DFFE_PN0P_  (.D(_01338_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[874] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[843]$_DFFE_PN0P_  (.D(_01339_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[875] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_6_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[844]$_DFFE_PN0P_  (.D(_01340_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[876] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_82_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[845]$_DFFE_PN0P_  (.D(_01341_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[877] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_42_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[846]$_DFFE_PN0P_  (.D(_01342_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[878] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_4_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[847]$_DFFE_PN0P_  (.D(_01343_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[879] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[848]$_DFFE_PN0P_  (.D(_01344_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[880] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_46_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[849]$_DFFE_PN0P_  (.D(_01345_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[881] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_52_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[84]$_DFFE_PN0P_  (.D(_01346_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[116] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_15_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[850]$_DFFE_PN0P_  (.D(_01347_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[882] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_70_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[851]$_DFFE_PN0P_  (.D(_01348_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[883] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_73_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[852]$_DFFE_PN0P_  (.D(_01349_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[884] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_5_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[853]$_DFFE_PN0P_  (.D(_01350_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[885] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_85_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[854]$_DFFE_PN0P_  (.D(_01351_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[886] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[855]$_DFFE_PN0P_  (.D(_01352_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[887] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_94_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[856]$_DFFE_PN0P_  (.D(_01353_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[888] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_11_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[857]$_DFFE_PN0P_  (.D(_01354_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[889] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[858]$_DFFE_PN0P_  (.D(_01355_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[890] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_83_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[859]$_DFFE_PN0P_  (.D(_01356_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[891] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_85_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[85]$_DFFE_PN0P_  (.D(_01357_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[117] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_25_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[860]$_DFFE_PN0P_  (.D(_01358_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[892] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_79_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[861]$_DFFE_PN0P_  (.D(_01359_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[893] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_40_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[862]$_DFFE_PN0P_  (.D(_01360_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[894] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_71_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[863]$_DFFE_PN0P_  (.D(_01361_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[895] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_46_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[864]$_DFFE_PN0P_  (.D(_01362_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[896] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[865]$_DFFE_PN0P_  (.D(_01363_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[897] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_45_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[866]$_DFFE_PN0P_  (.D(_01364_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[898] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_44_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[867]$_DFFE_PN0P_  (.D(_01365_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[899] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_76_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[868]$_DFFE_PN0P_  (.D(_01366_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[900] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_83_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[869]$_DFFE_PN0P_  (.D(_01367_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[901] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_3_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[86]$_DFFE_PN0P_  (.D(_01368_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[118] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_15_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[870]$_DFFE_PN0P_  (.D(_01369_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[902] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_97_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[871]$_DFFE_PN0P_  (.D(_01370_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[903] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[872]$_DFFE_PN0P_  (.D(_01371_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[904] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_71_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[873]$_DFFE_PN0P_  (.D(_01372_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[905] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_43_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[874]$_DFFE_PN0P_  (.D(_01373_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[906] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_1_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[875]$_DFFE_PN0P_  (.D(_01374_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[907] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_7_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[876]$_DFFE_PN0P_  (.D(_01375_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[908] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[877]$_DFFE_PN0P_  (.D(_01376_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[909] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_42_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[878]$_DFFE_PN0P_  (.D(_01377_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[910] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[879]$_DFFE_PN0P_  (.D(_01378_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[911] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_61_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[87]$_DFFE_PN0P_  (.D(_01379_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[119] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_23_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[880]$_DFFE_PN0P_  (.D(_01380_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[912] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_48_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[881]$_DFFE_PN0P_  (.D(_01381_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[913] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_52_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[882]$_DFFE_PN0P_  (.D(_01382_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[914] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_71_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[883]$_DFFE_PN0P_  (.D(_01383_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[915] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[884]$_DFFE_PN0P_  (.D(_01384_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[916] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_5_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[885]$_DFFE_PN0P_  (.D(_01385_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[917] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[886]$_DFFE_PN0P_  (.D(_01386_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[918] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[887]$_DFFE_PN0P_  (.D(_01387_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[919] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_93_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[888]$_DFFE_PN0P_  (.D(_01388_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[920] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_10_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[889]$_DFFE_PN0P_  (.D(_01389_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[921] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[88]$_DFFE_PN0P_  (.D(_01390_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[120] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_26_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[890]$_DFFE_PN0P_  (.D(_01391_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[922] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[891]$_DFFE_PN0P_  (.D(_01392_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[923] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_85_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[892]$_DFFE_PN0P_  (.D(_01393_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[924] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_12_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[893]$_DFFE_PN0P_  (.D(_01394_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[925] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_42_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[894]$_DFFE_PN0P_  (.D(_01395_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[926] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_69_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[895]$_DFFE_PN0P_  (.D(_01396_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[927] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_46_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[896]$_DFFE_PN0P_  (.D(_01397_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[928] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_32_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[897]$_DFFE_PN0P_  (.D(_01398_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[929] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_45_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[898]$_DFFE_PN0P_  (.D(_01399_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[930] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_44_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[899]$_DFFE_PN0P_  (.D(_01400_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[931] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_77_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[89]$_DFFE_PN0P_  (.D(_01401_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[121] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_27_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[8]$_DFFE_PN0P_  (.D(_01402_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[40] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_37_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[900]$_DFFE_PN0P_  (.D(_01403_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[932] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_83_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[901]$_DFFE_PN0P_  (.D(_01404_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[933] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[902]$_DFFE_PN0P_  (.D(_01405_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[934] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_97_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[903]$_DFFE_PN0P_  (.D(_01406_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[935] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[904]$_DFFE_PN0P_  (.D(_01407_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[936] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_63_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[905]$_DFFE_PN0P_  (.D(_01408_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[937] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_74_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[906]$_DFFE_PN0P_  (.D(_01409_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[938] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[907]$_DFFE_PN0P_  (.D(_01410_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[939] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_6_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[908]$_DFFE_PN0P_  (.D(_01411_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[940] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_82_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[909]$_DFFE_PN0P_  (.D(_01412_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[941] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_42_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[90]$_DFFE_PN0P_  (.D(_01413_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[122] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_13_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[910]$_DFFE_PN0P_  (.D(_01414_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[942] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_20_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[911]$_DFFE_PN0P_  (.D(_01415_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[943] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_60_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[912]$_DFFE_PN0P_  (.D(_01416_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[944] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[913]$_DFFE_PN0P_  (.D(_01417_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[945] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_52_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[914]$_DFFE_PN0P_  (.D(_01418_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[946] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_70_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[915]$_DFFE_PN0P_  (.D(_01419_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[947] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_72_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[916]$_DFFE_PN0P_  (.D(_01420_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[948] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_6_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[917]$_DFFE_PN0P_  (.D(_01421_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[949] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[918]$_DFFE_PN0P_  (.D(_01422_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[950] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[919]$_DFFE_PN0P_  (.D(_01423_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[951] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_94_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[91]$_DFFE_PN0P_  (.D(_01424_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[123] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_26_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[920]$_DFFE_PN0P_  (.D(_01425_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[952] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_10_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[921]$_DFFE_PN0P_  (.D(_01426_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[953] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[922]$_DFFE_PN0P_  (.D(_01427_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[954] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[923]$_DFFE_PN0P_  (.D(_01428_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[955] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_85_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[924]$_DFFE_PN0P_  (.D(_01429_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[956] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_11_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[925]$_DFFE_PN0P_  (.D(_01430_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[957] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_43_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[926]$_DFFE_PN0P_  (.D(_01431_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[958] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[927]$_DFFE_PN0P_  (.D(_01432_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[959] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_42_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[928]$_DFFE_PN0P_  (.D(_01433_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[960] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[929]$_DFFE_PN0P_  (.D(_01434_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[961] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_51_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[92]$_DFFE_PN0P_  (.D(_01435_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[124] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_25_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[930]$_DFFE_PN0P_  (.D(_01436_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[962] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_44_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[931]$_DFFE_PN0P_  (.D(_01437_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[963] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_77_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[932]$_DFFE_PN0P_  (.D(_01438_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[964] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_83_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[933]$_DFFE_PN0P_  (.D(_01439_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[965] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[934]$_DFFE_PN0P_  (.D(_01440_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[966] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_97_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[935]$_DFFE_PN0P_  (.D(_01441_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[967] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[936]$_DFFE_PN0P_  (.D(_01442_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[968] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_71_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[937]$_DFFE_PN0P_  (.D(_01443_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[969] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_40_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[938]$_DFFE_PN0P_  (.D(_01444_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[970] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_1_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[939]$_DFFE_PN0P_  (.D(_01445_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[971] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_6_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[93]$_DFFE_PN0P_  (.D(_01446_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[125] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_37_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[940]$_DFFE_PN0P_  (.D(_01447_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[972] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[941]$_DFFE_PN0P_  (.D(_01448_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[973] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_42_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[942]$_DFFE_PN0P_  (.D(_01449_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[974] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[943]$_DFFE_PN0P_  (.D(_01450_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[975] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_61_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[944]$_DFFE_PN0P_  (.D(_01451_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[976] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[945]$_DFFE_PN0P_  (.D(_01452_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[977] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[946]$_DFFE_PN0P_  (.D(_01453_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[978] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_69_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[947]$_DFFE_PN0P_  (.D(_01454_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[979] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_73_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[948]$_DFFE_PN0P_  (.D(_01455_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[980] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_5_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[949]$_DFFE_PN0P_  (.D(_01456_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[981] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[94]$_DFFE_PN0P_  (.D(_01457_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[126] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_37_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[950]$_DFFE_PN0P_  (.D(_01458_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[982] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[951]$_DFFE_PN0P_  (.D(_01459_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[983] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_95_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[952]$_DFFE_PN0P_  (.D(_01460_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[984] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_10_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[953]$_DFFE_PN0P_  (.D(_01461_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[985] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_70_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[954]$_DFFE_PN0P_  (.D(_01462_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[986] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[955]$_DFFE_PN0P_  (.D(_01463_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[987] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_83_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[956]$_DFFE_PN0P_  (.D(_01464_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[988] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_78_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[957]$_DFFE_PN0P_  (.D(_01465_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[989] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_40_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[958]$_DFFE_PN0P_  (.D(_01466_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[990] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_69_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[959]$_DFFE_PN0P_  (.D(_01467_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[991] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[95]$_DFFE_PN0P_  (.D(_01468_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[127] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_33_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[960]$_DFFE_PN0P_  (.D(_01469_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[992] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[961]$_DFFE_PN0P_  (.D(_01470_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[993] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_45_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[962]$_DFFE_PN0P_  (.D(_01471_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[994] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_45_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[963]$_DFFE_PN0P_  (.D(_01472_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[995] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_77_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[964]$_DFFE_PN0P_  (.D(_01473_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[996] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_82_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[965]$_DFFE_PN0P_  (.D(_01474_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[997] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[966]$_DFFE_PN0P_  (.D(_01475_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[998] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_97_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[967]$_DFFE_PN0P_  (.D(_01476_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[999] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[968]$_DFFE_PN0P_  (.D(_01477_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1000] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_71_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[969]$_DFFE_PN0P_  (.D(_01478_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1001] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_77_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[96]$_DFFE_PN0P_  (.D(_01479_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[128] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_32_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[970]$_DFFE_PN0P_  (.D(_01480_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1002] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_1_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[971]$_DFFE_PN0P_  (.D(_01481_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1003] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_6_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[972]$_DFFE_PN0P_  (.D(_01482_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1004] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_82_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[973]$_DFFE_PN0P_  (.D(_01483_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1005] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_42_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[974]$_DFFE_PN0P_  (.D(_01484_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1006] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_20_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[975]$_DFFE_PN0P_  (.D(_01485_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1007] ),
    .RESET_B(net468),
    .CLK(clknet_leaf_61_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[976]$_DFFE_PN0P_  (.D(_01486_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1008] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_31_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[977]$_DFFE_PN0P_  (.D(_01487_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1009] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_52_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[978]$_DFFE_PN0P_  (.D(_01488_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1010] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_70_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[979]$_DFFE_PN0P_  (.D(_01489_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1011] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_73_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[97]$_DFFE_PN0P_  (.D(_01490_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[129] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_30_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[980]$_DFFE_PN0P_  (.D(_01491_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1012] ),
    .RESET_B(net458),
    .CLK(clknet_leaf_5_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[981]$_DFFE_PN0P_  (.D(_01492_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1013] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[982]$_DFFE_PN0P_  (.D(_01493_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1014] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_1_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[983]$_DFFE_PN0P_  (.D(_01494_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1015] ),
    .RESET_B(net466),
    .CLK(clknet_leaf_95_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[984]$_DFFE_PN0P_  (.D(_01495_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1016] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_8_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[985]$_DFFE_PN0P_  (.D(_01496_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1017] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[986]$_DFFE_PN0P_  (.D(_01497_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1018] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_93_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[987]$_DFFE_PN0P_  (.D(_01498_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1019] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_83_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[988]$_DFFE_PN0P_  (.D(_01499_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1020] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_78_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[989]$_DFFE_PN0P_  (.D(_01500_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1021] ),
    .RESET_B(net465),
    .CLK(clknet_leaf_40_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[98]$_DFFE_PN0P_  (.D(_01501_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[130] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_41_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[990]$_DFFE_PN0P_  (.D(_01502_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1022] ),
    .RESET_B(net467),
    .CLK(clknet_leaf_69_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[991]$_DFFE_PN0P_  (.D(_01503_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[1023] ),
    .RESET_B(net464),
    .CLK(clknet_leaf_46_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[99]$_DFFE_PN0P_  (.D(_01504_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[131] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_38_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_1 \gen_regfile_ff.register_file_i.rf_reg_q[9]$_DFFE_PN0P_  (.D(_01505_),
    .Q(\gen_regfile_ff.register_file_i.rf_reg[41] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_37_clk_i_regs));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.controller_i.ctrl_fsm_cs[0]$_DFFE_PN0P_  (.D(_01506_),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs[0] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.controller_i.ctrl_fsm_cs[1]$_DFFE_PN0P_  (.D(_01507_),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs[1] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.controller_i.ctrl_fsm_cs[2]$_DFFE_PN0P_  (.D(_01508_),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs[2] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.controller_i.ctrl_fsm_cs[3]$_DFFE_PN0P_  (.D(_01509_),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs[3] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.controller_i.debug_mode_q$_DFFE_PN0P_  (.D(_01510_),
    .Q(\cs_registers_i.debug_mode_i ),
    .RESET_B(net455),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.controller_i.exc_req_q$_DFF_PN0_  (.D(\id_stage_i.controller_i.exc_req_d ),
    .Q(\id_stage_i.controller_i.exc_req_q ),
    .RESET_B(net455),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.controller_i.illegal_insn_q$_DFF_PN0_  (.D(\id_stage_i.controller_i.illegal_insn_d ),
    .Q(\id_stage_i.controller_i.illegal_insn_q ),
    .RESET_B(net455),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.controller_i.load_err_q$_DFF_PN0_  (.D(\id_stage_i.controller_i.load_err_d ),
    .Q(\id_stage_i.controller_i.load_err_q ),
    .RESET_B(net455),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_2 \id_stage_i.controller_i.nmi_mode_q$_DFFE_PN0P_  (.D(_01511_),
    .Q(\cs_registers_i.nmi_mode_i ),
    .RESET_B(net452),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.controller_i.store_err_q$_DFF_PN0_  (.D(\id_stage_i.controller_i.store_err_d ),
    .Q(\id_stage_i.controller_i.store_err_q ),
    .RESET_B(net455),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.g_branch_set_flop.branch_set_q$_DFF_PN0_  (.D(\id_stage_i.branch_set_d ),
    .Q(\id_stage_i.branch_set ),
    .RESET_B(net456),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.id_fsm_q$_DFFE_PN0P_  (.D(_01512_),
    .Q(\id_stage_i.id_fsm_q ),
    .RESET_B(net456),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[0]$_DFFE_PN0P_  (.D(_01513_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[0] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[10]$_DFFE_PN0P_  (.D(_01514_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[10] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[11]$_DFFE_PN0P_  (.D(_01515_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[11] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[12]$_DFFE_PN0P_  (.D(_01516_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[12] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[13]$_DFFE_PN0P_  (.D(_01517_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[13] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[14]$_DFFE_PN0P_  (.D(_01518_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[14] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[15]$_DFFE_PN0P_  (.D(_01519_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[15] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[16]$_DFFE_PN0P_  (.D(_01520_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[16] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[17]$_DFFE_PN0P_  (.D(_01521_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[17] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[18]$_DFFE_PN0P_  (.D(_01522_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[18] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[19]$_DFFE_PN0P_  (.D(_01523_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[19] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[1]$_DFFE_PN0P_  (.D(_01524_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[1] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[20]$_DFFE_PN0P_  (.D(_01525_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[20] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[21]$_DFFE_PN0P_  (.D(_01526_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[21] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[22]$_DFFE_PN0P_  (.D(_01527_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[22] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[23]$_DFFE_PN0P_  (.D(_01528_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[23] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[24]$_DFFE_PN0P_  (.D(_01529_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[24] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[25]$_DFFE_PN0P_  (.D(_01530_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[25] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[26]$_DFFE_PN0P_  (.D(_01531_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[26] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[27]$_DFFE_PN0P_  (.D(_01532_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[27] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[28]$_DFFE_PN0P_  (.D(_01533_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[28] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[29]$_DFFE_PN0P_  (.D(_01534_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[29] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[2]$_DFFE_PN0P_  (.D(_01535_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[2] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[30]$_DFFE_PN0P_  (.D(_01536_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[30] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[31]$_DFFE_PN0P_  (.D(_01537_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[31] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[34]$_DFFE_PN0P_  (.D(_01538_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[32] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[35]$_DFFE_PN0P_  (.D(_01539_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[33] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[36]$_DFFE_PN0P_  (.D(_01540_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[34] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[37]$_DFFE_PN0P_  (.D(_01541_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[35] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[38]$_DFFE_PN0P_  (.D(_01542_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[36] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[39]$_DFFE_PN0P_  (.D(_01543_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[37] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[3]$_DFFE_PN0P_  (.D(_01544_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[3] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[40]$_DFFE_PN0P_  (.D(_01545_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[38] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[41]$_DFFE_PN0P_  (.D(_01546_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[39] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[42]$_DFFE_PN0P_  (.D(_01547_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[40] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[43]$_DFFE_PN0P_  (.D(_01548_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[41] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[44]$_DFFE_PN0P_  (.D(_01549_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[42] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[45]$_DFFE_PN0P_  (.D(_01550_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[43] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[46]$_DFFE_PN0P_  (.D(_01551_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[44] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[47]$_DFFE_PN0P_  (.D(_01552_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[45] ),
    .RESET_B(net463),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[48]$_DFFE_PN0P_  (.D(_01553_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[46] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[49]$_DFFE_PN0P_  (.D(_01554_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[47] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[4]$_DFFE_PN0P_  (.D(_01555_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[4] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[50]$_DFFE_PN0P_  (.D(_01556_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[48] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[51]$_DFFE_PN0P_  (.D(_01557_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[49] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[52]$_DFFE_PN0P_  (.D(_01558_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[50] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[53]$_DFFE_PN0P_  (.D(_01559_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[51] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[54]$_DFFE_PN0P_  (.D(_01560_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[52] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[55]$_DFFE_PN0P_  (.D(_01561_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[53] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[56]$_DFFE_PN0P_  (.D(_01562_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[54] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[57]$_DFFE_PN0P_  (.D(_01563_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[55] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[58]$_DFFE_PN0P_  (.D(_01564_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[56] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[59]$_DFFE_PN0P_  (.D(_01565_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[57] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[5]$_DFFE_PN0P_  (.D(_01566_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[5] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[60]$_DFFE_PN0P_  (.D(_01567_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[58] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[61]$_DFFE_PN0P_  (.D(_01568_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[59] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[62]$_DFFE_PN0P_  (.D(_01569_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[60] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[63]$_DFFE_PN0P_  (.D(_01570_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[61] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[64]$_DFFE_PN0P_  (.D(_01571_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[62] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfrtp_4 \id_stage_i.imd_val_q[65]$_DFFE_PN0P_  (.D(_01572_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[63] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfrtp_2 \id_stage_i.imd_val_q[66]$_DFFE_PN0P_  (.D(_01573_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[66] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfrtp_2 \id_stage_i.imd_val_q[67]$_DFFE_PN0P_  (.D(_01574_),
    .Q(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.imd_val_q_i[67] ),
    .RESET_B(net462),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[6]$_DFFE_PN0P_  (.D(_01575_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[6] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[7]$_DFFE_PN0P_  (.D(_01576_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[7] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[8]$_DFFE_PN0P_  (.D(_01577_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[8] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfrtp_1 \id_stage_i.imd_val_q[9]$_DFFE_PN0P_  (.D(_01578_),
    .Q(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[9] ),
    .RESET_B(net459),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__dfrtp_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfrtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_q ),
    .RESET_B(net455),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[10] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[11] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[12] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[13] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[14] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[15] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[16] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[17] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[18] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[19] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[20] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[21] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[22] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[23] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[24] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[25] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[26] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[27] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[28] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[29] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[2] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[30] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[31] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[3] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[4] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[5] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[6] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[7] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[8] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[9] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_d[0] ),
    .DE(net1061),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_d[1] ),
    .DE(net990),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2]$_DFFE_PP_  (.D(net94),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[2] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[0]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[1] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(\cs_registers_i.pc_if_i[1] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[10]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[11] ),
    .DE(net254),
    .Q(\cs_registers_i.pc_if_i[11] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[11]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[12] ),
    .DE(net254),
    .Q(\cs_registers_i.pc_if_i[12] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[12]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[13] ),
    .DE(net254),
    .Q(\cs_registers_i.pc_if_i[13] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[13]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[14] ),
    .DE(net254),
    .Q(\cs_registers_i.pc_if_i[14] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[14]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[15] ),
    .DE(net254),
    .Q(\cs_registers_i.pc_if_i[15] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[15]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[16] ),
    .DE(net254),
    .Q(\cs_registers_i.pc_if_i[16] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[16]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[17] ),
    .DE(net254),
    .Q(\cs_registers_i.pc_if_i[17] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[17]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[18] ),
    .DE(net254),
    .Q(\cs_registers_i.pc_if_i[18] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[18]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[19] ),
    .DE(net254),
    .Q(\cs_registers_i.pc_if_i[19] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[19]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[20] ),
    .DE(net254),
    .Q(\cs_registers_i.pc_if_i[20] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[1]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[2] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(\cs_registers_i.pc_if_i[2] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[20]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[21] ),
    .DE(net254),
    .Q(\cs_registers_i.pc_if_i[21] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[21]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[22] ),
    .DE(net254),
    .Q(\cs_registers_i.pc_if_i[22] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[22]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[23] ),
    .DE(net254),
    .Q(\cs_registers_i.pc_if_i[23] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[23]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[24] ),
    .DE(net254),
    .Q(\cs_registers_i.pc_if_i[24] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[24]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[25] ),
    .DE(net254),
    .Q(\cs_registers_i.pc_if_i[25] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[25]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[26] ),
    .DE(net254),
    .Q(\cs_registers_i.pc_if_i[26] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[26]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[27] ),
    .DE(net254),
    .Q(\cs_registers_i.pc_if_i[27] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[27]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[28] ),
    .DE(net254),
    .Q(\cs_registers_i.pc_if_i[28] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[28]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[29] ),
    .DE(net254),
    .Q(\cs_registers_i.pc_if_i[29] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[29]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[30] ),
    .DE(net254),
    .Q(\cs_registers_i.pc_if_i[30] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[2]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[3] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(\cs_registers_i.pc_if_i[3] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[30]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[31] ),
    .DE(net254),
    .Q(\cs_registers_i.pc_if_i[31] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[3]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[4] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(\cs_registers_i.pc_if_i[4] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[4]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[5] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(\cs_registers_i.pc_if_i[5] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[5]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[6] ),
    .DE(net254),
    .Q(\cs_registers_i.pc_if_i[6] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[6]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[7] ),
    .DE(net254),
    .Q(\cs_registers_i.pc_if_i[7] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[7]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[8] ),
    .DE(net254),
    .Q(\cs_registers_i.pc_if_i[8] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[8]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[9] ),
    .DE(net254),
    .Q(\cs_registers_i.pc_if_i[9] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[9]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[10] ),
    .DE(net254),
    .Q(\cs_registers_i.pc_if_i[10] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[0] ),
    .DE(net1061),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[10] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[11] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[12] ),
    .DE(net1305),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[13] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[14] ),
    .DE(net1305),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[15] ),
    .DE(net1061),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[16] ),
    .DE(net1305),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[17] ),
    .DE(net1305),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[18] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[19] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[1] ),
    .DE(net1061),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[20] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[21] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[22] ),
    .DE(net1305),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[23] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[24] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[25] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[26] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[27] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[28] ),
    .DE(net1061),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[29] ),
    .DE(net1061),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[2] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[30] ),
    .DE(net1061),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[31] ),
    .DE(net1061),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[32] ),
    .DE(net990),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[33] ),
    .DE(net1039),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[34] ),
    .DE(net990),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[35] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[36] ),
    .DE(net1039),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[37] ),
    .DE(net1039),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[38] ),
    .DE(net1303),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[39] ),
    .DE(net1303),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[3] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[40] ),
    .DE(net990),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[41] ),
    .DE(net1039),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[42] ),
    .DE(net1039),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[43] ),
    .DE(net1303),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[44] ),
    .DE(net1303),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[45] ),
    .DE(net1460),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[46] ),
    .DE(net1039),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[47] ),
    .DE(net990),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[48] ),
    .DE(net1303),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[49] ),
    .DE(net1303),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[4] ),
    .DE(net1305),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[50] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[51] ),
    .DE(net1460),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[52] ),
    .DE(net1460),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[53] ),
    .DE(net990),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[54] ),
    .DE(net1303),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[55] ),
    .DE(net990),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[56] ),
    .DE(net990),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[57] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[58] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[59] ),
    .DE(net1039),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[5] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[60] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[61] ),
    .DE(net1460),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[62] ),
    .DE(net1039),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[63] ),
    .DE(net1303),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64]$_DFFE_PP_  (.D(net96),
    .DE(net317),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65]$_DFFE_PP_  (.D(net107),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[2] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66]$_DFFE_PP_  (.D(net118),
    .DE(net317),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67]$_DFFE_PP_  (.D(net121),
    .DE(net317),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68]$_DFFE_PP_  (.D(net122),
    .DE(net317),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69]$_DFFE_PP_  (.D(net123),
    .DE(net317),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[6] ),
    .DE(net1305),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70]$_DFFE_PP_  (.D(net124),
    .DE(net317),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71]$_DFFE_PP_  (.D(net125),
    .DE(net317),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72]$_DFFE_PP_  (.D(net126),
    .DE(net317),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73]$_DFFE_PP_  (.D(net127),
    .DE(net317),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74]$_DFFE_PP_  (.D(net97),
    .DE(net317),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75]$_DFFE_PP_  (.D(net98),
    .DE(net317),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76]$_DFFE_PP_  (.D(net99),
    .DE(net318),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77]$_DFFE_PP_  (.D(net100),
    .DE(net318),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78]$_DFFE_PP_  (.D(net101),
    .DE(net317),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79]$_DFFE_PP_  (.D(net102),
    .DE(net317),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[7] ),
    .DE(net1305),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80]$_DFFE_PP_  (.D(net103),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[2] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81]$_DFFE_PP_  (.D(net104),
    .DE(net318),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82]$_DFFE_PP_  (.D(net105),
    .DE(net318),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83]$_DFFE_PP_  (.D(net106),
    .DE(net318),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84]$_DFFE_PP_  (.D(net108),
    .DE(net318),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85]$_DFFE_PP_  (.D(net109),
    .DE(net318),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86]$_DFFE_PP_  (.D(net110),
    .DE(net317),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87]$_DFFE_PP_  (.D(net111),
    .DE(net318),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88]$_DFFE_PP_  (.D(net112),
    .DE(net318),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89]$_DFFE_PP_  (.D(net113),
    .DE(net318),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[8] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90]$_DFFE_PP_  (.D(net114),
    .DE(net318),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91]$_DFFE_PP_  (.D(net115),
    .DE(net318),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92]$_DFFE_PP_  (.D(net116),
    .DE(net318),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93]$_DFFE_PP_  (.D(net117),
    .DE(net318),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94]$_DFFE_PP_  (.D(net119),
    .DE(net318),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95]$_DFFE_PP_  (.D(net120),
    .DE(net318),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9]$_DFFE_PP_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[9] ),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfrtp_4 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_4 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[1]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_4 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[2]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfrtp_2 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1]$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10]$_DFFE_PP_  (.D(net219),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11]$_DFFE_PP_  (.D(net220),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12]$_DFFE_PP_  (.D(net221),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13]$_DFFE_PP_  (.D(net222),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14]$_DFFE_PP_  (.D(net223),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15]$_DFFE_PP_  (.D(net224),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16]$_DFFE_PP_  (.D(net225),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17]$_DFFE_PP_  (.D(net226),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18]$_DFFE_PP_  (.D(net227),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19]$_DFFE_PP_  (.D(net228),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20]$_DFFE_PP_  (.D(net229),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21]$_DFFE_PP_  (.D(net230),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22]$_DFFE_PP_  (.D(net231),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23]$_DFFE_PP_  (.D(net232),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24]$_DFFE_PP_  (.D(net233),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25]$_DFFE_PP_  (.D(net234),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26]$_DFFE_PP_  (.D(net235),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27]$_DFFE_PP_  (.D(net236),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28]$_DFFE_PP_  (.D(net237),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29]$_DFFE_PP_  (.D(net238),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2]$_DFFE_PP_  (.D(net239),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30]$_DFFE_PP_  (.D(net240),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31]$_DFFE_PP_  (.D(net241),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3]$_DFFE_PP_  (.D(net242),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4]$_DFFE_PP_  (.D(net243),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5]$_DFFE_PP_  (.D(net244),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6]$_DFFE_PP_  (.D(net245),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7]$_DFFE_PP_  (.D(net246),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8]$_DFFE_PP_  (.D(net247),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9]$_DFFE_PP_  (.D(net248),
    .DE(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfrtp_4 \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q$_DFF_PN0_  (.D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ),
    .Q(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .RESET_B(net455),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.illegal_c_insn_id_o$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.illegal_instr_o ),
    .DE(net253),
    .Q(\id_stage_i.decoder_i.illegal_c_insn_i ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_fetch_err_o$_DFFE_PN_  (.D(\if_stage_i.fetch_err ),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_fetch_err_i ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_fetch_err_plus2_o$_SDFFCE_PN0N_  (.D(_01579_),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_is_compressed_id_o$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.is_compressed_o ),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_is_compressed_i ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[0]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[0] ),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_i[0] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[10]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[10] ),
    .DE(net253),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[3] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[11]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[11] ),
    .DE(net253),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[12]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[12] ),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_i[12] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[13]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[13] ),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_i[13] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[14]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[14] ),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_i[14] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[15]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[15] ),
    .DE(net253),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[0] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[16]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[16] ),
    .DE(net253),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[1] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[17]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[17] ),
    .DE(net253),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[2] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[18]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[18] ),
    .DE(net253),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[3] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[19]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[19] ),
    .DE(net253),
    .Q(\gen_regfile_ff.register_file_i.raddr_a_i[4] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[1]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[1] ),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_i[1] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[20]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[20] ),
    .DE(net253),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[0] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[21]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[21] ),
    .DE(net253),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[1] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[22]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[22] ),
    .DE(net253),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[2] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[23]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[23] ),
    .DE(net253),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[3] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[24]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[24] ),
    .DE(net253),
    .Q(\gen_regfile_ff.register_file_i.raddr_b_i[4] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[25]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[25] ),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_i[25] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[26]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[26] ),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_i[26] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[27]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[27] ),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_i[27] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[28]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[28] ),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_i[28] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[29]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[29] ),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_i[29] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[2]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[2] ),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_i[2] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[30]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[30] ),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_i[30] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[31]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[31] ),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_i[31] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[3]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[3] ),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_i[3] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[4]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[4] ),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_i[4] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[5]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[5] ),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_i[5] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[6]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[6] ),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_i[6] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[7]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[7] ),
    .DE(net253),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[8]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[8] ),
    .DE(net253),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_alu_id_o[9]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_o[9] ),
    .DE(net253),
    .Q(\gen_regfile_ff.register_file_i.waddr_a_i[2] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[0]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_i[0] ),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_compressed_i[0] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[10]$_DFFE_PN_  (.D(_11074_),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_compressed_i[10] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[11]$_DFFE_PN_  (.D(_11078_),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_compressed_i[11] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[12]$_DFFE_PN_  (.D(_11115_),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_compressed_i[12] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[13]$_DFFE_PN_  (.D(_11055_),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_compressed_i[13] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[14]$_DFFE_PN_  (.D(_11061_),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_compressed_i[14] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[15]$_DFFE_PN_  (.D(_11068_),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_compressed_i[15] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[1]$_DFFE_PN_  (.D(_10839_),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_compressed_i[1] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[2]$_DFFE_PN_  (.D(_11091_),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_compressed_i[2] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[3]$_DFFE_PN_  (.D(_11095_),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_compressed_i[3] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[4]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_i[4] ),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_compressed_i[4] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[5]$_DFFE_PN_  (.D(_11082_),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_compressed_i[5] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[6]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_i[6] ),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_compressed_i[6] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[7]$_DFFE_PN_  (.D(_11103_),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_compressed_i[7] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[8]$_DFFE_PN_  (.D(_11107_),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_compressed_i[8] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.instr_rdata_c_id_o[9]$_DFFE_PN_  (.D(\if_stage_i.compressed_decoder_i.instr_i[9] ),
    .DE(net253),
    .Q(\id_stage_i.controller_i.instr_compressed_i[9] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_4 \if_stage_i.instr_valid_id_q$_DFF_PN0_  (.D(\if_stage_i.instr_valid_id_d ),
    .Q(\id_stage_i.controller_i.instr_valid_i ),
    .RESET_B(net455),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[10]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[10] ),
    .DE(_00007_),
    .Q(\cs_registers_i.pc_id_i[10] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[11]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[11] ),
    .DE(_00007_),
    .Q(\cs_registers_i.pc_id_i[11] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[12]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[12] ),
    .DE(_00007_),
    .Q(\cs_registers_i.pc_id_i[12] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[13]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[13] ),
    .DE(_00007_),
    .Q(\cs_registers_i.pc_id_i[13] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[14]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[14] ),
    .DE(_00007_),
    .Q(\cs_registers_i.pc_id_i[14] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[15]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[15] ),
    .DE(_00007_),
    .Q(\cs_registers_i.pc_id_i[15] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[16]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[16] ),
    .DE(net1328),
    .Q(\cs_registers_i.pc_id_i[16] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[17]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[17] ),
    .DE(net1328),
    .Q(\cs_registers_i.pc_id_i[17] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[18]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[18] ),
    .DE(net1328),
    .Q(\cs_registers_i.pc_id_i[18] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[19]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[19] ),
    .DE(net1328),
    .Q(\cs_registers_i.pc_id_i[19] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[1]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[1] ),
    .DE(net253),
    .Q(\cs_registers_i.pc_id_i[1] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[20]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[20] ),
    .DE(net1328),
    .Q(\cs_registers_i.pc_id_i[20] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[21]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[21] ),
    .DE(net1328),
    .Q(\cs_registers_i.pc_id_i[21] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[22]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[22] ),
    .DE(net1328),
    .Q(\cs_registers_i.pc_id_i[22] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[23]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[23] ),
    .DE(net1328),
    .Q(\cs_registers_i.pc_id_i[23] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[24]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[24] ),
    .DE(net1328),
    .Q(\cs_registers_i.pc_id_i[24] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[25]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[25] ),
    .DE(net1328),
    .Q(\cs_registers_i.pc_id_i[25] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[26]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[26] ),
    .DE(net1328),
    .Q(\cs_registers_i.pc_id_i[26] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[27]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[27] ),
    .DE(net1328),
    .Q(\cs_registers_i.pc_id_i[27] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[28]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[28] ),
    .DE(_00007_),
    .Q(\cs_registers_i.pc_id_i[28] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[29]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[29] ),
    .DE(_00007_),
    .Q(\cs_registers_i.pc_id_i[29] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[2]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[2] ),
    .DE(net1328),
    .Q(\cs_registers_i.pc_id_i[2] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[30]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[30] ),
    .DE(_00007_),
    .Q(\cs_registers_i.pc_id_i[30] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[31]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[31] ),
    .DE(_00007_),
    .Q(\cs_registers_i.pc_id_i[31] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[3]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[3] ),
    .DE(net1328),
    .Q(\cs_registers_i.pc_id_i[3] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[4]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[4] ),
    .DE(net1328),
    .Q(\cs_registers_i.pc_id_i[4] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[5]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[5] ),
    .DE(_00007_),
    .Q(\cs_registers_i.pc_id_i[5] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[6]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[6] ),
    .DE(_00007_),
    .Q(\cs_registers_i.pc_id_i[6] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[7]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[7] ),
    .DE(_00007_),
    .Q(\cs_registers_i.pc_id_i[7] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[8]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[8] ),
    .DE(_00007_),
    .Q(\cs_registers_i.pc_id_i[8] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \if_stage_i.pc_id_o[9]$_DFFE_PN_  (.D(\cs_registers_i.pc_if_i[9] ),
    .DE(_00007_),
    .Q(\cs_registers_i.pc_id_i[9] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[0]$_DFFE_PN0P_  (.D(_01580_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[0] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[10]$_DFFE_PN0P_  (.D(_01581_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[10] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[11]$_DFFE_PN0P_  (.D(_01582_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[11] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[12]$_DFFE_PN0P_  (.D(_01583_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[12] ),
    .RESET_B(net454),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[13]$_DFFE_PN0P_  (.D(_01584_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[13] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[14]$_DFFE_PN0P_  (.D(_01585_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[14] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[15]$_DFFE_PN0P_  (.D(_01586_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[15] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[16]$_DFFE_PN0P_  (.D(_01587_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[16] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[17]$_DFFE_PN0P_  (.D(_01588_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[17] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[18]$_DFFE_PN0P_  (.D(_01589_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[18] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[19]$_DFFE_PN0P_  (.D(_01590_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[19] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[1]$_DFFE_PN0P_  (.D(_01591_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[1] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[20]$_DFFE_PN0P_  (.D(_01592_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[20] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[21]$_DFFE_PN0P_  (.D(_01593_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[21] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[22]$_DFFE_PN0P_  (.D(_01594_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[22] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[23]$_DFFE_PN0P_  (.D(_01595_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[23] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[24]$_DFFE_PN0P_  (.D(_01596_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[24] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[25]$_DFFE_PN0P_  (.D(_01597_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[25] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[26]$_DFFE_PN0P_  (.D(_01598_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[26] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[27]$_DFFE_PN0P_  (.D(_01599_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[27] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[28]$_DFFE_PN0P_  (.D(_01600_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[28] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[29]$_DFFE_PN0P_  (.D(_01601_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[29] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfrtp_2 \load_store_unit_i.addr_last_q[2]$_DFFE_PN0P_  (.D(_01602_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[2] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[30]$_DFFE_PN0P_  (.D(_01603_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[30] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[31]$_DFFE_PN0P_  (.D(_01604_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[31] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfrtp_2 \load_store_unit_i.addr_last_q[3]$_DFFE_PN0P_  (.D(_01605_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[3] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[4]$_DFFE_PN0P_  (.D(_01606_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[4] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[5]$_DFFE_PN0P_  (.D(_01607_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[5] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[6]$_DFFE_PN0P_  (.D(_01608_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[6] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[7]$_DFFE_PN0P_  (.D(_01609_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[7] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_2 \load_store_unit_i.addr_last_q[8]$_DFFE_PN0P_  (.D(_01610_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[8] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.addr_last_q[9]$_DFFE_PN0P_  (.D(_01611_),
    .Q(\id_stage_i.controller_i.lsu_addr_last_i[9] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.data_sign_ext_q$_DFFE_PN0P_  (.D(_01612_),
    .Q(\load_store_unit_i.data_sign_ext_q ),
    .RESET_B(net456),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.data_we_q$_DFFE_PN0P_  (.D(_01613_),
    .Q(\load_store_unit_i.data_we_q ),
    .RESET_B(net455),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.handle_misaligned_q$_DFFE_PN0P_  (.D(_01614_),
    .Q(\load_store_unit_i.handle_misaligned_q ),
    .RESET_B(net457),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.ls_fsm_cs[0]$_DFFE_PN0P_  (.D(_01615_),
    .Q(\load_store_unit_i.ls_fsm_cs[0] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.ls_fsm_cs[1]$_DFFE_PN0P_  (.D(_01616_),
    .Q(\load_store_unit_i.ls_fsm_cs[1] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.ls_fsm_cs[2]$_DFFE_PN0P_  (.D(_01617_),
    .Q(\load_store_unit_i.ls_fsm_cs[2] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.lsu_err_q$_DFFE_PN0P_  (.D(_01618_),
    .Q(\load_store_unit_i.lsu_err_q ),
    .RESET_B(net455),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.rdata_offset_q[0]$_DFFE_PN0P_  (.D(_01619_),
    .Q(\load_store_unit_i.rdata_offset_q[0] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfrtp_4 \load_store_unit_i.rdata_offset_q[1]$_DFFE_PN0P_  (.D(_01620_),
    .Q(\load_store_unit_i.rdata_offset_q[1] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[0]$_DFFE_PN0P_  (.D(_01621_),
    .Q(\load_store_unit_i.rdata_q[8] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[10]$_DFFE_PN0P_  (.D(_01622_),
    .Q(\load_store_unit_i.rdata_q[18] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[11]$_DFFE_PN0P_  (.D(_01623_),
    .Q(\load_store_unit_i.rdata_q[19] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[12]$_DFFE_PN0P_  (.D(_01624_),
    .Q(\load_store_unit_i.rdata_q[20] ),
    .RESET_B(net455),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[13]$_DFFE_PN0P_  (.D(_01625_),
    .Q(\load_store_unit_i.rdata_q[21] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[14]$_DFFE_PN0P_  (.D(_01626_),
    .Q(\load_store_unit_i.rdata_q[22] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[15]$_DFFE_PN0P_  (.D(_01627_),
    .Q(\load_store_unit_i.rdata_q[23] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[16]$_DFFE_PN0P_  (.D(_01628_),
    .Q(\load_store_unit_i.rdata_q[24] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[17]$_DFFE_PN0P_  (.D(_01629_),
    .Q(\load_store_unit_i.rdata_q[25] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[18]$_DFFE_PN0P_  (.D(_01630_),
    .Q(\load_store_unit_i.rdata_q[26] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[19]$_DFFE_PN0P_  (.D(_01631_),
    .Q(\load_store_unit_i.rdata_q[27] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[1]$_DFFE_PN0P_  (.D(_01632_),
    .Q(\load_store_unit_i.rdata_q[9] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[20]$_DFFE_PN0P_  (.D(_01633_),
    .Q(\load_store_unit_i.rdata_q[28] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[21]$_DFFE_PN0P_  (.D(_01634_),
    .Q(\load_store_unit_i.rdata_q[29] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[22]$_DFFE_PN0P_  (.D(_01635_),
    .Q(\load_store_unit_i.rdata_q[30] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[23]$_DFFE_PN0P_  (.D(_01636_),
    .Q(\load_store_unit_i.rdata_q[31] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[2]$_DFFE_PN0P_  (.D(_01637_),
    .Q(\load_store_unit_i.rdata_q[10] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[3]$_DFFE_PN0P_  (.D(_01638_),
    .Q(\load_store_unit_i.rdata_q[11] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[4]$_DFFE_PN0P_  (.D(_01639_),
    .Q(\load_store_unit_i.rdata_q[12] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[5]$_DFFE_PN0P_  (.D(_01640_),
    .Q(\load_store_unit_i.rdata_q[13] ),
    .RESET_B(net457),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[6]$_DFFE_PN0P_  (.D(_01641_),
    .Q(\load_store_unit_i.rdata_q[14] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[7]$_DFFE_PN0P_  (.D(_01642_),
    .Q(\load_store_unit_i.rdata_q[15] ),
    .RESET_B(net456),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[8]$_DFFE_PN0P_  (.D(_01643_),
    .Q(\load_store_unit_i.rdata_q[16] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfrtp_1 \load_store_unit_i.rdata_q[9]$_DFFE_PN0P_  (.D(_01644_),
    .Q(\load_store_unit_i.rdata_q[17] ),
    .RESET_B(net460),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4079 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(boot_addr_i[10]),
    .X(net1));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(boot_addr_i[11]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(boot_addr_i[12]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(boot_addr_i[13]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(boot_addr_i[14]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(boot_addr_i[15]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(boot_addr_i[16]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(boot_addr_i[17]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(boot_addr_i[18]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(boot_addr_i[19]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(boot_addr_i[20]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(boot_addr_i[21]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(boot_addr_i[22]),
    .X(net13));
 sky130_fd_sc_hd__dlymetal6s2s_1 input14 (.A(boot_addr_i[23]),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(boot_addr_i[24]),
    .X(net15));
 sky130_fd_sc_hd__dlymetal6s2s_1 input16 (.A(boot_addr_i[25]),
    .X(net16));
 sky130_fd_sc_hd__dlymetal6s2s_1 input17 (.A(boot_addr_i[26]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(boot_addr_i[27]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(boot_addr_i[28]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(boot_addr_i[29]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(boot_addr_i[30]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(boot_addr_i[31]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(boot_addr_i[8]),
    .X(net23));
 sky130_fd_sc_hd__dlymetal6s2s_1 input24 (.A(boot_addr_i[9]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_4 input25 (.A(data_err_i),
    .X(net25));
 sky130_fd_sc_hd__buf_4 input26 (.A(data_gnt_i),
    .X(net26));
 sky130_fd_sc_hd__buf_4 input27 (.A(data_rdata_i[0]),
    .X(net27));
 sky130_fd_sc_hd__buf_4 input28 (.A(data_rdata_i[10]),
    .X(net28));
 sky130_fd_sc_hd__buf_4 input29 (.A(data_rdata_i[11]),
    .X(net29));
 sky130_fd_sc_hd__buf_4 input30 (.A(data_rdata_i[12]),
    .X(net30));
 sky130_fd_sc_hd__buf_4 input31 (.A(data_rdata_i[13]),
    .X(net31));
 sky130_fd_sc_hd__buf_4 input32 (.A(data_rdata_i[14]),
    .X(net32));
 sky130_fd_sc_hd__buf_4 input33 (.A(data_rdata_i[15]),
    .X(net33));
 sky130_fd_sc_hd__buf_4 input34 (.A(data_rdata_i[16]),
    .X(net34));
 sky130_fd_sc_hd__buf_4 input35 (.A(data_rdata_i[17]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 input36 (.A(data_rdata_i[18]),
    .X(net36));
 sky130_fd_sc_hd__buf_4 input37 (.A(data_rdata_i[19]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_4 input38 (.A(data_rdata_i[1]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_4 input39 (.A(data_rdata_i[20]),
    .X(net39));
 sky130_fd_sc_hd__buf_4 input40 (.A(data_rdata_i[21]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_4 input41 (.A(data_rdata_i[22]),
    .X(net41));
 sky130_fd_sc_hd__buf_4 input42 (.A(data_rdata_i[23]),
    .X(net42));
 sky130_fd_sc_hd__buf_4 input43 (.A(data_rdata_i[24]),
    .X(net43));
 sky130_fd_sc_hd__buf_4 input44 (.A(data_rdata_i[25]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 input45 (.A(data_rdata_i[26]),
    .X(net45));
 sky130_fd_sc_hd__buf_4 input46 (.A(data_rdata_i[27]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 input47 (.A(data_rdata_i[28]),
    .X(net47));
 sky130_fd_sc_hd__buf_4 input48 (.A(data_rdata_i[29]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 input49 (.A(data_rdata_i[2]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_4 input50 (.A(data_rdata_i[30]),
    .X(net50));
 sky130_fd_sc_hd__buf_4 input51 (.A(data_rdata_i[31]),
    .X(net51));
 sky130_fd_sc_hd__buf_4 input52 (.A(data_rdata_i[3]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_4 input53 (.A(data_rdata_i[4]),
    .X(net53));
 sky130_fd_sc_hd__buf_4 input54 (.A(data_rdata_i[5]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_4 input55 (.A(data_rdata_i[6]),
    .X(net55));
 sky130_fd_sc_hd__buf_4 input56 (.A(data_rdata_i[7]),
    .X(net56));
 sky130_fd_sc_hd__buf_4 input57 (.A(data_rdata_i[8]),
    .X(net57));
 sky130_fd_sc_hd__buf_4 input58 (.A(data_rdata_i[9]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_4 input59 (.A(data_rvalid_i),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_4 input60 (.A(debug_req_i),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(fetch_enable_i),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(hart_id_i[0]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(hart_id_i[10]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(hart_id_i[11]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(hart_id_i[12]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(hart_id_i[13]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(hart_id_i[14]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(hart_id_i[15]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(hart_id_i[16]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(hart_id_i[17]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(hart_id_i[18]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(hart_id_i[19]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_2 input73 (.A(hart_id_i[1]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 input74 (.A(hart_id_i[20]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 input75 (.A(hart_id_i[21]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(hart_id_i[22]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(hart_id_i[23]),
    .X(net77));
 sky130_fd_sc_hd__dlymetal6s2s_1 input78 (.A(hart_id_i[24]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input79 (.A(hart_id_i[25]),
    .X(net79));
 sky130_fd_sc_hd__dlymetal6s2s_1 input80 (.A(hart_id_i[26]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 input81 (.A(hart_id_i[27]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 input82 (.A(hart_id_i[28]),
    .X(net82));
 sky130_fd_sc_hd__dlymetal6s2s_1 input83 (.A(hart_id_i[29]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 input84 (.A(hart_id_i[2]),
    .X(net84));
 sky130_fd_sc_hd__dlymetal6s2s_1 input85 (.A(hart_id_i[30]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 input86 (.A(hart_id_i[31]),
    .X(net86));
 sky130_fd_sc_hd__dlymetal6s2s_1 input87 (.A(hart_id_i[3]),
    .X(net87));
 sky130_fd_sc_hd__dlymetal6s2s_1 input88 (.A(hart_id_i[4]),
    .X(net88));
 sky130_fd_sc_hd__dlymetal6s2s_1 input89 (.A(hart_id_i[5]),
    .X(net89));
 sky130_fd_sc_hd__dlymetal6s2s_1 input90 (.A(hart_id_i[6]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(hart_id_i[7]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 input92 (.A(hart_id_i[8]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 input93 (.A(hart_id_i[9]),
    .X(net93));
 sky130_fd_sc_hd__buf_2 input94 (.A(instr_err_i),
    .X(net94));
 sky130_fd_sc_hd__buf_4 input95 (.A(instr_gnt_i),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 input96 (.A(instr_rdata_i[0]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 input97 (.A(instr_rdata_i[10]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 input98 (.A(instr_rdata_i[11]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 input99 (.A(instr_rdata_i[12]),
    .X(net99));
 sky130_fd_sc_hd__dlymetal6s2s_1 input100 (.A(instr_rdata_i[13]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_2 input101 (.A(instr_rdata_i[14]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 input102 (.A(instr_rdata_i[15]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_2 input103 (.A(instr_rdata_i[16]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_2 input104 (.A(instr_rdata_i[17]),
    .X(net104));
 sky130_fd_sc_hd__dlymetal6s2s_1 input105 (.A(instr_rdata_i[18]),
    .X(net105));
 sky130_fd_sc_hd__dlymetal6s2s_1 input106 (.A(instr_rdata_i[19]),
    .X(net106));
 sky130_fd_sc_hd__buf_2 input107 (.A(instr_rdata_i[1]),
    .X(net107));
 sky130_fd_sc_hd__dlymetal6s2s_1 input108 (.A(instr_rdata_i[20]),
    .X(net108));
 sky130_fd_sc_hd__dlymetal6s2s_1 input109 (.A(instr_rdata_i[21]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 input110 (.A(instr_rdata_i[22]),
    .X(net110));
 sky130_fd_sc_hd__dlymetal6s2s_1 input111 (.A(instr_rdata_i[23]),
    .X(net111));
 sky130_fd_sc_hd__dlymetal6s2s_1 input112 (.A(instr_rdata_i[24]),
    .X(net112));
 sky130_fd_sc_hd__dlymetal6s2s_1 input113 (.A(instr_rdata_i[25]),
    .X(net113));
 sky130_fd_sc_hd__dlymetal6s2s_1 input114 (.A(instr_rdata_i[26]),
    .X(net114));
 sky130_fd_sc_hd__dlymetal6s2s_1 input115 (.A(instr_rdata_i[27]),
    .X(net115));
 sky130_fd_sc_hd__dlymetal6s2s_1 input116 (.A(instr_rdata_i[28]),
    .X(net116));
 sky130_fd_sc_hd__dlymetal6s2s_1 input117 (.A(instr_rdata_i[29]),
    .X(net117));
 sky130_fd_sc_hd__buf_2 input118 (.A(instr_rdata_i[2]),
    .X(net118));
 sky130_fd_sc_hd__dlymetal6s2s_1 input119 (.A(instr_rdata_i[30]),
    .X(net119));
 sky130_fd_sc_hd__dlymetal6s2s_1 input120 (.A(instr_rdata_i[31]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 input121 (.A(instr_rdata_i[3]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_2 input122 (.A(instr_rdata_i[4]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 input123 (.A(instr_rdata_i[5]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 input124 (.A(instr_rdata_i[6]),
    .X(net124));
 sky130_fd_sc_hd__buf_2 input125 (.A(instr_rdata_i[7]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_2 input126 (.A(instr_rdata_i[8]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 input127 (.A(instr_rdata_i[9]),
    .X(net127));
 sky130_fd_sc_hd__buf_2 input128 (.A(instr_rvalid_i),
    .X(net128));
 sky130_fd_sc_hd__dlymetal6s2s_1 input129 (.A(irq_external_i),
    .X(net129));
 sky130_fd_sc_hd__dlymetal6s2s_1 input130 (.A(irq_fast_i[0]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 input131 (.A(irq_fast_i[10]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_2 input132 (.A(irq_fast_i[11]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 input133 (.A(irq_fast_i[12]),
    .X(net133));
 sky130_fd_sc_hd__dlymetal6s2s_1 input134 (.A(irq_fast_i[13]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_2 input135 (.A(irq_fast_i[14]),
    .X(net135));
 sky130_fd_sc_hd__dlymetal6s2s_1 input136 (.A(irq_fast_i[1]),
    .X(net136));
 sky130_fd_sc_hd__dlymetal6s2s_1 input137 (.A(irq_fast_i[2]),
    .X(net137));
 sky130_fd_sc_hd__dlymetal6s2s_1 input138 (.A(irq_fast_i[3]),
    .X(net138));
 sky130_fd_sc_hd__buf_2 input139 (.A(irq_fast_i[4]),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_2 input140 (.A(irq_fast_i[5]),
    .X(net140));
 sky130_fd_sc_hd__dlymetal6s2s_1 input141 (.A(irq_fast_i[6]),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_2 input142 (.A(irq_fast_i[7]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_2 input143 (.A(irq_fast_i[8]),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_2 input144 (.A(irq_fast_i[9]),
    .X(net144));
 sky130_fd_sc_hd__buf_2 input145 (.A(irq_nm_i),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_2 input146 (.A(irq_software_i),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_2 input147 (.A(irq_timer_i),
    .X(net147));
 sky130_fd_sc_hd__buf_16 input148 (.A(rst_ni),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 input149 (.A(test_en_i),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_1 output150 (.A(net150),
    .X(core_sleep_o));
 sky130_fd_sc_hd__clkbuf_1 output151 (.A(net1578),
    .X(data_addr_o[10]));
 sky130_fd_sc_hd__clkbuf_1 output152 (.A(net152),
    .X(data_addr_o[11]));
 sky130_fd_sc_hd__clkbuf_1 output153 (.A(net1558),
    .X(data_addr_o[12]));
 sky130_fd_sc_hd__clkbuf_1 output154 (.A(net1571),
    .X(data_addr_o[13]));
 sky130_fd_sc_hd__clkbuf_1 output155 (.A(net1274),
    .X(data_addr_o[14]));
 sky130_fd_sc_hd__clkbuf_1 output156 (.A(net719),
    .X(data_addr_o[15]));
 sky130_fd_sc_hd__clkbuf_1 output157 (.A(net1582),
    .X(data_addr_o[16]));
 sky130_fd_sc_hd__clkbuf_1 output158 (.A(net1561),
    .X(data_addr_o[17]));
 sky130_fd_sc_hd__clkbuf_1 output159 (.A(net1241),
    .X(data_addr_o[18]));
 sky130_fd_sc_hd__clkbuf_1 output160 (.A(net1261),
    .X(data_addr_o[19]));
 sky130_fd_sc_hd__clkbuf_1 output161 (.A(net690),
    .X(data_addr_o[20]));
 sky130_fd_sc_hd__clkbuf_1 output162 (.A(net1258),
    .X(data_addr_o[21]));
 sky130_fd_sc_hd__clkbuf_1 output163 (.A(net1548),
    .X(data_addr_o[22]));
 sky130_fd_sc_hd__clkbuf_1 output164 (.A(net1244),
    .X(data_addr_o[23]));
 sky130_fd_sc_hd__clkbuf_1 output165 (.A(net774),
    .X(data_addr_o[24]));
 sky130_fd_sc_hd__clkbuf_1 output166 (.A(net166),
    .X(data_addr_o[25]));
 sky130_fd_sc_hd__clkbuf_1 output167 (.A(net167),
    .X(data_addr_o[26]));
 sky130_fd_sc_hd__clkbuf_1 output168 (.A(net687),
    .X(data_addr_o[27]));
 sky130_fd_sc_hd__clkbuf_1 output169 (.A(net492),
    .X(data_addr_o[28]));
 sky130_fd_sc_hd__clkbuf_1 output170 (.A(net170),
    .X(data_addr_o[29]));
 sky130_fd_sc_hd__clkbuf_1 output171 (.A(net171),
    .X(data_addr_o[2]));
 sky130_fd_sc_hd__clkbuf_1 output172 (.A(net172),
    .X(data_addr_o[30]));
 sky130_fd_sc_hd__clkbuf_1 output173 (.A(net481),
    .X(data_addr_o[31]));
 sky130_fd_sc_hd__clkbuf_1 output174 (.A(net1526),
    .X(data_addr_o[3]));
 sky130_fd_sc_hd__clkbuf_1 output175 (.A(net175),
    .X(data_addr_o[4]));
 sky130_fd_sc_hd__clkbuf_1 output176 (.A(net1040),
    .X(data_addr_o[5]));
 sky130_fd_sc_hd__clkbuf_1 output177 (.A(net177),
    .X(data_addr_o[6]));
 sky130_fd_sc_hd__clkbuf_1 output178 (.A(net178),
    .X(data_addr_o[7]));
 sky130_fd_sc_hd__clkbuf_1 output179 (.A(net179),
    .X(data_addr_o[8]));
 sky130_fd_sc_hd__clkbuf_1 output180 (.A(net1589),
    .X(data_addr_o[9]));
 sky130_fd_sc_hd__clkbuf_1 output181 (.A(net181),
    .X(data_be_o[0]));
 sky130_fd_sc_hd__clkbuf_1 output182 (.A(net182),
    .X(data_be_o[1]));
 sky130_fd_sc_hd__clkbuf_1 output183 (.A(net183),
    .X(data_be_o[2]));
 sky130_fd_sc_hd__clkbuf_1 output184 (.A(net184),
    .X(data_be_o[3]));
 sky130_fd_sc_hd__clkbuf_1 output185 (.A(net185),
    .X(data_req_o));
 sky130_fd_sc_hd__clkbuf_1 output186 (.A(net186),
    .X(data_wdata_o[0]));
 sky130_fd_sc_hd__clkbuf_1 output187 (.A(net187),
    .X(data_wdata_o[10]));
 sky130_fd_sc_hd__clkbuf_1 output188 (.A(net188),
    .X(data_wdata_o[11]));
 sky130_fd_sc_hd__clkbuf_1 output189 (.A(net189),
    .X(data_wdata_o[12]));
 sky130_fd_sc_hd__clkbuf_1 output190 (.A(net190),
    .X(data_wdata_o[13]));
 sky130_fd_sc_hd__clkbuf_1 output191 (.A(net191),
    .X(data_wdata_o[14]));
 sky130_fd_sc_hd__clkbuf_1 output192 (.A(net192),
    .X(data_wdata_o[15]));
 sky130_fd_sc_hd__clkbuf_1 output193 (.A(net193),
    .X(data_wdata_o[16]));
 sky130_fd_sc_hd__clkbuf_1 output194 (.A(net194),
    .X(data_wdata_o[17]));
 sky130_fd_sc_hd__clkbuf_1 output195 (.A(net195),
    .X(data_wdata_o[18]));
 sky130_fd_sc_hd__clkbuf_1 output196 (.A(net196),
    .X(data_wdata_o[19]));
 sky130_fd_sc_hd__clkbuf_1 output197 (.A(net197),
    .X(data_wdata_o[1]));
 sky130_fd_sc_hd__clkbuf_1 output198 (.A(net198),
    .X(data_wdata_o[20]));
 sky130_fd_sc_hd__clkbuf_1 output199 (.A(net199),
    .X(data_wdata_o[21]));
 sky130_fd_sc_hd__clkbuf_1 output200 (.A(net200),
    .X(data_wdata_o[22]));
 sky130_fd_sc_hd__clkbuf_1 output201 (.A(net201),
    .X(data_wdata_o[23]));
 sky130_fd_sc_hd__clkbuf_1 output202 (.A(net202),
    .X(data_wdata_o[24]));
 sky130_fd_sc_hd__clkbuf_1 output203 (.A(net203),
    .X(data_wdata_o[25]));
 sky130_fd_sc_hd__clkbuf_1 output204 (.A(net204),
    .X(data_wdata_o[26]));
 sky130_fd_sc_hd__clkbuf_1 output205 (.A(net205),
    .X(data_wdata_o[27]));
 sky130_fd_sc_hd__clkbuf_1 output206 (.A(net206),
    .X(data_wdata_o[28]));
 sky130_fd_sc_hd__clkbuf_1 output207 (.A(net207),
    .X(data_wdata_o[29]));
 sky130_fd_sc_hd__clkbuf_1 output208 (.A(net208),
    .X(data_wdata_o[2]));
 sky130_fd_sc_hd__clkbuf_1 output209 (.A(net209),
    .X(data_wdata_o[30]));
 sky130_fd_sc_hd__clkbuf_1 output210 (.A(net210),
    .X(data_wdata_o[31]));
 sky130_fd_sc_hd__clkbuf_1 output211 (.A(net211),
    .X(data_wdata_o[3]));
 sky130_fd_sc_hd__clkbuf_1 output212 (.A(net212),
    .X(data_wdata_o[4]));
 sky130_fd_sc_hd__clkbuf_1 output213 (.A(net213),
    .X(data_wdata_o[5]));
 sky130_fd_sc_hd__clkbuf_1 output214 (.A(net214),
    .X(data_wdata_o[6]));
 sky130_fd_sc_hd__clkbuf_1 output215 (.A(net215),
    .X(data_wdata_o[7]));
 sky130_fd_sc_hd__clkbuf_1 output216 (.A(net216),
    .X(data_wdata_o[8]));
 sky130_fd_sc_hd__clkbuf_1 output217 (.A(net217),
    .X(data_wdata_o[9]));
 sky130_fd_sc_hd__clkbuf_1 output218 (.A(net218),
    .X(data_we_o));
 sky130_fd_sc_hd__clkbuf_1 output219 (.A(net219),
    .X(instr_addr_o[10]));
 sky130_fd_sc_hd__clkbuf_1 output220 (.A(net220),
    .X(instr_addr_o[11]));
 sky130_fd_sc_hd__clkbuf_1 output221 (.A(net221),
    .X(instr_addr_o[12]));
 sky130_fd_sc_hd__clkbuf_1 output222 (.A(net222),
    .X(instr_addr_o[13]));
 sky130_fd_sc_hd__clkbuf_1 output223 (.A(net223),
    .X(instr_addr_o[14]));
 sky130_fd_sc_hd__clkbuf_1 output224 (.A(net224),
    .X(instr_addr_o[15]));
 sky130_fd_sc_hd__clkbuf_1 output225 (.A(net225),
    .X(instr_addr_o[16]));
 sky130_fd_sc_hd__clkbuf_1 output226 (.A(net226),
    .X(instr_addr_o[17]));
 sky130_fd_sc_hd__clkbuf_1 output227 (.A(net227),
    .X(instr_addr_o[18]));
 sky130_fd_sc_hd__clkbuf_1 output228 (.A(net228),
    .X(instr_addr_o[19]));
 sky130_fd_sc_hd__clkbuf_1 output229 (.A(net229),
    .X(instr_addr_o[20]));
 sky130_fd_sc_hd__clkbuf_1 output230 (.A(net230),
    .X(instr_addr_o[21]));
 sky130_fd_sc_hd__clkbuf_1 output231 (.A(net231),
    .X(instr_addr_o[22]));
 sky130_fd_sc_hd__clkbuf_1 output232 (.A(net232),
    .X(instr_addr_o[23]));
 sky130_fd_sc_hd__clkbuf_1 output233 (.A(net233),
    .X(instr_addr_o[24]));
 sky130_fd_sc_hd__clkbuf_1 output234 (.A(net234),
    .X(instr_addr_o[25]));
 sky130_fd_sc_hd__clkbuf_1 output235 (.A(net235),
    .X(instr_addr_o[26]));
 sky130_fd_sc_hd__clkbuf_1 output236 (.A(net236),
    .X(instr_addr_o[27]));
 sky130_fd_sc_hd__clkbuf_1 output237 (.A(net237),
    .X(instr_addr_o[28]));
 sky130_fd_sc_hd__clkbuf_1 output238 (.A(net238),
    .X(instr_addr_o[29]));
 sky130_fd_sc_hd__clkbuf_1 output239 (.A(net239),
    .X(instr_addr_o[2]));
 sky130_fd_sc_hd__clkbuf_1 output240 (.A(net240),
    .X(instr_addr_o[30]));
 sky130_fd_sc_hd__clkbuf_1 output241 (.A(net241),
    .X(instr_addr_o[31]));
 sky130_fd_sc_hd__clkbuf_1 output242 (.A(net242),
    .X(instr_addr_o[3]));
 sky130_fd_sc_hd__clkbuf_1 output243 (.A(net243),
    .X(instr_addr_o[4]));
 sky130_fd_sc_hd__clkbuf_1 output244 (.A(net244),
    .X(instr_addr_o[5]));
 sky130_fd_sc_hd__clkbuf_1 output245 (.A(net245),
    .X(instr_addr_o[6]));
 sky130_fd_sc_hd__clkbuf_1 output246 (.A(net246),
    .X(instr_addr_o[7]));
 sky130_fd_sc_hd__clkbuf_1 output247 (.A(net247),
    .X(instr_addr_o[8]));
 sky130_fd_sc_hd__clkbuf_1 output248 (.A(net248),
    .X(instr_addr_o[9]));
 sky130_fd_sc_hd__clkbuf_1 output249 (.A(net249),
    .X(instr_req_o));
 sky130_fd_sc_hd__buf_12 load_slew250 (.A(net1295),
    .X(net250));
 sky130_fd_sc_hd__buf_12 wire251 (.A(_04763_),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_16 load_slew252 (.A(_04661_),
    .X(net252));
 sky130_fd_sc_hd__buf_16 max_cap253 (.A(_00007_),
    .X(net253));
 sky130_fd_sc_hd__buf_12 wire254 (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .X(net254));
 sky130_fd_sc_hd__buf_16 max_cap255 (.A(_05502_),
    .X(net255));
 sky130_fd_sc_hd__buf_8 wire256 (.A(_05433_),
    .X(net256));
 sky130_fd_sc_hd__buf_16 max_cap257 (.A(_05268_),
    .X(net257));
 sky130_fd_sc_hd__buf_6 wire258 (.A(_01908_),
    .X(net258));
 sky130_fd_sc_hd__buf_16 load_slew259 (.A(net260),
    .X(net259));
 sky130_fd_sc_hd__buf_16 load_slew260 (.A(_05770_),
    .X(net260));
 sky130_fd_sc_hd__buf_6 load_slew261 (.A(_05706_),
    .X(net261));
 sky130_fd_sc_hd__buf_16 load_slew262 (.A(_05706_),
    .X(net262));
 sky130_fd_sc_hd__buf_16 load_slew263 (.A(_05640_),
    .X(net263));
 sky130_fd_sc_hd__buf_16 load_slew264 (.A(_05640_),
    .X(net264));
 sky130_fd_sc_hd__buf_8 load_slew265 (.A(net266),
    .X(net265));
 sky130_fd_sc_hd__buf_16 max_cap266 (.A(net267),
    .X(net266));
 sky130_fd_sc_hd__buf_8 load_slew267 (.A(_01665_),
    .X(net267));
 sky130_fd_sc_hd__buf_16 max_cap268 (.A(_11833_),
    .X(net268));
 sky130_fd_sc_hd__buf_16 load_slew269 (.A(_12760_),
    .X(net269));
 sky130_fd_sc_hd__buf_16 load_slew270 (.A(_12760_),
    .X(net270));
 sky130_fd_sc_hd__buf_16 load_slew271 (.A(_11243_),
    .X(net271));
 sky130_fd_sc_hd__buf_8 load_slew272 (.A(_12131_),
    .X(net272));
 sky130_fd_sc_hd__buf_8 wire273 (.A(_11328_),
    .X(net273));
 sky130_fd_sc_hd__buf_16 load_slew274 (.A(_11238_),
    .X(net274));
 sky130_fd_sc_hd__buf_16 load_slew275 (.A(net276),
    .X(net275));
 sky130_fd_sc_hd__buf_16 load_slew276 (.A(_13394_),
    .X(net276));
 sky130_fd_sc_hd__buf_16 load_slew277 (.A(net283),
    .X(net277));
 sky130_fd_sc_hd__buf_8 wire278 (.A(net279),
    .X(net278));
 sky130_fd_sc_hd__buf_8 load_slew279 (.A(net280),
    .X(net279));
 sky130_fd_sc_hd__buf_16 load_slew280 (.A(net282),
    .X(net280));
 sky130_fd_sc_hd__buf_16 load_slew281 (.A(net282),
    .X(net281));
 sky130_fd_sc_hd__buf_8 load_slew282 (.A(net283),
    .X(net282));
 sky130_fd_sc_hd__buf_8 load_slew283 (.A(_12685_),
    .X(net283));
 sky130_fd_sc_hd__buf_12 load_slew284 (.A(net285),
    .X(net284));
 sky130_fd_sc_hd__buf_16 wire285 (.A(_11267_),
    .X(net285));
 sky130_fd_sc_hd__buf_16 wire286 (.A(net287),
    .X(net286));
 sky130_fd_sc_hd__buf_16 load_slew287 (.A(_10970_),
    .X(net287));
 sky130_fd_sc_hd__buf_16 load_slew288 (.A(_10968_),
    .X(net288));
 sky130_fd_sc_hd__buf_12 wire289 (.A(_10968_),
    .X(net289));
 sky130_fd_sc_hd__buf_6 wire290 (.A(net291),
    .X(net290));
 sky130_fd_sc_hd__buf_6 wire291 (.A(net292),
    .X(net291));
 sky130_fd_sc_hd__buf_6 load_slew292 (.A(net293),
    .X(net292));
 sky130_fd_sc_hd__buf_6 load_slew293 (.A(_07330_),
    .X(net293));
 sky130_fd_sc_hd__buf_8 load_slew294 (.A(net295),
    .X(net294));
 sky130_fd_sc_hd__buf_8 load_slew295 (.A(_01762_),
    .X(net295));
 sky130_fd_sc_hd__buf_16 load_slew296 (.A(net694),
    .X(net296));
 sky130_fd_sc_hd__buf_16 load_slew297 (.A(net697),
    .X(net297));
 sky130_fd_sc_hd__buf_8 wire298 (.A(_12694_),
    .X(net298));
 sky130_fd_sc_hd__buf_16 load_slew299 (.A(net300),
    .X(net299));
 sky130_fd_sc_hd__buf_8 load_slew300 (.A(net637),
    .X(net300));
 sky130_fd_sc_hd__buf_8 load_slew301 (.A(net1206),
    .X(net301));
 sky130_fd_sc_hd__buf_8 load_slew302 (.A(net734),
    .X(net302));
 sky130_fd_sc_hd__buf_8 load_slew303 (.A(net304),
    .X(net303));
 sky130_fd_sc_hd__buf_6 load_slew304 (.A(net747),
    .X(net304));
 sky130_fd_sc_hd__buf_8 load_slew305 (.A(net306),
    .X(net305));
 sky130_fd_sc_hd__buf_6 wire306 (.A(_09928_),
    .X(net306));
 sky130_fd_sc_hd__buf_8 wire307 (.A(net931),
    .X(net307));
 sky130_fd_sc_hd__buf_12 load_slew308 (.A(net476),
    .X(net308));
 sky130_fd_sc_hd__buf_12 load_slew309 (.A(net480),
    .X(net309));
 sky130_fd_sc_hd__buf_12 load_slew310 (.A(_08370_),
    .X(net310));
 sky130_fd_sc_hd__buf_8 load_slew311 (.A(_03424_),
    .X(net311));
 sky130_fd_sc_hd__buf_8 load_slew312 (.A(net314),
    .X(net312));
 sky130_fd_sc_hd__buf_8 load_slew313 (.A(net314),
    .X(net313));
 sky130_fd_sc_hd__buf_8 load_slew314 (.A(net1103),
    .X(net314));
 sky130_fd_sc_hd__buf_6 wire315 (.A(net316),
    .X(net315));
 sky130_fd_sc_hd__bufbuf_16 wire316 (.A(_08284_),
    .X(net316));
 sky130_fd_sc_hd__buf_6 load_slew317 (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[2] ),
    .X(net317));
 sky130_fd_sc_hd__buf_6 wire318 (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[2] ),
    .X(net318));
 sky130_fd_sc_hd__buf_16 max_cap319 (.A(_08107_),
    .X(net319));
 sky130_fd_sc_hd__buf_12 load_slew320 (.A(_01712_),
    .X(net320));
 sky130_fd_sc_hd__buf_16 load_slew321 (.A(net322),
    .X(net321));
 sky130_fd_sc_hd__buf_16 wire322 (.A(_01702_),
    .X(net322));
 sky130_fd_sc_hd__buf_16 load_slew323 (.A(net1150),
    .X(net323));
 sky130_fd_sc_hd__buf_12 load_slew324 (.A(_08484_),
    .X(net324));
 sky130_fd_sc_hd__buf_12 load_slew325 (.A(_08464_),
    .X(net325));
 sky130_fd_sc_hd__buf_16 load_slew326 (.A(net1014),
    .X(net326));
 sky130_fd_sc_hd__buf_16 max_cap327 (.A(net1014),
    .X(net327));
 sky130_fd_sc_hd__buf_16 load_slew328 (.A(_08453_),
    .X(net328));
 sky130_fd_sc_hd__buf_12 load_slew329 (.A(net1202),
    .X(net329));
 sky130_fd_sc_hd__buf_12 load_slew330 (.A(_08331_),
    .X(net330));
 sky130_fd_sc_hd__buf_16 wire331 (.A(\gen_regfile_ff.register_file_i.waddr_a_i[0] ),
    .X(net331));
 sky130_fd_sc_hd__buf_8 load_slew332 (.A(net334),
    .X(net332));
 sky130_fd_sc_hd__buf_16 load_slew333 (.A(net334),
    .X(net333));
 sky130_fd_sc_hd__buf_16 wire334 (.A(\gen_regfile_ff.register_file_i.raddr_b_i[4] ),
    .X(net334));
 sky130_fd_sc_hd__buf_16 max_cap335 (.A(net336),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_16 wire336 (.A(net337),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_16 wire337 (.A(\gen_regfile_ff.register_file_i.raddr_b_i[3] ),
    .X(net337));
 sky130_fd_sc_hd__buf_16 load_slew338 (.A(net339),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_16 load_slew339 (.A(net343),
    .X(net339));
 sky130_fd_sc_hd__buf_16 load_slew340 (.A(net341),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_16 wire341 (.A(net343),
    .X(net341));
 sky130_fd_sc_hd__buf_16 load_slew342 (.A(net343),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_16 wire343 (.A(\gen_regfile_ff.register_file_i.raddr_b_i[2] ),
    .X(net343));
 sky130_fd_sc_hd__buf_16 load_slew344 (.A(net345),
    .X(net344));
 sky130_fd_sc_hd__buf_16 load_slew345 (.A(net346),
    .X(net345));
 sky130_fd_sc_hd__buf_8 load_slew346 (.A(net367),
    .X(net346));
 sky130_fd_sc_hd__buf_16 max_cap347 (.A(net348),
    .X(net347));
 sky130_fd_sc_hd__buf_16 load_slew348 (.A(net355),
    .X(net348));
 sky130_fd_sc_hd__buf_16 load_slew349 (.A(net352),
    .X(net349));
 sky130_fd_sc_hd__buf_16 load_slew350 (.A(net351),
    .X(net350));
 sky130_fd_sc_hd__buf_12 load_slew351 (.A(net352),
    .X(net351));
 sky130_fd_sc_hd__buf_16 load_slew352 (.A(net354),
    .X(net352));
 sky130_fd_sc_hd__buf_16 load_slew353 (.A(net354),
    .X(net353));
 sky130_fd_sc_hd__buf_16 load_slew354 (.A(net356),
    .X(net354));
 sky130_fd_sc_hd__buf_16 load_slew355 (.A(net356),
    .X(net355));
 sky130_fd_sc_hd__buf_16 load_slew356 (.A(net367),
    .X(net356));
 sky130_fd_sc_hd__buf_16 load_slew357 (.A(net358),
    .X(net357));
 sky130_fd_sc_hd__buf_16 load_slew358 (.A(net359),
    .X(net358));
 sky130_fd_sc_hd__buf_16 load_slew359 (.A(net364),
    .X(net359));
 sky130_fd_sc_hd__buf_16 load_slew360 (.A(net362),
    .X(net360));
 sky130_fd_sc_hd__buf_8 load_slew361 (.A(net362),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_16 wire362 (.A(net363),
    .X(net362));
 sky130_fd_sc_hd__buf_16 load_slew363 (.A(net365),
    .X(net363));
 sky130_fd_sc_hd__buf_16 max_cap364 (.A(net365),
    .X(net364));
 sky130_fd_sc_hd__buf_16 wire365 (.A(net366),
    .X(net365));
 sky130_fd_sc_hd__buf_16 load_slew366 (.A(net367),
    .X(net366));
 sky130_fd_sc_hd__buf_16 load_slew367 (.A(net511),
    .X(net367));
 sky130_fd_sc_hd__buf_16 load_slew368 (.A(net370),
    .X(net368));
 sky130_fd_sc_hd__buf_8 load_slew369 (.A(net370),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_16 wire370 (.A(net371),
    .X(net370));
 sky130_fd_sc_hd__buf_16 load_slew371 (.A(net512),
    .X(net371));
 sky130_fd_sc_hd__buf_16 load_slew372 (.A(net787),
    .X(net372));
 sky130_fd_sc_hd__buf_8 load_slew373 (.A(net375),
    .X(net373));
 sky130_fd_sc_hd__buf_16 load_slew374 (.A(net375),
    .X(net374));
 sky130_fd_sc_hd__buf_16 load_slew375 (.A(net381),
    .X(net375));
 sky130_fd_sc_hd__buf_16 load_slew376 (.A(net377),
    .X(net376));
 sky130_fd_sc_hd__buf_16 load_slew377 (.A(net378),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_16 load_slew378 (.A(net380),
    .X(net378));
 sky130_fd_sc_hd__buf_16 max_cap379 (.A(net654),
    .X(net379));
 sky130_fd_sc_hd__buf_16 max_cap380 (.A(net654),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_16 load_slew381 (.A(net653),
    .X(net381));
 sky130_fd_sc_hd__buf_6 load_slew382 (.A(net655),
    .X(net382));
 sky130_fd_sc_hd__buf_8 load_slew383 (.A(net386),
    .X(net383));
 sky130_fd_sc_hd__buf_16 load_slew384 (.A(net385),
    .X(net384));
 sky130_fd_sc_hd__buf_16 max_cap385 (.A(net386),
    .X(net385));
 sky130_fd_sc_hd__buf_16 wire386 (.A(\gen_regfile_ff.register_file_i.raddr_a_i[4] ),
    .X(net386));
 sky130_fd_sc_hd__buf_16 load_slew387 (.A(net388),
    .X(net387));
 sky130_fd_sc_hd__buf_16 max_cap388 (.A(net389),
    .X(net388));
 sky130_fd_sc_hd__buf_16 load_slew389 (.A(net390),
    .X(net389));
 sky130_fd_sc_hd__buf_16 load_slew390 (.A(net391),
    .X(net390));
 sky130_fd_sc_hd__buf_16 load_slew391 (.A(net392),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_16 wire392 (.A(\gen_regfile_ff.register_file_i.raddr_a_i[3] ),
    .X(net392));
 sky130_fd_sc_hd__buf_16 max_cap393 (.A(net394),
    .X(net393));
 sky130_fd_sc_hd__buf_16 load_slew394 (.A(net399),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_16 wire395 (.A(net396),
    .X(net395));
 sky130_fd_sc_hd__buf_12 load_slew396 (.A(net398),
    .X(net396));
 sky130_fd_sc_hd__buf_8 load_slew397 (.A(net398),
    .X(net397));
 sky130_fd_sc_hd__buf_16 load_slew398 (.A(net400),
    .X(net398));
 sky130_fd_sc_hd__buf_16 max_cap399 (.A(net400),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_16 load_slew400 (.A(\gen_regfile_ff.register_file_i.raddr_a_i[2] ),
    .X(net400));
 sky130_fd_sc_hd__buf_16 load_slew401 (.A(net402),
    .X(net401));
 sky130_fd_sc_hd__buf_16 load_slew402 (.A(net403),
    .X(net402));
 sky130_fd_sc_hd__buf_16 load_slew403 (.A(net415),
    .X(net403));
 sky130_fd_sc_hd__buf_16 load_slew404 (.A(net409),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_16 wire405 (.A(net410),
    .X(net405));
 sky130_fd_sc_hd__buf_8 load_slew406 (.A(net410),
    .X(net406));
 sky130_fd_sc_hd__buf_16 load_slew407 (.A(net408),
    .X(net407));
 sky130_fd_sc_hd__buf_16 load_slew408 (.A(net410),
    .X(net408));
 sky130_fd_sc_hd__buf_16 max_cap409 (.A(net410),
    .X(net409));
 sky130_fd_sc_hd__buf_16 max_cap410 (.A(net411),
    .X(net410));
 sky130_fd_sc_hd__buf_16 load_slew411 (.A(net414),
    .X(net411));
 sky130_fd_sc_hd__buf_6 load_slew412 (.A(net414),
    .X(net412));
 sky130_fd_sc_hd__buf_6 load_slew413 (.A(net414),
    .X(net413));
 sky130_fd_sc_hd__buf_16 max_cap414 (.A(net415),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_16 wire415 (.A(\gen_regfile_ff.register_file_i.raddr_a_i[1] ),
    .X(net415));
 sky130_fd_sc_hd__buf_16 max_cap416 (.A(net419),
    .X(net416));
 sky130_fd_sc_hd__buf_16 load_slew417 (.A(net418),
    .X(net417));
 sky130_fd_sc_hd__buf_16 load_slew418 (.A(net420),
    .X(net418));
 sky130_fd_sc_hd__buf_16 load_slew419 (.A(net420),
    .X(net419));
 sky130_fd_sc_hd__buf_16 load_slew420 (.A(net440),
    .X(net420));
 sky130_fd_sc_hd__buf_16 load_slew421 (.A(net422),
    .X(net421));
 sky130_fd_sc_hd__buf_16 max_cap422 (.A(net423),
    .X(net422));
 sky130_fd_sc_hd__clkbuf_16 wire423 (.A(net425),
    .X(net423));
 sky130_fd_sc_hd__buf_16 load_slew424 (.A(net425),
    .X(net424));
 sky130_fd_sc_hd__buf_16 max_cap425 (.A(net426),
    .X(net425));
 sky130_fd_sc_hd__buf_16 load_slew426 (.A(net427),
    .X(net426));
 sky130_fd_sc_hd__buf_16 load_slew427 (.A(net439),
    .X(net427));
 sky130_fd_sc_hd__buf_16 load_slew428 (.A(net430),
    .X(net428));
 sky130_fd_sc_hd__buf_16 load_slew429 (.A(net430),
    .X(net429));
 sky130_fd_sc_hd__buf_16 load_slew430 (.A(net431),
    .X(net430));
 sky130_fd_sc_hd__buf_16 load_slew431 (.A(net437),
    .X(net431));
 sky130_fd_sc_hd__buf_16 load_slew432 (.A(net433),
    .X(net432));
 sky130_fd_sc_hd__buf_12 load_slew433 (.A(net434),
    .X(net433));
 sky130_fd_sc_hd__buf_16 max_cap434 (.A(net435),
    .X(net434));
 sky130_fd_sc_hd__buf_16 load_slew435 (.A(net438),
    .X(net435));
 sky130_fd_sc_hd__buf_16 load_slew436 (.A(net438),
    .X(net436));
 sky130_fd_sc_hd__buf_16 load_slew437 (.A(net438),
    .X(net437));
 sky130_fd_sc_hd__buf_16 max_cap438 (.A(net439),
    .X(net438));
 sky130_fd_sc_hd__buf_16 max_cap439 (.A(net440),
    .X(net439));
 sky130_fd_sc_hd__clkbuf_16 wire440 (.A(\gen_regfile_ff.register_file_i.raddr_a_i[0] ),
    .X(net440));
 sky130_fd_sc_hd__buf_8 load_slew441 (.A(net443),
    .X(net441));
 sky130_fd_sc_hd__buf_16 load_slew442 (.A(net443),
    .X(net442));
 sky130_fd_sc_hd__buf_16 load_slew443 (.A(net444),
    .X(net443));
 sky130_fd_sc_hd__buf_16 load_slew444 (.A(net1087),
    .X(net444));
 sky130_fd_sc_hd__buf_8 load_slew445 (.A(net680),
    .X(net445));
 sky130_fd_sc_hd__buf_16 load_slew446 (.A(net447),
    .X(net446));
 sky130_fd_sc_hd__buf_16 load_slew447 (.A(net448),
    .X(net447));
 sky130_fd_sc_hd__buf_8 load_slew448 (.A(\gen_regfile_ff.register_file_i.waddr_a_i[4] ),
    .X(net448));
 sky130_fd_sc_hd__buf_16 load_slew449 (.A(net450),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_16 load_slew450 (.A(net451),
    .X(net450));
 sky130_fd_sc_hd__buf_16 load_slew451 (.A(\cs_registers_i.pc_if_i[1] ),
    .X(net451));
 sky130_fd_sc_hd__buf_16 wire452 (.A(net455),
    .X(net452));
 sky130_fd_sc_hd__buf_16 load_slew453 (.A(net454),
    .X(net453));
 sky130_fd_sc_hd__buf_16 load_slew454 (.A(net456),
    .X(net454));
 sky130_fd_sc_hd__buf_16 load_slew455 (.A(net456),
    .X(net455));
 sky130_fd_sc_hd__buf_16 load_slew456 (.A(net457),
    .X(net456));
 sky130_fd_sc_hd__buf_16 load_slew457 (.A(net458),
    .X(net457));
 sky130_fd_sc_hd__buf_16 load_slew458 (.A(net466),
    .X(net458));
 sky130_fd_sc_hd__buf_16 load_slew459 (.A(net460),
    .X(net459));
 sky130_fd_sc_hd__buf_16 wire460 (.A(net466),
    .X(net460));
 sky130_fd_sc_hd__buf_16 load_slew461 (.A(net463),
    .X(net461));
 sky130_fd_sc_hd__buf_16 load_slew462 (.A(net463),
    .X(net462));
 sky130_fd_sc_hd__buf_16 load_slew463 (.A(net464),
    .X(net463));
 sky130_fd_sc_hd__buf_16 load_slew464 (.A(net465),
    .X(net464));
 sky130_fd_sc_hd__buf_16 load_slew465 (.A(net466),
    .X(net465));
 sky130_fd_sc_hd__buf_16 load_slew466 (.A(net148),
    .X(net466));
 sky130_fd_sc_hd__buf_16 load_slew467 (.A(net468),
    .X(net467));
 sky130_fd_sc_hd__buf_16 load_slew468 (.A(net469),
    .X(net468));
 sky130_fd_sc_hd__buf_16 load_slew469 (.A(net148),
    .X(net469));
 sky130_fd_sc_hd__conb_1 ibex_core_470 (.LO(net470));
 sky130_fd_sc_hd__conb_1 _27319__471 (.LO(net471));
 sky130_fd_sc_hd__conb_1 _27320__472 (.LO(net472));
 sky130_fd_sc_hd__conb_1 _27321__473 (.LO(net473));
 sky130_fd_sc_hd__conb_1 _27352__474 (.LO(net474));
 sky130_fd_sc_hd__conb_1 _27353__475 (.LO(net475));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk_i (.A(clk_i),
    .X(clknet_0_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_1_0__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk_i_regs (.A(clknet_3_4__leaf_clk_i_regs),
    .X(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk_i_regs (.A(clknet_3_1__leaf_clk_i_regs),
    .X(clknet_leaf_1_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk_i_regs (.A(clknet_3_4__leaf_clk_i_regs),
    .X(clknet_leaf_2_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk_i_regs (.A(clknet_3_4__leaf_clk_i_regs),
    .X(clknet_leaf_3_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk_i_regs (.A(clknet_3_5__leaf_clk_i_regs),
    .X(clknet_leaf_4_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk_i_regs (.A(clknet_3_4__leaf_clk_i_regs),
    .X(clknet_leaf_5_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk_i_regs (.A(clknet_3_4__leaf_clk_i_regs),
    .X(clknet_leaf_6_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk_i_regs (.A(clknet_3_4__leaf_clk_i_regs),
    .X(clknet_leaf_7_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk_i_regs (.A(clknet_3_4__leaf_clk_i_regs),
    .X(clknet_leaf_8_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk_i_regs (.A(clknet_3_4__leaf_clk_i_regs),
    .X(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk_i_regs (.A(clknet_3_4__leaf_clk_i_regs),
    .X(clknet_leaf_10_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk_i_regs (.A(clknet_3_4__leaf_clk_i_regs),
    .X(clknet_leaf_11_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk_i_regs (.A(clknet_3_7__leaf_clk_i_regs),
    .X(clknet_leaf_12_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk_i_regs (.A(clknet_3_7__leaf_clk_i_regs),
    .X(clknet_leaf_13_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk_i_regs (.A(clknet_3_5__leaf_clk_i_regs),
    .X(clknet_leaf_14_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk_i_regs (.A(clknet_3_7__leaf_clk_i_regs),
    .X(clknet_leaf_15_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk_i_regs (.A(clknet_3_5__leaf_clk_i_regs),
    .X(clknet_leaf_16_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk_i_regs (.A(clknet_3_5__leaf_clk_i_regs),
    .X(clknet_leaf_17_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk_i_regs (.A(clknet_3_5__leaf_clk_i_regs),
    .X(clknet_leaf_18_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk_i_regs (.A(clknet_3_5__leaf_clk_i_regs),
    .X(clknet_leaf_19_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk_i_regs (.A(clknet_3_5__leaf_clk_i_regs),
    .X(clknet_leaf_20_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk_i_regs (.A(clknet_3_5__leaf_clk_i_regs),
    .X(clknet_leaf_21_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk_i_regs (.A(clknet_3_7__leaf_clk_i_regs),
    .X(clknet_leaf_22_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk_i_regs (.A(clknet_3_7__leaf_clk_i_regs),
    .X(clknet_leaf_23_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk_i_regs (.A(clknet_3_7__leaf_clk_i_regs),
    .X(clknet_leaf_24_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk_i_regs (.A(clknet_3_7__leaf_clk_i_regs),
    .X(clknet_leaf_25_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk_i_regs (.A(clknet_3_7__leaf_clk_i_regs),
    .X(clknet_leaf_26_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk_i_regs (.A(clknet_3_6__leaf_clk_i_regs),
    .X(clknet_leaf_27_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk_i_regs (.A(clknet_3_6__leaf_clk_i_regs),
    .X(clknet_leaf_28_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk_i_regs (.A(clknet_3_7__leaf_clk_i_regs),
    .X(clknet_leaf_29_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk_i_regs (.A(clknet_3_6__leaf_clk_i_regs),
    .X(clknet_leaf_30_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk_i_regs (.A(clknet_3_6__leaf_clk_i_regs),
    .X(clknet_leaf_31_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk_i_regs (.A(clknet_3_6__leaf_clk_i_regs),
    .X(clknet_leaf_32_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk_i_regs (.A(clknet_3_6__leaf_clk_i_regs),
    .X(clknet_leaf_33_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk_i_regs (.A(clknet_3_6__leaf_clk_i_regs),
    .X(clknet_leaf_34_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk_i_regs (.A(clknet_3_6__leaf_clk_i_regs),
    .X(clknet_leaf_35_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk_i_regs (.A(clknet_3_6__leaf_clk_i_regs),
    .X(clknet_leaf_36_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk_i_regs (.A(clknet_3_6__leaf_clk_i_regs),
    .X(clknet_leaf_37_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk_i_regs (.A(clknet_3_6__leaf_clk_i_regs),
    .X(clknet_leaf_38_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk_i_regs (.A(clknet_3_1__leaf_clk_i_regs),
    .X(clknet_leaf_39_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_40_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_41_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_42_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_43_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_44_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_45_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_46_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_48_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_49_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_50_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_51_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_52_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_54_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_55_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_57_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_58_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_59_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_60_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_61_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_63_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_64_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_69_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk_i_regs (.A(clknet_3_1__leaf_clk_i_regs),
    .X(clknet_leaf_70_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_71_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk_i_regs (.A(clknet_3_2__leaf_clk_i_regs),
    .X(clknet_leaf_72_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_73_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk_i_regs (.A(clknet_3_3__leaf_clk_i_regs),
    .X(clknet_leaf_74_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk_i_regs (.A(clknet_3_1__leaf_clk_i_regs),
    .X(clknet_leaf_75_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk_i_regs (.A(clknet_3_1__leaf_clk_i_regs),
    .X(clknet_leaf_76_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk_i_regs (.A(clknet_3_1__leaf_clk_i_regs),
    .X(clknet_leaf_77_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk_i_regs (.A(clknet_3_7__leaf_clk_i_regs),
    .X(clknet_leaf_78_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk_i_regs (.A(clknet_3_1__leaf_clk_i_regs),
    .X(clknet_leaf_79_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk_i_regs (.A(clknet_3_1__leaf_clk_i_regs),
    .X(clknet_leaf_80_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk_i_regs (.A(clknet_3_1__leaf_clk_i_regs),
    .X(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk_i_regs (.A(clknet_3_4__leaf_clk_i_regs),
    .X(clknet_leaf_82_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_83_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk_i_regs (.A(clknet_3_1__leaf_clk_i_regs),
    .X(clknet_leaf_85_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk_i_regs (.A(clknet_3_1__leaf_clk_i_regs),
    .X(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_88_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_90_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_91_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_92_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_93_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_94_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_95_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_96_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_97_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_98_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk_i_regs (.A(clknet_3_0__leaf_clk_i_regs),
    .X(clknet_leaf_99_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk_i_regs (.A(clk_i_regs),
    .X(clknet_0_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk_i_regs (.A(clknet_0_clk_i_regs),
    .X(clknet_3_0__leaf_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk_i_regs (.A(clknet_0_clk_i_regs),
    .X(clknet_3_1__leaf_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk_i_regs (.A(clknet_0_clk_i_regs),
    .X(clknet_3_2__leaf_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk_i_regs (.A(clknet_0_clk_i_regs),
    .X(clknet_3_3__leaf_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk_i_regs (.A(clknet_0_clk_i_regs),
    .X(clknet_3_4__leaf_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk_i_regs (.A(clknet_0_clk_i_regs),
    .X(clknet_3_5__leaf_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk_i_regs (.A(clknet_0_clk_i_regs),
    .X(clknet_3_6__leaf_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk_i_regs (.A(clknet_0_clk_i_regs),
    .X(clknet_3_7__leaf_clk_i_regs));
 sky130_fd_sc_hd__clkinv_16 clkload0 (.A(clknet_3_1__leaf_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkload1 (.A(clknet_3_2__leaf_clk_i_regs));
 sky130_fd_sc_hd__inv_16 clkload2 (.A(clknet_3_3__leaf_clk_i_regs));
 sky130_fd_sc_hd__clkinv_16 clkload3 (.A(clknet_3_4__leaf_clk_i_regs));
 sky130_fd_sc_hd__clkinv_16 clkload4 (.A(clknet_3_5__leaf_clk_i_regs));
 sky130_fd_sc_hd__clkinv_16 clkload5 (.A(clknet_3_6__leaf_clk_i_regs));
 sky130_fd_sc_hd__clkinv_16 clkload6 (.A(clknet_3_7__leaf_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload7 (.A(clknet_leaf_67_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload8 (.A(clknet_leaf_68_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload9 (.A(clknet_leaf_83_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload10 (.A(clknet_leaf_84_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload11 (.A(clknet_leaf_87_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload12 (.A(clknet_leaf_88_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload13 (.A(clknet_leaf_89_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload14 (.A(clknet_leaf_90_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload15 (.A(clknet_leaf_91_clk_i_regs));
 sky130_fd_sc_hd__clkinv_2 clkload16 (.A(clknet_leaf_92_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload17 (.A(clknet_leaf_93_clk_i_regs));
 sky130_fd_sc_hd__clkinv_2 clkload18 (.A(clknet_leaf_94_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload19 (.A(clknet_leaf_95_clk_i_regs));
 sky130_fd_sc_hd__bufinv_16 clkload20 (.A(clknet_leaf_96_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload21 (.A(clknet_leaf_98_clk_i_regs));
 sky130_fd_sc_hd__inv_6 clkload22 (.A(clknet_leaf_99_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload23 (.A(clknet_leaf_1_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload24 (.A(clknet_leaf_39_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload25 (.A(clknet_leaf_70_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload26 (.A(clknet_leaf_75_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload27 (.A(clknet_leaf_80_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload28 (.A(clknet_leaf_81_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload29 (.A(clknet_leaf_85_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload30 (.A(clknet_leaf_86_clk_i_regs));
 sky130_fd_sc_hd__clkinv_2 clkload31 (.A(clknet_leaf_52_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload32 (.A(clknet_leaf_53_clk_i_regs));
 sky130_fd_sc_hd__bufinv_16 clkload33 (.A(clknet_leaf_54_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload34 (.A(clknet_leaf_55_clk_i_regs));
 sky130_fd_sc_hd__clkinv_2 clkload35 (.A(clknet_leaf_56_clk_i_regs));
 sky130_fd_sc_hd__bufinv_16 clkload36 (.A(clknet_leaf_57_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload37 (.A(clknet_leaf_58_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload38 (.A(clknet_leaf_59_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload39 (.A(clknet_leaf_60_clk_i_regs));
 sky130_fd_sc_hd__bufinv_16 clkload40 (.A(clknet_leaf_61_clk_i_regs));
 sky130_fd_sc_hd__bufinv_16 clkload41 (.A(clknet_leaf_62_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload42 (.A(clknet_leaf_63_clk_i_regs));
 sky130_fd_sc_hd__clkinv_2 clkload43 (.A(clknet_leaf_64_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload44 (.A(clknet_leaf_65_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload45 (.A(clknet_leaf_66_clk_i_regs));
 sky130_fd_sc_hd__clkinv_2 clkload46 (.A(clknet_leaf_72_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload47 (.A(clknet_leaf_42_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload48 (.A(clknet_leaf_43_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload49 (.A(clknet_leaf_44_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload50 (.A(clknet_leaf_45_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload51 (.A(clknet_leaf_46_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload52 (.A(clknet_leaf_47_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload53 (.A(clknet_leaf_48_clk_i_regs));
 sky130_fd_sc_hd__bufinv_16 clkload54 (.A(clknet_leaf_49_clk_i_regs));
 sky130_fd_sc_hd__clkinv_2 clkload55 (.A(clknet_leaf_50_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload56 (.A(clknet_leaf_73_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload57 (.A(clknet_leaf_0_clk_i_regs));
 sky130_fd_sc_hd__clkinv_2 clkload58 (.A(clknet_leaf_3_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload59 (.A(clknet_leaf_5_clk_i_regs));
 sky130_fd_sc_hd__clkinv_2 clkload60 (.A(clknet_leaf_6_clk_i_regs));
 sky130_fd_sc_hd__clkinv_2 clkload61 (.A(clknet_leaf_7_clk_i_regs));
 sky130_fd_sc_hd__clkinv_2 clkload62 (.A(clknet_leaf_8_clk_i_regs));
 sky130_fd_sc_hd__clkinv_2 clkload63 (.A(clknet_leaf_9_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload64 (.A(clknet_leaf_10_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload65 (.A(clknet_leaf_11_clk_i_regs));
 sky130_fd_sc_hd__bufinv_16 clkload66 (.A(clknet_leaf_82_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload67 (.A(clknet_leaf_4_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload68 (.A(clknet_leaf_14_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload69 (.A(clknet_leaf_16_clk_i_regs));
 sky130_fd_sc_hd__bufinv_16 clkload70 (.A(clknet_leaf_17_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload71 (.A(clknet_leaf_19_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload72 (.A(clknet_leaf_20_clk_i_regs));
 sky130_fd_sc_hd__inv_6 clkload73 (.A(clknet_leaf_21_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload74 (.A(clknet_leaf_30_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload75 (.A(clknet_leaf_32_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload76 (.A(clknet_leaf_33_clk_i_regs));
 sky130_fd_sc_hd__clkinv_2 clkload77 (.A(clknet_leaf_36_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload78 (.A(clknet_leaf_37_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload79 (.A(clknet_leaf_38_clk_i_regs));
 sky130_fd_sc_hd__bufinv_16 clkload80 (.A(clknet_leaf_12_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_1 clkload81 (.A(clknet_leaf_13_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload82 (.A(clknet_leaf_15_clk_i_regs));
 sky130_fd_sc_hd__clkinv_2 clkload83 (.A(clknet_leaf_22_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload84 (.A(clknet_leaf_23_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload85 (.A(clknet_leaf_24_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_8 clkload86 (.A(clknet_leaf_25_clk_i_regs));
 sky130_fd_sc_hd__inv_6 clkload87 (.A(clknet_leaf_29_clk_i_regs));
 sky130_fd_sc_hd__clkinv_2 clkload88 (.A(clknet_leaf_78_clk_i_regs));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sky130_fd_sc_hd__inv_16 clkload89 (.A(clknet_3_0_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload90 (.A(clknet_3_1_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload91 (.A(clknet_3_2_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload92 (.A(clknet_3_3_0_clk));
 sky130_fd_sc_hd__clkinv_16 clkload93 (.A(clknet_3_4_0_clk));
 sky130_fd_sc_hd__inv_6 clkload94 (.A(clknet_3_5_0_clk));
 sky130_fd_sc_hd__inv_6 clkload95 (.A(clknet_3_7_0_clk));
 sky130_fd_sc_hd__clkinv_1 clkload96 (.A(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkinv_1 clkload97 (.A(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkinv_2 clkload98 (.A(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkinv_2 clkload99 (.A(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkinv_1 clkload100 (.A(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkinv_2 clkload101 (.A(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkinv_2 clkload102 (.A(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkinv_2 clkload103 (.A(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload104 (.A(clknet_leaf_6_clk));
 sky130_fd_sc_hd__bufinv_16 clkload105 (.A(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkinv_4 clkload106 (.A(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload107 (.A(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload108 (.A(clknet_leaf_77_clk));
 sky130_fd_sc_hd__bufinv_16 clkload109 (.A(clknet_leaf_78_clk));
 sky130_fd_sc_hd__inv_8 clkload110 (.A(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload111 (.A(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload112 (.A(clknet_leaf_10_clk));
 sky130_fd_sc_hd__inv_4 clkload113 (.A(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload114 (.A(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload115 (.A(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload116 (.A(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload117 (.A(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload118 (.A(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload119 (.A(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload120 (.A(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload121 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload122 (.A(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkinv_2 clkload123 (.A(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload124 (.A(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkinv_2 clkload125 (.A(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload126 (.A(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload127 (.A(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkinv_4 clkload128 (.A(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload129 (.A(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload130 (.A(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload131 (.A(clknet_leaf_66_clk));
 sky130_fd_sc_hd__bufinv_16 clkload132 (.A(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkinv_2 clkload133 (.A(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkinv_2 clkload134 (.A(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkinv_4 clkload135 (.A(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload136 (.A(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkinv_2 clkload137 (.A(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkinv_2 clkload138 (.A(clknet_leaf_55_clk));
 sky130_fd_sc_hd__bufinv_16 clkload139 (.A(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkinv_2 clkload140 (.A(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload141 (.A(clknet_leaf_64_clk));
 sky130_fd_sc_hd__bufinv_16 clkload142 (.A(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload143 (.A(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkinv_2 clkload144 (.A(clknet_leaf_68_clk));
 sky130_fd_sc_hd__bufinv_16 clkload145 (.A(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkinv_1 clkload146 (.A(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload147 (.A(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkinv_1 clkload148 (.A(clknet_leaf_34_clk));
 sky130_fd_sc_hd__bufinv_16 clkload149 (.A(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload150 (.A(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkinv_1 clkload151 (.A(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkinv_2 clkload152 (.A(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload153 (.A(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkinv_1 clkload154 (.A(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload155 (.A(clknet_leaf_42_clk));
 sky130_fd_sc_hd__bufinv_16 clkload156 (.A(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkinv_1 clkload157 (.A(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload158 (.A(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload159 (.A(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload160 (.A(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload161 (.A(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload162 (.A(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload163 (.A(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload164 (.A(clknet_leaf_51_clk));
 sky130_fd_sc_hd__bufinv_16 clkload165 (.A(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload166 (.A(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 delaybuf_0_core_clock (.A(delaynet_0_core_clock),
    .X(delaynet_1_core_clock));
 sky130_fd_sc_hd__clkbuf_16 delaybuf_1_core_clock (.A(delaynet_1_core_clock),
    .X(clk_i_regs));
 sky130_fd_sc_hd__buf_6 rebuffer1 (.A(_08743_),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net476),
    .X(net477));
 sky130_fd_sc_hd__clkbuf_16 clone879 (.A(net1014),
    .X(net1474));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(net476),
    .X(net479));
 sky130_fd_sc_hd__clkbuf_2 rebuffer5 (.A(net476),
    .X(net480));
 sky130_fd_sc_hd__buf_2 rebuffer6 (.A(net173),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer7 (.A(net481),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer8 (.A(net482),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net481),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer10 (.A(_08261_),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer11 (.A(net485),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer12 (.A(net486),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer13 (.A(_08261_),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer14 (.A(net488),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer15 (.A(net489),
    .X(net490));
 sky130_fd_sc_hd__buf_8 split16 (.A(net965),
    .X(net491));
 sky130_fd_sc_hd__buf_6 rebuffer17 (.A(net169),
    .X(net492));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer18 (.A(net492),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer19 (.A(net493),
    .X(net494));
 sky130_fd_sc_hd__buf_6 rebuffer20 (.A(_08895_),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer21 (.A(net495),
    .X(net496));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer22 (.A(net496),
    .X(net497));
 sky130_fd_sc_hd__buf_6 rebuffer23 (.A(_09147_),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer24 (.A(net498),
    .X(net499));
 sky130_fd_sc_hd__o211ai_4 clone25 (.A1(_05193_),
    .A2(_05252_),
    .B1(_05260_),
    .C1(_11824_),
    .Y(net500));
 sky130_fd_sc_hd__clkbuf_4 rebuffer26 (.A(_08476_),
    .X(net501));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer27 (.A(net501),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer28 (.A(net501),
    .X(net503));
 sky130_fd_sc_hd__buf_2 rebuffer29 (.A(net501),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer30 (.A(net504),
    .X(net505));
 sky130_fd_sc_hd__buf_12 rebuffer31 (.A(_08476_),
    .X(net506));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer32 (.A(net506),
    .X(net507));
 sky130_fd_sc_hd__buf_12 rebuffer33 (.A(net507),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer34 (.A(net508),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer35 (.A(net508),
    .X(net510));
 sky130_fd_sc_hd__buf_6 rebuffer36 (.A(\gen_regfile_ff.register_file_i.raddr_b_i[1] ),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer37 (.A(net511),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer38 (.A(net511),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer39 (.A(net513),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer40 (.A(net514),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer41 (.A(net514),
    .X(net516));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer42 (.A(_08471_),
    .X(net517));
 sky130_fd_sc_hd__buf_6 rebuffer43 (.A(net517),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer44 (.A(net518),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer45 (.A(net518),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer46 (.A(net1280),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer47 (.A(net521),
    .X(net522));
 sky130_fd_sc_hd__clkbuf_4 rebuffer48 (.A(_08471_),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer49 (.A(net523),
    .X(net524));
 sky130_fd_sc_hd__buf_8 rebuffer50 (.A(net523),
    .X(net525));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer51 (.A(net525),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer52 (.A(_08258_),
    .X(net527));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer53 (.A(_08258_),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer54 (.A(_08258_),
    .X(net529));
 sky130_fd_sc_hd__buf_2 rebuffer55 (.A(_08331_),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer56 (.A(_08331_),
    .X(net531));
 sky130_fd_sc_hd__buf_2 rebuffer57 (.A(_08331_),
    .X(net532));
 sky130_fd_sc_hd__buf_4 rebuffer58 (.A(net532),
    .X(net533));
 sky130_fd_sc_hd__buf_6 rebuffer59 (.A(net533),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer60 (.A(_08590_),
    .X(net535));
 sky130_fd_sc_hd__buf_6 rebuffer61 (.A(net715),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer62 (.A(net956),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer63 (.A(_08321_),
    .X(net538));
 sky130_fd_sc_hd__buf_2 rebuffer64 (.A(_08321_),
    .X(net539));
 sky130_fd_sc_hd__buf_2 rebuffer65 (.A(net539),
    .X(net540));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer66 (.A(net539),
    .X(net541));
 sky130_fd_sc_hd__buf_2 rebuffer67 (.A(_08321_),
    .X(net542));
 sky130_fd_sc_hd__buf_2 rebuffer68 (.A(net542),
    .X(net543));
 sky130_fd_sc_hd__buf_6 rebuffer69 (.A(net542),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer70 (.A(\gen_regfile_ff.register_file_i.raddr_b_i[3] ),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer71 (.A(net545),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer72 (.A(net546),
    .X(net547));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer73 (.A(net545),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer74 (.A(_08610_),
    .X(net549));
 sky130_fd_sc_hd__buf_6 rebuffer75 (.A(net712),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer76 (.A(\gen_regfile_ff.register_file_i.raddr_b_i[2] ),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer77 (.A(net551),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer78 (.A(net552),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer79 (.A(net552),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer80 (.A(net554),
    .X(net555));
 sky130_fd_sc_hd__buf_6 rebuffer81 (.A(_08597_),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer82 (.A(net556),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer83 (.A(net557),
    .X(net558));
 sky130_fd_sc_hd__buf_12 rebuffer84 (.A(_09035_),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer85 (.A(net559),
    .X(net560));
 sky130_fd_sc_hd__buf_4 rebuffer86 (.A(net560),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer87 (.A(_09035_),
    .X(net562));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer88 (.A(net562),
    .X(net563));
 sky130_fd_sc_hd__buf_6 split89 (.A(net994),
    .X(net564));
 sky130_fd_sc_hd__and2_4 clone90 (.A(net1225),
    .B(net394),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer91 (.A(net1118),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer92 (.A(net566),
    .X(net567));
 sky130_fd_sc_hd__buf_6 rebuffer93 (.A(net1118),
    .X(net568));
 sky130_fd_sc_hd__buf_2 rebuffer94 (.A(net568),
    .X(net569));
 sky130_fd_sc_hd__clkbuf_2 rebuffer95 (.A(net1118),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer96 (.A(\gen_regfile_ff.register_file_i.raddr_a_i[0] ),
    .X(net571));
 sky130_fd_sc_hd__clkbuf_2 rebuffer97 (.A(net1285),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer98 (.A(net572),
    .X(net573));
 sky130_fd_sc_hd__buf_4 rebuffer99 (.A(net573),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer100 (.A(net1032),
    .X(net575));
 sky130_fd_sc_hd__clkbuf_2 rebuffer101 (.A(net1032),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer102 (.A(net576),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer103 (.A(net577),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer104 (.A(net577),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer105 (.A(net579),
    .X(net580));
 sky130_fd_sc_hd__buf_2 rebuffer106 (.A(net580),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer107 (.A(net581),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer108 (.A(net581),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer109 (.A(net576),
    .X(net584));
 sky130_fd_sc_hd__buf_1 rebuffer110 (.A(net864),
    .X(net585));
 sky130_fd_sc_hd__clkbuf_2 rebuffer111 (.A(_08599_),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer112 (.A(\gen_regfile_ff.register_file_i.raddr_a_i[3] ),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer113 (.A(net587),
    .X(net588));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer114 (.A(_08457_),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer115 (.A(net589),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer116 (.A(net589),
    .X(net591));
 sky130_fd_sc_hd__buf_2 rebuffer117 (.A(net1014),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer118 (.A(net592),
    .X(net593));
 sky130_fd_sc_hd__buf_6 rebuffer119 (.A(_08202_),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer120 (.A(net594),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer121 (.A(net594),
    .X(net596));
 sky130_fd_sc_hd__buf_6 rebuffer122 (.A(net594),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer123 (.A(net597),
    .X(net598));
 sky130_fd_sc_hd__buf_4 rebuffer124 (.A(net597),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer125 (.A(net597),
    .X(net600));
 sky130_fd_sc_hd__buf_4 rebuffer126 (.A(_08901_),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer127 (.A(net601),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer128 (.A(net601),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer129 (.A(net601),
    .X(net604));
 sky130_fd_sc_hd__clkbuf_2 rebuffer130 (.A(_08901_),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer131 (.A(net605),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer132 (.A(net605),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer133 (.A(net1247),
    .X(net608));
 sky130_fd_sc_hd__buf_2 rebuffer134 (.A(_08344_),
    .X(net609));
 sky130_fd_sc_hd__buf_2 rebuffer135 (.A(net609),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer136 (.A(net610),
    .X(net611));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer137 (.A(net609),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer138 (.A(_08807_),
    .X(net613));
 sky130_fd_sc_hd__buf_12 rebuffer139 (.A(_08807_),
    .X(net614));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer140 (.A(net614),
    .X(net615));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer141 (.A(net615),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer142 (.A(net614),
    .X(net617));
 sky130_fd_sc_hd__buf_2 rebuffer143 (.A(_08606_),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer144 (.A(net618),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer145 (.A(net619),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer146 (.A(net1002),
    .X(net621));
 sky130_fd_sc_hd__buf_4 rebuffer147 (.A(_08799_),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer148 (.A(net622),
    .X(net623));
 sky130_fd_sc_hd__buf_8 rebuffer149 (.A(net622),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer150 (.A(net624),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer151 (.A(net624),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer152 (.A(\gen_regfile_ff.register_file_i.raddr_a_i[1] ),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer153 (.A(_08910_),
    .X(net628));
 sky130_fd_sc_hd__buf_2 rebuffer154 (.A(_08910_),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer155 (.A(net629),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer156 (.A(net629),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer157 (.A(net629),
    .X(net632));
 sky130_fd_sc_hd__clkbuf_2 rebuffer158 (.A(_08910_),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer159 (.A(net633),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer160 (.A(net633),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer161 (.A(_08949_),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer162 (.A(net636),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer163 (.A(net637),
    .X(net638));
 sky130_fd_sc_hd__buf_1 rebuffer164 (.A(net636),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer165 (.A(net639),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer166 (.A(net640),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer167 (.A(net641),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer168 (.A(net636),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer169 (.A(_08414_),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer170 (.A(_08414_),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer171 (.A(_08414_),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer172 (.A(net646),
    .X(net647));
 sky130_fd_sc_hd__buf_2 rebuffer173 (.A(net834),
    .X(net648));
 sky130_fd_sc_hd__nor2_8 clone174 (.A(net405),
    .B(net393),
    .Y(net649));
 sky130_fd_sc_hd__nor2_4 clone175 (.A(net338),
    .B(net377),
    .Y(net650));
 sky130_fd_sc_hd__buf_12 rebuffer983 (.A(net151),
    .X(net1578));
 sky130_fd_sc_hd__o211ai_4 clone177 (.A1(_05193_),
    .A2(_05252_),
    .B1(_05260_),
    .C1(_11824_),
    .Y(net652));
 sky130_fd_sc_hd__buf_4 rebuffer178 (.A(net809),
    .X(net653));
 sky130_fd_sc_hd__buf_6 rebuffer179 (.A(\gen_regfile_ff.register_file_i.raddr_b_i[0] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer180 (.A(net1059),
    .X(net655));
 sky130_fd_sc_hd__buf_12 rebuffer181 (.A(_10216_),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer182 (.A(net656),
    .X(net657));
 sky130_fd_sc_hd__clkbuf_2 rebuffer183 (.A(net982),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer184 (.A(net658),
    .X(net659));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer185 (.A(net658),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer186 (.A(\gen_regfile_ff.register_file_i.raddr_a_i[2] ),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer187 (.A(net661),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer188 (.A(\id_stage_i.controller_i.instr_i[26] ),
    .X(net663));
 sky130_fd_sc_hd__buf_6 rebuffer189 (.A(\id_stage_i.controller_i.instr_i[26] ),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer190 (.A(net664),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer191 (.A(net664),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer192 (.A(net664),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer193 (.A(net667),
    .X(net668));
 sky130_fd_sc_hd__buf_6 rebuffer194 (.A(\id_stage_i.controller_i.instr_i[29] ),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer195 (.A(net669),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer196 (.A(net670),
    .X(net671));
 sky130_fd_sc_hd__buf_6 rebuffer197 (.A(net669),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer198 (.A(net672),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer199 (.A(net672),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer200 (.A(net674),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer201 (.A(\id_stage_i.controller_i.instr_i[13] ),
    .X(net676));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer202 (.A(\id_stage_i.controller_i.instr_i[13] ),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer203 (.A(net677),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer204 (.A(\id_stage_i.controller_i.instr_i[13] ),
    .X(net679));
 sky130_fd_sc_hd__buf_6 rebuffer205 (.A(\id_stage_i.controller_i.instr_i[13] ),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer206 (.A(net680),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer207 (.A(\id_stage_i.controller_i.instr_i[13] ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer208 (.A(net682),
    .X(net683));
 sky130_fd_sc_hd__buf_12 rebuffer209 (.A(_10407_),
    .X(net684));
 sky130_fd_sc_hd__a31oi_4 clone210 (.A1(net686),
    .A2(net266),
    .A3(_05186_),
    .B1(_05190_),
    .Y(net685));
 sky130_fd_sc_hd__buf_12 rebuffer211 (.A(net860),
    .X(net686));
 sky130_fd_sc_hd__buf_12 rebuffer212 (.A(net168),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer213 (.A(net687),
    .X(net688));
 sky130_fd_sc_hd__clkbuf_4 rebuffer214 (.A(net161),
    .X(net689));
 sky130_fd_sc_hd__buf_2 rebuffer215 (.A(net689),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer216 (.A(net690),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer217 (.A(net689),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer218 (.A(net692),
    .X(net693));
 sky130_fd_sc_hd__buf_8 rebuffer219 (.A(_08431_),
    .X(net694));
 sky130_fd_sc_hd__buf_2 rebuffer220 (.A(net694),
    .X(net695));
 sky130_fd_sc_hd__buf_4 rebuffer221 (.A(net695),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer222 (.A(net694),
    .X(net697));
 sky130_fd_sc_hd__nor2_4 clone223 (.A(net337),
    .B(_08161_),
    .Y(net698));
 sky130_fd_sc_hd__and4_2 clone224 (.A(net861),
    .B(net980),
    .C(net986),
    .D(net985),
    .X(net699));
 sky130_fd_sc_hd__buf_12 rebuffer225 (.A(_08734_),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer226 (.A(net700),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer227 (.A(net700),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer228 (.A(net702),
    .X(net703));
 sky130_fd_sc_hd__buf_4 rebuffer229 (.A(net702),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer230 (.A(net704),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer231 (.A(_08734_),
    .X(net706));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer232 (.A(net706),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer233 (.A(_08796_),
    .X(net708));
 sky130_fd_sc_hd__buf_6 rebuffer234 (.A(net708),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer235 (.A(net709),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer236 (.A(net709),
    .X(net711));
 sky130_fd_sc_hd__clkbuf_2 rebuffer237 (.A(_08610_),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer238 (.A(net712),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer239 (.A(net713),
    .X(net714));
 sky130_fd_sc_hd__buf_2 rebuffer240 (.A(_08590_),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer241 (.A(net715),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer242 (.A(net716),
    .X(net717));
 sky130_fd_sc_hd__buf_12 rebuffer982 (.A(_03736_),
    .X(net1577));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer244 (.A(net721),
    .X(net719));
 sky130_fd_sc_hd__a21oi_2 clone981 (.A1(net1577),
    .A2(net266),
    .B1(_03738_),
    .Y(net1576));
 sky130_fd_sc_hd__buf_12 rebuffer246 (.A(net156),
    .X(net721));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer247 (.A(_08999_),
    .X(net722));
 sky130_fd_sc_hd__bufbuf_16 rebuffer248 (.A(_08999_),
    .X(net723));
 sky130_fd_sc_hd__buf_4 rebuffer249 (.A(net723),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer250 (.A(net724),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer251 (.A(net725),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer252 (.A(net726),
    .X(net727));
 sky130_fd_sc_hd__buf_2 rebuffer253 (.A(_08999_),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer254 (.A(net728),
    .X(net729));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer255 (.A(net729),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer256 (.A(_08897_),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer257 (.A(net731),
    .X(net732));
 sky130_fd_sc_hd__buf_2 rebuffer258 (.A(net423),
    .X(net733));
 sky130_fd_sc_hd__buf_6 rebuffer259 (.A(_02009_),
    .X(net734));
 sky130_fd_sc_hd__buf_2 rebuffer260 (.A(net734),
    .X(net735));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer261 (.A(net735),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer262 (.A(_09450_),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer263 (.A(_09450_),
    .X(net738));
 sky130_fd_sc_hd__or3_4 clone264 (.A(_08293_),
    .B(_08294_),
    .C(_08265_),
    .X(net739));
 sky130_fd_sc_hd__buf_12 rebuffer265 (.A(_05261_),
    .X(net740));
 sky130_fd_sc_hd__buf_8 rebuffer266 (.A(_01966_),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer267 (.A(net741),
    .X(net742));
 sky130_fd_sc_hd__buf_6 rebuffer268 (.A(_10254_),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer269 (.A(net743),
    .X(net744));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer270 (.A(net743),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer271 (.A(_09995_),
    .X(net746));
 sky130_fd_sc_hd__buf_6 rebuffer272 (.A(_09995_),
    .X(net747));
 sky130_fd_sc_hd__clkbuf_2 rebuffer273 (.A(net747),
    .X(net748));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer274 (.A(net748),
    .X(net749));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer275 (.A(net748),
    .X(net750));
 sky130_fd_sc_hd__buf_2 rebuffer276 (.A(_08839_),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer277 (.A(net853),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer278 (.A(net853),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer279 (.A(\gen_regfile_ff.register_file_i.raddr_b_i[4] ),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer280 (.A(net754),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer281 (.A(net755),
    .X(net756));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer282 (.A(_08606_),
    .X(net757));
 sky130_fd_sc_hd__clkbuf_2 rebuffer283 (.A(_08606_),
    .X(net758));
 sky130_fd_sc_hd__buf_6 rebuffer284 (.A(_09060_),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer285 (.A(net759),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer286 (.A(net759),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer287 (.A(net759),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer288 (.A(net759),
    .X(net763));
 sky130_fd_sc_hd__buf_2 rebuffer289 (.A(_09060_),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer290 (.A(net764),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer291 (.A(net764),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer292 (.A(_08359_),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer293 (.A(net767),
    .X(net768));
 sky130_fd_sc_hd__buf_2 rebuffer294 (.A(_09651_),
    .X(net769));
 sky130_fd_sc_hd__buf_6 rebuffer295 (.A(_09054_),
    .X(net770));
 sky130_fd_sc_hd__buf_2 rebuffer296 (.A(net770),
    .X(net771));
 sky130_fd_sc_hd__buf_12 rebuffer297 (.A(_09054_),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer298 (.A(net772),
    .X(net773));
 sky130_fd_sc_hd__buf_12 rebuffer299 (.A(net165),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer300 (.A(net774),
    .X(net775));
 sky130_fd_sc_hd__buf_12 rebuffer301 (.A(_09751_),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer302 (.A(net776),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer303 (.A(_09044_),
    .X(net778));
 sky130_fd_sc_hd__buf_6 rebuffer304 (.A(_10806_),
    .X(net779));
 sky130_fd_sc_hd__buf_4 rebuffer305 (.A(net1209),
    .X(net780));
 sky130_fd_sc_hd__and2_2 clone306 (.A(net929),
    .B(net1208),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer307 (.A(_09086_),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer308 (.A(net782),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer309 (.A(net783),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer310 (.A(_08693_),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer311 (.A(net415),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer312 (.A(\gen_regfile_ff.register_file_i.raddr_b_i[1] ),
    .X(net787));
 sky130_fd_sc_hd__buf_8 rebuffer313 (.A(_01978_),
    .X(net788));
 sky130_fd_sc_hd__buf_6 rebuffer314 (.A(net788),
    .X(net789));
 sky130_fd_sc_hd__buf_8 rebuffer315 (.A(net789),
    .X(net790));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer316 (.A(net790),
    .X(net791));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer317 (.A(net791),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer318 (.A(_13466_),
    .X(net793));
 sky130_fd_sc_hd__buf_6 clone319 (.A(net795),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer320 (.A(\gen_regfile_ff.register_file_i.raddr_a_i[1] ),
    .X(net795));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer321 (.A(_09104_),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer322 (.A(net796),
    .X(net797));
 sky130_fd_sc_hd__buf_4 rebuffer323 (.A(net797),
    .X(net798));
 sky130_fd_sc_hd__clkbuf_16 clone324 (.A(net856),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer325 (.A(_09148_),
    .X(net800));
 sky130_fd_sc_hd__buf_6 rebuffer326 (.A(\id_stage_i.controller_i.instr_i[27] ),
    .X(net801));
 sky130_fd_sc_hd__buf_6 rebuffer327 (.A(net801),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer328 (.A(net802),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer329 (.A(net802),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer330 (.A(net804),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer331 (.A(net801),
    .X(net806));
 sky130_fd_sc_hd__buf_4 rebuffer332 (.A(_09054_),
    .X(net807));
 sky130_fd_sc_hd__buf_6 rebuffer333 (.A(_09054_),
    .X(net808));
 sky130_fd_sc_hd__clkbuf_2 rebuffer334 (.A(\gen_regfile_ff.register_file_i.raddr_b_i[0] ),
    .X(net809));
 sky130_fd_sc_hd__buf_2 rebuffer335 (.A(\gen_regfile_ff.register_file_i.raddr_b_i[0] ),
    .X(net810));
 sky130_fd_sc_hd__buf_6 rebuffer336 (.A(\id_stage_i.controller_i.instr_i[28] ),
    .X(net811));
 sky130_fd_sc_hd__buf_6 rebuffer337 (.A(net811),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer338 (.A(net812),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer339 (.A(net812),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer340 (.A(net814),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer341 (.A(net811),
    .X(net816));
 sky130_fd_sc_hd__buf_2 rebuffer342 (.A(_08497_),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer343 (.A(net817),
    .X(net818));
 sky130_fd_sc_hd__buf_4 rebuffer344 (.A(net818),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer345 (.A(net819),
    .X(net820));
 sky130_fd_sc_hd__buf_6 rebuffer346 (.A(\id_stage_i.controller_i.instr_i[31] ),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer347 (.A(net821),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer348 (.A(net821),
    .X(net823));
 sky130_fd_sc_hd__buf_6 rebuffer349 (.A(net823),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer350 (.A(net824),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer351 (.A(net824),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer352 (.A(net826),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer353 (.A(net827),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer354 (.A(net827),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer355 (.A(net829),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer356 (.A(net823),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer357 (.A(net821),
    .X(net832));
 sky130_fd_sc_hd__buf_4 rebuffer358 (.A(net848),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer359 (.A(net833),
    .X(net834));
 sky130_fd_sc_hd__buf_6 rebuffer360 (.A(_09675_),
    .X(net835));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer361 (.A(net835),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer362 (.A(net836),
    .X(net837));
 sky130_fd_sc_hd__buf_6 rebuffer363 (.A(net837),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer364 (.A(_08630_),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer365 (.A(\id_stage_i.controller_i.instr_i[3] ),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer366 (.A(net840),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer367 (.A(\id_stage_i.controller_i.instr_i[3] ),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer368 (.A(net842),
    .X(net843));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer369 (.A(\id_stage_i.controller_i.instr_i[3] ),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer370 (.A(net844),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer371 (.A(net845),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer372 (.A(net844),
    .X(net847));
 sky130_fd_sc_hd__clkbuf_2 rebuffer373 (.A(_09445_),
    .X(net848));
 sky130_fd_sc_hd__buf_6 rebuffer374 (.A(_09445_),
    .X(net849));
 sky130_fd_sc_hd__buf_6 rebuffer375 (.A(_10665_),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer376 (.A(net850),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer377 (.A(net850),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer378 (.A(net440),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer379 (.A(net853),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer380 (.A(net1293),
    .X(net855));
 sky130_fd_sc_hd__clkbuf_16 clone381 (.A(net427),
    .X(net856));
 sky130_fd_sc_hd__a21o_2 clone382 (.A1(net658),
    .A2(_01712_),
    .B1(net1268),
    .X(net857));
 sky130_fd_sc_hd__buf_2 rebuffer383 (.A(_03963_),
    .X(net858));
 sky130_fd_sc_hd__a31oi_4 clone384 (.A1(net686),
    .A2(net266),
    .A3(_05186_),
    .B1(_05190_),
    .Y(net859));
 sky130_fd_sc_hd__buf_6 rebuffer385 (.A(_05167_),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer386 (.A(_08967_),
    .X(net861));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer387 (.A(_08599_),
    .X(net862));
 sky130_fd_sc_hd__buf_4 rebuffer388 (.A(net862),
    .X(net863));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer389 (.A(net863),
    .X(net864));
 sky130_fd_sc_hd__clkbuf_16 clone390 (.A(net963),
    .X(net865));
 sky130_fd_sc_hd__buf_6 rebuffer391 (.A(_08469_),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer392 (.A(net866),
    .X(net867));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer393 (.A(net866),
    .X(net868));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer394 (.A(net868),
    .X(net869));
 sky130_fd_sc_hd__buf_4 rebuffer395 (.A(_08469_),
    .X(net870));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer396 (.A(net870),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer397 (.A(net870),
    .X(net872));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer398 (.A(net870),
    .X(net873));
 sky130_fd_sc_hd__nor3_4 clone399 (.A(_04397_),
    .B(_04406_),
    .C(net1262),
    .Y(net874));
 sky130_fd_sc_hd__buf_6 rebuffer400 (.A(_08610_),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer401 (.A(net875),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer402 (.A(_09357_),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer403 (.A(net877),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer404 (.A(_09357_),
    .X(net879));
 sky130_fd_sc_hd__clkbuf_2 rebuffer405 (.A(_09053_),
    .X(net880));
 sky130_fd_sc_hd__buf_2 rebuffer406 (.A(net880),
    .X(net881));
 sky130_fd_sc_hd__buf_2 rebuffer407 (.A(net1223),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer408 (.A(_09054_),
    .X(net883));
 sky130_fd_sc_hd__buf_6 rebuffer409 (.A(_10436_),
    .X(net884));
 sky130_fd_sc_hd__clkbuf_16 clone410 (.A(net1296),
    .X(net885));
 sky130_fd_sc_hd__buf_6 clone411 (.A(net1296),
    .X(net886));
 sky130_fd_sc_hd__or2_2 clone412 (.A(net1215),
    .B(_01976_),
    .X(net887));
 sky130_fd_sc_hd__clkbuf_2 rebuffer413 (.A(_02797_),
    .X(net888));
 sky130_fd_sc_hd__clkbuf_2 rebuffer414 (.A(_08453_),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer415 (.A(net889),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer416 (.A(net889),
    .X(net891));
 sky130_fd_sc_hd__buf_6 rebuffer417 (.A(_08474_),
    .X(net892));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer418 (.A(net892),
    .X(net893));
 sky130_fd_sc_hd__buf_2 rebuffer419 (.A(net892),
    .X(net894));
 sky130_fd_sc_hd__buf_2 rebuffer420 (.A(_08474_),
    .X(net895));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer421 (.A(net895),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer422 (.A(net895),
    .X(net897));
 sky130_fd_sc_hd__nor2_4 clone423 (.A(_02300_),
    .B(_02299_),
    .Y(net898));
 sky130_fd_sc_hd__and2_2 clone424 (.A(_02931_),
    .B(net900),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer425 (.A(net1223),
    .X(net900));
 sky130_fd_sc_hd__clkbuf_16 clone426 (.A(net422),
    .X(net901));
 sky130_fd_sc_hd__buf_1 rebuffer427 (.A(net1174),
    .X(net902));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer428 (.A(_03177_),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer429 (.A(net984),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer430 (.A(net904),
    .X(net905));
 sky130_fd_sc_hd__buf_2 rebuffer431 (.A(_02308_),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer432 (.A(net906),
    .X(net907));
 sky130_fd_sc_hd__buf_2 rebuffer433 (.A(net906),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer434 (.A(net1286),
    .X(net909));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer435 (.A(net909),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer436 (.A(net910),
    .X(net911));
 sky130_fd_sc_hd__clkbuf_16 clone437 (.A(net1311),
    .X(net912));
 sky130_fd_sc_hd__buf_6 rebuffer438 (.A(_09085_),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer439 (.A(net913),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer440 (.A(net913),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer441 (.A(_09413_),
    .X(net916));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer442 (.A(\id_stage_i.controller_i.instr_i[30] ),
    .X(net917));
 sky130_fd_sc_hd__buf_2 rebuffer443 (.A(net917),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer444 (.A(net918),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer445 (.A(net919),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer446 (.A(net920),
    .X(net921));
 sky130_fd_sc_hd__buf_2 rebuffer447 (.A(net917),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer448 (.A(net917),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer449 (.A(net917),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer450 (.A(_09149_),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer451 (.A(net925),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer452 (.A(net926),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer453 (.A(net925),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer454 (.A(_01966_),
    .X(net929));
 sky130_fd_sc_hd__clkbuf_2 rebuffer455 (.A(net1281),
    .X(net930));
 sky130_fd_sc_hd__buf_6 rebuffer456 (.A(_09331_),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer457 (.A(net931),
    .X(net932));
 sky130_fd_sc_hd__nand3_2 clone458 (.A(net1034),
    .B(_08306_),
    .C(_08300_),
    .Y(net933));
 sky130_fd_sc_hd__buf_2 rebuffer459 (.A(_08901_),
    .X(net934));
 sky130_fd_sc_hd__buf_1 rebuffer460 (.A(net934),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer461 (.A(_02715_),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer462 (.A(_10331_),
    .X(net937));
 sky130_fd_sc_hd__clkbuf_16 clone463 (.A(net1012),
    .X(net938));
 sky130_fd_sc_hd__nor2_4 clone464 (.A(net1166),
    .B(net1058),
    .Y(net939));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer465 (.A(_08370_),
    .X(net940));
 sky130_fd_sc_hd__buf_6 rebuffer466 (.A(_08370_),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer467 (.A(net941),
    .X(net942));
 sky130_fd_sc_hd__buf_2 rebuffer468 (.A(net941),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer469 (.A(net943),
    .X(net944));
 sky130_fd_sc_hd__buf_6 rebuffer470 (.A(_01717_),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer471 (.A(net945),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer472 (.A(net945),
    .X(net947));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer473 (.A(net945),
    .X(net948));
 sky130_fd_sc_hd__buf_4 rebuffer474 (.A(net948),
    .X(net949));
 sky130_fd_sc_hd__buf_1 rebuffer475 (.A(net949),
    .X(net950));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer476 (.A(net950),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer477 (.A(_09111_),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer478 (.A(net952),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer479 (.A(net1506),
    .X(net954));
 sky130_fd_sc_hd__clkbuf_2 rebuffer480 (.A(_08590_),
    .X(net955));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer481 (.A(net955),
    .X(net956));
 sky130_fd_sc_hd__clkbuf_16 clone482 (.A(_05261_),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer483 (.A(_02057_),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer484 (.A(_02512_),
    .X(net959));
 sky130_fd_sc_hd__buf_12 rebuffer485 (.A(_09895_),
    .X(net960));
 sky130_fd_sc_hd__buf_6 rebuffer486 (.A(net960),
    .X(net961));
 sky130_fd_sc_hd__clkbuf_16 clone487 (.A(net437),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer488 (.A(net1147),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer489 (.A(net1191),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer490 (.A(\id_stage_i.controller_i.instr_i[12] ),
    .X(net965));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer491 (.A(\id_stage_i.controller_i.instr_i[12] ),
    .X(net966));
 sky130_fd_sc_hd__buf_6 rebuffer492 (.A(\id_stage_i.controller_i.instr_i[12] ),
    .X(net967));
 sky130_fd_sc_hd__buf_6 rebuffer493 (.A(net967),
    .X(net968));
 sky130_fd_sc_hd__buf_1 rebuffer494 (.A(net968),
    .X(net969));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer495 (.A(net968),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer496 (.A(net968),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer497 (.A(net968),
    .X(net972));
 sky130_fd_sc_hd__buf_2 rebuffer498 (.A(net967),
    .X(net973));
 sky130_fd_sc_hd__o22a_2 clone499 (.A1(_08639_),
    .A2(_08703_),
    .B1(net308),
    .B2(_08436_),
    .X(net974));
 sky130_fd_sc_hd__bufbuf_16 rebuffer500 (.A(net392),
    .X(net975));
 sky130_fd_sc_hd__buf_2 rebuffer501 (.A(net975),
    .X(net976));
 sky130_fd_sc_hd__buf_6 rebuffer502 (.A(net975),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer503 (.A(net975),
    .X(net978));
 sky130_fd_sc_hd__o211ai_2 clone504 (.A1(_09684_),
    .A2(_09686_),
    .B1(_09706_),
    .C1(net1056),
    .Y(net979));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer505 (.A(_08994_),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer506 (.A(_08995_),
    .X(net981));
 sky130_fd_sc_hd__buf_2 rebuffer507 (.A(_08995_),
    .X(net982));
 sky130_fd_sc_hd__clkbuf_16 clone508 (.A(net1029),
    .X(net983));
 sky130_fd_sc_hd__a21oi_2 clone509 (.A1(_01712_),
    .A2(net660),
    .B1(net1268),
    .Y(net984));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer510 (.A(_08978_),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer511 (.A(_08986_),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer512 (.A(_09039_),
    .X(net987));
 sky130_fd_sc_hd__clkbuf_16 clone513 (.A(net365),
    .X(net988));
 sky130_fd_sc_hd__clkbuf_16 clone514 (.A(net1162),
    .X(net989));
 sky130_fd_sc_hd__a22o_4 clone515 (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .A2(net991),
    .B1(_07641_),
    .B2(_11139_),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer516 (.A(_07636_),
    .X(net991));
 sky130_fd_sc_hd__buf_2 rebuffer517 (.A(net163),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer518 (.A(net992),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer519 (.A(\id_stage_i.controller_i.instr_i[5] ),
    .X(net994));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer520 (.A(\id_stage_i.controller_i.instr_i[5] ),
    .X(net995));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer521 (.A(net995),
    .X(net996));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer522 (.A(net996),
    .X(net997));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer523 (.A(net997),
    .X(net998));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer524 (.A(net996),
    .X(net999));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer525 (.A(\id_stage_i.controller_i.instr_i[5] ),
    .X(net1000));
 sky130_fd_sc_hd__buf_6 rebuffer526 (.A(_09174_),
    .X(net1001));
 sky130_fd_sc_hd__buf_6 rebuffer527 (.A(net1276),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer528 (.A(_08597_),
    .X(net1003));
 sky130_fd_sc_hd__and2_2 clone529 (.A(net1035),
    .B(_02503_),
    .X(net1004));
 sky130_fd_sc_hd__xnor3_2 clone530 (.A(_02493_),
    .B(_02496_),
    .C(_02531_),
    .X(net1005));
 sky130_fd_sc_hd__clkbuf_2 rebuffer531 (.A(_02132_),
    .X(net1006));
 sky130_fd_sc_hd__buf_4 rebuffer532 (.A(net161),
    .X(net1007));
 sky130_fd_sc_hd__clkbuf_16 clone533 (.A(net423),
    .X(net1008));
 sky130_fd_sc_hd__clkbuf_16 clone534 (.A(net1070),
    .X(net1009));
 sky130_fd_sc_hd__nand2_4 clone535 (.A(net1011),
    .B(_02424_),
    .Y(net1010));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer536 (.A(_02425_),
    .X(net1011));
 sky130_fd_sc_hd__buf_6 clone537 (.A(net425),
    .X(net1012));
 sky130_fd_sc_hd__clkbuf_16 clone538 (.A(net1015),
    .X(net1013));
 sky130_fd_sc_hd__buf_12 rebuffer539 (.A(_08457_),
    .X(net1014));
 sky130_fd_sc_hd__buf_2 rebuffer540 (.A(net1014),
    .X(net1015));
 sky130_fd_sc_hd__clkbuf_16 clone541 (.A(net426),
    .X(net1016));
 sky130_fd_sc_hd__buf_6 clone554 (.A(net653),
    .X(net1029));
 sky130_fd_sc_hd__buf_6 clone555 (.A(net363),
    .X(net1030));
 sky130_fd_sc_hd__clkbuf_16 clone595 (.A(net1114),
    .X(net1070));
 sky130_fd_sc_hd__buf_6 rebuffer596 (.A(_10478_),
    .X(net1071));
 sky130_fd_sc_hd__clkbuf_16 clone597 (.A(net415),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer598 (.A(_08520_),
    .X(net1073));
 sky130_fd_sc_hd__clkbuf_16 clone599 (.A(net433),
    .X(net1074));
 sky130_fd_sc_hd__clkbuf_16 clone600 (.A(net1152),
    .X(net1075));
 sky130_fd_sc_hd__clkbuf_16 clone601 (.A(net427),
    .X(net1076));
 sky130_fd_sc_hd__clkbuf_16 clone602 (.A(net366),
    .X(net1077));
 sky130_fd_sc_hd__clkbuf_16 clone603 (.A(net408),
    .X(net1078));
 sky130_fd_sc_hd__buf_6 rebuffer604 (.A(_09405_),
    .X(net1079));
 sky130_fd_sc_hd__clkbuf_16 clone605 (.A(net1147),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer606 (.A(_10259_),
    .X(net1081));
 sky130_fd_sc_hd__clkbuf_16 clone607 (.A(net388),
    .X(net1082));
 sky130_fd_sc_hd__clkbuf_16 clone608 (.A(net1112),
    .X(net1083));
 sky130_fd_sc_hd__clkbuf_16 clone609 (.A(net1147),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer610 (.A(_08950_),
    .X(net1085));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer611 (.A(\id_stage_i.controller_i.instr_i[14] ),
    .X(net1086));
 sky130_fd_sc_hd__buf_6 rebuffer612 (.A(\id_stage_i.controller_i.instr_i[14] ),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer613 (.A(net1087),
    .X(net1088));
 sky130_fd_sc_hd__buf_6 rebuffer614 (.A(net1087),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer615 (.A(net1089),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer616 (.A(net1090),
    .X(net1091));
 sky130_fd_sc_hd__buf_1 rebuffer617 (.A(net1089),
    .X(net1092));
 sky130_fd_sc_hd__clkbuf_16 clone618 (.A(net358),
    .X(net1093));
 sky130_fd_sc_hd__buf_6 rebuffer619 (.A(\id_stage_i.controller_i.instr_i[6] ),
    .X(net1094));
 sky130_fd_sc_hd__buf_4 rebuffer620 (.A(net1094),
    .X(net1095));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer621 (.A(net1095),
    .X(net1096));
 sky130_fd_sc_hd__buf_2 rebuffer622 (.A(\id_stage_i.controller_i.instr_i[6] ),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer623 (.A(net1097),
    .X(net1098));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer624 (.A(net1097),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer625 (.A(net1099),
    .X(net1100));
 sky130_fd_sc_hd__buf_2 rebuffer626 (.A(_08586_),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer627 (.A(net1101),
    .X(net1102));
 sky130_fd_sc_hd__buf_6 rebuffer628 (.A(_08586_),
    .X(net1103));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer629 (.A(net1103),
    .X(net1104));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer630 (.A(net1103),
    .X(net1105));
 sky130_fd_sc_hd__buf_6 rebuffer631 (.A(net1103),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer632 (.A(net1103),
    .X(net1107));
 sky130_fd_sc_hd__clkbuf_16 clone633 (.A(net389),
    .X(net1108));
 sky130_fd_sc_hd__buf_2 rebuffer634 (.A(net418),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer635 (.A(_08957_),
    .X(net1110));
 sky130_fd_sc_hd__clkbuf_16 clone636 (.A(net1130),
    .X(net1111));
 sky130_fd_sc_hd__clkbuf_16 clone637 (.A(net411),
    .X(net1112));
 sky130_fd_sc_hd__clkbuf_16 clone638 (.A(net1114),
    .X(net1113));
 sky130_fd_sc_hd__clkbuf_2 rebuffer639 (.A(net414),
    .X(net1114));
 sky130_fd_sc_hd__buf_4 rebuffer640 (.A(_08307_),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer641 (.A(net1115),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer642 (.A(net1115),
    .X(net1117));
 sky130_fd_sc_hd__buf_6 rebuffer643 (.A(_08613_),
    .X(net1118));
 sky130_fd_sc_hd__clkbuf_16 clone644 (.A(net1014),
    .X(net1119));
 sky130_fd_sc_hd__clkbuf_16 clone645 (.A(net367),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer646 (.A(_09283_),
    .X(net1121));
 sky130_fd_sc_hd__clkbuf_16 clone647 (.A(net1123),
    .X(net1122));
 sky130_fd_sc_hd__clkbuf_16 clone648 (.A(net437),
    .X(net1123));
 sky130_fd_sc_hd__buf_6 rebuffer649 (.A(\id_stage_i.controller_i.instr_i[4] ),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer650 (.A(net1124),
    .X(net1125));
 sky130_fd_sc_hd__buf_2 rebuffer651 (.A(net1125),
    .X(net1126));
 sky130_fd_sc_hd__buf_4 rebuffer652 (.A(\id_stage_i.controller_i.instr_i[4] ),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer653 (.A(net1127),
    .X(net1128));
 sky130_fd_sc_hd__clkbuf_16 clone654 (.A(net1130),
    .X(net1129));
 sky130_fd_sc_hd__clkbuf_16 clone655 (.A(net439),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer656 (.A(_08694_),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer657 (.A(net1131),
    .X(net1132));
 sky130_fd_sc_hd__clkbuf_16 clone658 (.A(net1154),
    .X(net1133));
 sky130_fd_sc_hd__or3_2 clone659 (.A(_08293_),
    .B(_08294_),
    .C(_08265_),
    .X(net1134));
 sky130_fd_sc_hd__clkbuf_16 clone660 (.A(net418),
    .X(net1135));
 sky130_fd_sc_hd__buf_1 rebuffer661 (.A(_09333_),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer662 (.A(net1136),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer663 (.A(net1136),
    .X(net1138));
 sky130_fd_sc_hd__buf_2 rebuffer664 (.A(_09333_),
    .X(net1139));
 sky130_fd_sc_hd__clkbuf_16 clone665 (.A(net390),
    .X(net1140));
 sky130_fd_sc_hd__clkbuf_16 clone666 (.A(net365),
    .X(net1141));
 sky130_fd_sc_hd__clkbuf_16 clone667 (.A(net1148),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer668 (.A(_09222_),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer669 (.A(_09606_),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer670 (.A(_09414_),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer671 (.A(net1145),
    .X(net1146));
 sky130_fd_sc_hd__clkbuf_16 clone672 (.A(net1162),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer673 (.A(net511),
    .X(net1148));
 sky130_fd_sc_hd__clkbuf_16 clone674 (.A(net1151),
    .X(net1149));
 sky130_fd_sc_hd__buf_4 rebuffer675 (.A(_08799_),
    .X(net1150));
 sky130_fd_sc_hd__buf_1 rebuffer676 (.A(_08799_),
    .X(net1151));
 sky130_fd_sc_hd__clkbuf_16 clone677 (.A(net392),
    .X(net1152));
 sky130_fd_sc_hd__and2_4 clone678 (.A(net343),
    .B(net810),
    .X(net1153));
 sky130_fd_sc_hd__clkbuf_16 clone679 (.A(net381),
    .X(net1154));
 sky130_fd_sc_hd__buf_2 rebuffer685 (.A(_03148_),
    .X(net1160));
 sky130_fd_sc_hd__mux2_4 clone686 (.A0(net1184),
    .A1(net1211),
    .S(net322),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer687 (.A(net440),
    .X(net1162));
 sky130_fd_sc_hd__buf_6 rebuffer688 (.A(_10762_),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer689 (.A(net1163),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer690 (.A(net1163),
    .X(net1165));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer691 (.A(_01991_),
    .X(net1166));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer692 (.A(net1182),
    .X(net1167));
 sky130_fd_sc_hd__buf_2 rebuffer693 (.A(net1167),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer694 (.A(net1168),
    .X(net1169));
 sky130_fd_sc_hd__buf_1 rebuffer695 (.A(_02132_),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer696 (.A(_02132_),
    .X(net1171));
 sky130_fd_sc_hd__and2_2 clone697 (.A(_01966_),
    .B(net1200),
    .X(net1172));
 sky130_fd_sc_hd__a21o_4 clone698 (.A1(_02619_),
    .A2(_01712_),
    .B1(net1293),
    .X(net1173));
 sky130_fd_sc_hd__buf_6 rebuffer699 (.A(_10102_),
    .X(net1174));
 sky130_fd_sc_hd__clkbuf_16 clone700 (.A(net430),
    .X(net1175));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer701 (.A(net1155),
    .X(net1176));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer702 (.A(net1156),
    .X(net1177));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer703 (.A(net1155),
    .X(net1178));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer704 (.A(net1178),
    .X(net1179));
 sky130_fd_sc_hd__buf_6 rebuffer705 (.A(_02132_),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer706 (.A(net1180),
    .X(net1181));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer707 (.A(net1181),
    .X(net1182));
 sky130_fd_sc_hd__buf_1 rebuffer708 (.A(_03013_),
    .X(net1183));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer709 (.A(_09217_),
    .X(net1184));
 sky130_fd_sc_hd__clkbuf_16 clone710 (.A(net408),
    .X(net1185));
 sky130_fd_sc_hd__clkbuf_16 clone726 (.A(net1203),
    .X(net1201));
 sky130_fd_sc_hd__buf_2 rebuffer727 (.A(_08453_),
    .X(net1202));
 sky130_fd_sc_hd__buf_2 rebuffer728 (.A(net1202),
    .X(net1203));
 sky130_fd_sc_hd__clkbuf_16 clone729 (.A(net1234),
    .X(net1204));
 sky130_fd_sc_hd__buf_6 rebuffer730 (.A(_03375_),
    .X(net1205));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer731 (.A(net1205),
    .X(net1206));
 sky130_fd_sc_hd__buf_4 rebuffer732 (.A(net1206),
    .X(net1207));
 sky130_fd_sc_hd__nand2_4 clone741 (.A(net1036),
    .B(_02424_),
    .Y(net1216));
 sky130_fd_sc_hd__buf_6 rebuffer742 (.A(_10201_),
    .X(net1217));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer743 (.A(net1217),
    .X(net1218));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer744 (.A(_02525_),
    .X(net1219));
 sky130_fd_sc_hd__buf_6 clone745 (.A(net380),
    .X(net1220));
 sky130_fd_sc_hd__clkbuf_2 rebuffer750 (.A(net391),
    .X(net1225));
 sky130_fd_sc_hd__buf_12 rebuffer751 (.A(_08324_),
    .X(net1226));
 sky130_fd_sc_hd__buf_6 rebuffer752 (.A(_08324_),
    .X(net1227));
 sky130_fd_sc_hd__nand4_2 clone753 (.A(_02391_),
    .B(_02392_),
    .C(net1025),
    .D(_02395_),
    .Y(net1228));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer754 (.A(_10915_),
    .X(net1229));
 sky130_fd_sc_hd__buf_6 rebuffer755 (.A(net1229),
    .X(net1230));
 sky130_fd_sc_hd__buf_6 rebuffer756 (.A(net1230),
    .X(net1231));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer757 (.A(net1231),
    .X(net1232));
 sky130_fd_sc_hd__clkbuf_16 clone758 (.A(net1234),
    .X(net1233));
 sky130_fd_sc_hd__buf_4 rebuffer759 (.A(net410),
    .X(net1234));
 sky130_fd_sc_hd__buf_4 rebuffer760 (.A(net411),
    .X(net1235));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer761 (.A(_10272_),
    .X(net1236));
 sky130_fd_sc_hd__buf_12 rebuffer762 (.A(_05191_),
    .X(net1237));
 sky130_fd_sc_hd__clkbuf_16 clone763 (.A(_05191_),
    .X(net1238));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer764 (.A(net1335),
    .X(net1239));
 sky130_fd_sc_hd__dlymetal6s4s_1 rebuffer765 (.A(net1239),
    .X(net1240));
 sky130_fd_sc_hd__buf_12 rebuffer766 (.A(net159),
    .X(net1241));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer767 (.A(net1241),
    .X(net1242));
 sky130_fd_sc_hd__buf_4 rebuffer769 (.A(net164),
    .X(net1244));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer770 (.A(net164),
    .X(net1245));
 sky130_fd_sc_hd__o221ai_4 clone771 (.A1(_05060_),
    .A2(net1505),
    .B1(_05061_),
    .B2(_05078_),
    .C1(net265),
    .Y(net1246));
 sky130_fd_sc_hd__buf_2 rebuffer772 (.A(_08344_),
    .X(net1247));
 sky130_fd_sc_hd__and2_2 clone773 (.A(net1225),
    .B(net394),
    .X(net1248));
 sky130_fd_sc_hd__o221ai_4 clone774 (.A1(_05060_),
    .A2(net1505),
    .B1(_05061_),
    .B2(_05078_),
    .C1(net265),
    .Y(net1249));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer775 (.A(_05577_),
    .X(net1250));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer776 (.A(_05577_),
    .X(net1251));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer777 (.A(_05577_),
    .X(net1252));
 sky130_fd_sc_hd__buf_6 rebuffer778 (.A(_05577_),
    .X(net1253));
 sky130_fd_sc_hd__o221ai_4 clone779 (.A1(_05060_),
    .A2(net1505),
    .B1(_05061_),
    .B2(_05078_),
    .C1(net265),
    .Y(net1254));
 sky130_fd_sc_hd__clkbuf_2 rebuffer780 (.A(net162),
    .X(net1255));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer781 (.A(net1255),
    .X(net1256));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer782 (.A(net1255),
    .X(net1257));
 sky130_fd_sc_hd__buf_6 rebuffer783 (.A(net1257),
    .X(net1258));
 sky130_fd_sc_hd__buf_12 rebuffer784 (.A(net162),
    .X(net1259));
 sky130_fd_sc_hd__buf_12 rebuffer785 (.A(net160),
    .X(net1260));
 sky130_fd_sc_hd__buf_2 rebuffer786 (.A(net1260),
    .X(net1261));
 sky130_fd_sc_hd__buf_6 rebuffer787 (.A(_04534_),
    .X(net1262));
 sky130_fd_sc_hd__buf_6 rebuffer795 (.A(net874),
    .X(net1270));
 sky130_fd_sc_hd__buf_6 rebuffer796 (.A(net874),
    .X(net1271));
 sky130_fd_sc_hd__buf_12 rebuffer798 (.A(net155),
    .X(net1273));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer799 (.A(net1273),
    .X(net1274));
 sky130_fd_sc_hd__a31oi_4 clone813 (.A1(_02646_),
    .A2(_03478_),
    .A3(_04256_),
    .B1(net1289),
    .Y(net1288));
 sky130_fd_sc_hd__buf_8 rebuffer814 (.A(_04389_),
    .X(net1289));
 sky130_fd_sc_hd__buf_6 rebuffer815 (.A(net1288),
    .X(net1290));
 sky130_fd_sc_hd__buf_12 rebuffer816 (.A(net1288),
    .X(net1291));
 sky130_fd_sc_hd__nor3_2 clone817 (.A(_11164_),
    .B(_07635_),
    .C(_11201_),
    .Y(net1292));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer818 (.A(_02621_),
    .X(net1293));
 sky130_fd_sc_hd__clkbuf_16 clone819 (.A(net1296),
    .X(net1294));
 sky130_fd_sc_hd__buf_2 rebuffer820 (.A(_04975_),
    .X(net1295));
 sky130_fd_sc_hd__buf_6 rebuffer821 (.A(_04975_),
    .X(net1296));
 sky130_fd_sc_hd__nand3_4 clone825 (.A(net1020),
    .B(net331),
    .C(net1325),
    .Y(net1300));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer848 (.A(_05956_),
    .X(net1323));
 sky130_fd_sc_hd__buf_6 rebuffer849 (.A(_05956_),
    .X(net1324));
 sky130_fd_sc_hd__buf_4 rebuffer850 (.A(net1324),
    .X(net1325));
 sky130_fd_sc_hd__o31a_4 clone851 (.A1(_11641_),
    .A2(_02646_),
    .A3(_04248_),
    .B1(_04251_),
    .X(net1326));
 sky130_fd_sc_hd__o31a_4 clone852 (.A1(_11641_),
    .A2(_02646_),
    .A3(_04248_),
    .B1(_04251_),
    .X(net1327));
 sky130_fd_sc_hd__nor2_4 clone853 (.A(_11201_),
    .B(_11164_),
    .Y(net1328));
 sky130_fd_sc_hd__buf_12 load_slew1 (.A(net1585),
    .X(net1017));
 sky130_fd_sc_hd__buf_12 load_slew2 (.A(_13251_),
    .X(net1018));
 sky130_fd_sc_hd__clkbuf_4 wire3 (.A(_11348_),
    .X(net1019));
 sky130_fd_sc_hd__buf_16 load_slew4 (.A(net1021),
    .X(net1020));
 sky130_fd_sc_hd__buf_16 wire5 (.A(\gen_regfile_ff.register_file_i.waddr_a_i[1] ),
    .X(net1021));
 sky130_fd_sc_hd__buf_12 rebuffer16 (.A(_09157_),
    .X(net1022));
 sky130_fd_sc_hd__buf_2 rebuffer25 (.A(_09157_),
    .X(net1023));
 sky130_fd_sc_hd__and2_4 clone26 (.A(net343),
    .B(net810),
    .X(net1024));
 sky130_fd_sc_hd__buf_2 rebuffer89 (.A(_02393_),
    .X(net1025));
 sky130_fd_sc_hd__a2111o_2 clone91 (.A1(_10996_),
    .A2(_11004_),
    .B1(_11042_),
    .C1(_11034_),
    .D1(_11011_),
    .X(net1026));
 sky130_fd_sc_hd__buf_2 rebuffer174 (.A(_02396_),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer175 (.A(net1027),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer177 (.A(net1027),
    .X(net1031));
 sky130_fd_sc_hd__buf_6 rebuffer210 (.A(\id_stage_i.controller_i.instr_i[25] ),
    .X(net1032));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer223 (.A(net1032),
    .X(net1033));
 sky130_fd_sc_hd__buf_2 rebuffer224 (.A(_08299_),
    .X(net1034));
 sky130_fd_sc_hd__buf_12 rebuffer264 (.A(_02502_),
    .X(net1035));
 sky130_fd_sc_hd__buf_6 rebuffer306 (.A(_02425_),
    .X(net1036));
 sky130_fd_sc_hd__clkbuf_2 rebuffer319 (.A(_09159_),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer324 (.A(net1037),
    .X(net1038));
 sky130_fd_sc_hd__a22o_4 clone325 (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .A2(net1292),
    .B1(_11139_),
    .B2(_07641_),
    .X(net1039));
 sky130_fd_sc_hd__buf_2 rebuffer381 (.A(net176),
    .X(net1040));
 sky130_fd_sc_hd__buf_6 rebuffer382 (.A(_10535_),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer384 (.A(net1041),
    .X(net1042));
 sky130_fd_sc_hd__buf_6 rebuffer390 (.A(_08464_),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer399 (.A(net1043),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer410 (.A(net1043),
    .X(net1045));
 sky130_fd_sc_hd__buf_8 rebuffer411 (.A(net1043),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer412 (.A(net1046),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer423 (.A(_08405_),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer424 (.A(_09928_),
    .X(net1049));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer426 (.A(_01992_),
    .X(net1050));
 sky130_fd_sc_hd__buf_6 rebuffer437 (.A(_02003_),
    .X(net1051));
 sky130_fd_sc_hd__buf_2 rebuffer458 (.A(_02003_),
    .X(net1052));
 sky130_fd_sc_hd__buf_6 rebuffer463 (.A(_02003_),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer464 (.A(net1053),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer482 (.A(net1053),
    .X(net1055));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer487 (.A(_09699_),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer499 (.A(_01990_),
    .X(net1057));
 sky130_fd_sc_hd__buf_4 rebuffer504 (.A(net1057),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer508 (.A(\gen_regfile_ff.register_file_i.raddr_b_i[0] ),
    .X(net1059));
 sky130_fd_sc_hd__buf_2 rebuffer509 (.A(_01992_),
    .X(net1060));
 sky130_fd_sc_hd__nand2_8 clone510 (.A(_07639_),
    .B(_07640_),
    .Y(net1061));
 sky130_fd_sc_hd__xnor2_2 clone511 (.A(_10959_),
    .B(_09118_),
    .Y(net1062));
 sky130_fd_sc_hd__buf_12 rebuffer513 (.A(_03118_),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer514 (.A(net1063),
    .X(net1064));
 sky130_fd_sc_hd__buf_12 rebuffer515 (.A(_09303_),
    .X(net1065));
 sky130_fd_sc_hd__clkbuf_2 rebuffer529 (.A(net1065),
    .X(net1066));
 sky130_fd_sc_hd__clkbuf_2 rebuffer530 (.A(_02138_),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer533 (.A(_02138_),
    .X(net1068));
 sky130_fd_sc_hd__buf_6 rebuffer534 (.A(_02331_),
    .X(net1069));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer535 (.A(_01725_),
    .X(net1155));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer537 (.A(net1155),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer538 (.A(_02725_),
    .X(net1157));
 sky130_fd_sc_hd__or2_2 clone539 (.A(_02725_),
    .B(_02723_),
    .X(net1158));
 sky130_fd_sc_hd__clkbuf_2 rebuffer541 (.A(_02599_),
    .X(net1159));
 sky130_fd_sc_hd__clkbuf_16 clone542 (.A(net480),
    .X(net1186));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer543 (.A(_09349_),
    .X(net1187));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer544 (.A(net1187),
    .X(net1188));
 sky130_fd_sc_hd__buf_6 rebuffer545 (.A(net1188),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer546 (.A(_01711_),
    .X(net1190));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer547 (.A(_08745_),
    .X(net1191));
 sky130_fd_sc_hd__buf_2 rebuffer548 (.A(_02622_),
    .X(net1192));
 sky130_fd_sc_hd__buf_1 rebuffer549 (.A(_02622_),
    .X(net1193));
 sky130_fd_sc_hd__a21o_2 clone550 (.A1(_02619_),
    .A2(_01712_),
    .B1(_02621_),
    .X(net1194));
 sky130_fd_sc_hd__buf_4 rebuffer551 (.A(_08187_),
    .X(net1195));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer552 (.A(net1195),
    .X(net1196));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer553 (.A(net1195),
    .X(net1197));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer554 (.A(net1195),
    .X(net1198));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer555 (.A(net1195),
    .X(net1199));
 sky130_fd_sc_hd__buf_4 rebuffer556 (.A(_01970_),
    .X(net1200));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer557 (.A(net1200),
    .X(net1208));
 sky130_fd_sc_hd__buf_2 rebuffer558 (.A(_01980_),
    .X(net1209));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer559 (.A(_08910_),
    .X(net1210));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer560 (.A(_10392_),
    .X(net1211));
 sky130_fd_sc_hd__buf_2 rebuffer561 (.A(_10392_),
    .X(net1212));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer562 (.A(_02730_),
    .X(net1213));
 sky130_fd_sc_hd__clkbuf_4 rebuffer563 (.A(_01977_),
    .X(net1214));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer564 (.A(net1214),
    .X(net1215));
 sky130_fd_sc_hd__buf_6 rebuffer565 (.A(_02773_),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer566 (.A(net1221),
    .X(net1222));
 sky130_fd_sc_hd__buf_6 rebuffer567 (.A(_02930_),
    .X(net1223));
 sky130_fd_sc_hd__buf_4 rebuffer568 (.A(_01978_),
    .X(net1224));
 sky130_fd_sc_hd__buf_4 rebuffer569 (.A(_03165_),
    .X(net1243));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer570 (.A(net1243),
    .X(net1263));
 sky130_fd_sc_hd__buf_2 rebuffer571 (.A(net1263),
    .X(net1264));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer572 (.A(net1264),
    .X(net1265));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer573 (.A(net1265),
    .X(net1266));
 sky130_fd_sc_hd__buf_1 rebuffer574 (.A(_02746_),
    .X(net1267));
 sky130_fd_sc_hd__and4b_2 clone575 (.A_N(_09763_),
    .B(net1269),
    .C(_09783_),
    .D(net321),
    .X(net1268));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer576 (.A(net1304),
    .X(net1269));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer577 (.A(_09784_),
    .X(net1272));
 sky130_fd_sc_hd__buf_1 rebuffer578 (.A(_02630_),
    .X(net1275));
 sky130_fd_sc_hd__buf_2 rebuffer579 (.A(_08606_),
    .X(net1276));
 sky130_fd_sc_hd__buf_6 rebuffer580 (.A(_02504_),
    .X(net1277));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer581 (.A(_08752_),
    .X(net1278));
 sky130_fd_sc_hd__a21oi_2 clone582 (.A1(_01719_),
    .A2(_01720_),
    .B1(_01724_),
    .Y(net1279));
 sky130_fd_sc_hd__buf_8 rebuffer583 (.A(_08471_),
    .X(net1280));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer584 (.A(net1280),
    .X(net1281));
 sky130_fd_sc_hd__clkbuf_16 clone585 (.A(net390),
    .X(net1282));
 sky130_fd_sc_hd__clkbuf_16 clone586 (.A(net422),
    .X(net1283));
 sky130_fd_sc_hd__clkbuf_4 rebuffer587 (.A(net426),
    .X(net1284));
 sky130_fd_sc_hd__buf_12 rebuffer588 (.A(_08544_),
    .X(net1285));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer589 (.A(_02308_),
    .X(net1286));
 sky130_fd_sc_hd__nor2_4 clone590 (.A(net1214),
    .B(_01976_),
    .Y(net1287));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer591 (.A(_02435_),
    .X(net1297));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer592 (.A(_08159_),
    .X(net1298));
 sky130_fd_sc_hd__buf_4 rebuffer593 (.A(_08159_),
    .X(net1299));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer594 (.A(net1299),
    .X(net1301));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer595 (.A(net1301),
    .X(net1302));
 sky130_fd_sc_hd__a22o_4 clone596 (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .A2(net991),
    .B1(_07641_),
    .B2(_11139_),
    .X(net1303));
 sky130_fd_sc_hd__buf_6 rebuffer597 (.A(_09776_),
    .X(net1304));
 sky130_fd_sc_hd__nand2_4 clone598 (.A(_07639_),
    .B(_07640_),
    .Y(net1305));
 sky130_fd_sc_hd__buf_2 rebuffer599 (.A(_09051_),
    .X(net1306));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer600 (.A(_02301_),
    .X(net1307));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer601 (.A(net1307),
    .X(net1308));
 sky130_fd_sc_hd__clkbuf_16 clone604 (.A(net378),
    .X(net1309));
 sky130_fd_sc_hd__buf_6 clone606 (.A(net380),
    .X(net1310));
 sky130_fd_sc_hd__buf_2 rebuffer607 (.A(net431),
    .X(net1311));
 sky130_fd_sc_hd__clkbuf_16 clone610 (.A(net354),
    .X(net1312));
 sky130_fd_sc_hd__buf_12 rebuffer618 (.A(_10222_),
    .X(net1313));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer633 (.A(net1313),
    .X(net1314));
 sky130_fd_sc_hd__buf_6 rebuffer636 (.A(_04535_),
    .X(net1315));
 sky130_fd_sc_hd__buf_6 rebuffer637 (.A(net1315),
    .X(net1316));
 sky130_fd_sc_hd__buf_6 clone639 (.A(_04535_),
    .X(net1317));
 sky130_fd_sc_hd__buf_6 rebuffer666 (.A(_02800_),
    .X(net1335));
 sky130_fd_sc_hd__dlygate4sd3_1 rebuffer667 (.A(_02800_),
    .X(net1336));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer810 (.A(_02692_),
    .X(net1413));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer811 (.A(net1413),
    .X(net1414));
 sky130_fd_sc_hd__buf_12 rebuffer860 (.A(_08575_),
    .X(net1455));
 sky130_fd_sc_hd__buf_2 rebuffer861 (.A(net1455),
    .X(net1456));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer862 (.A(net1456),
    .X(net1457));
 sky130_fd_sc_hd__buf_6 rebuffer863 (.A(net1457),
    .X(net1458));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer864 (.A(net1458),
    .X(net1459));
 sky130_fd_sc_hd__a22o_4 clone865 (.A1(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .A2(net1292),
    .B1(_11139_),
    .B2(_07641_),
    .X(net1460));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer866 (.A(_08424_),
    .X(net1461));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer867 (.A(net1461),
    .X(net1462));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer868 (.A(_08424_),
    .X(net1463));
 sky130_fd_sc_hd__buf_1 rebuffer869 (.A(_10974_),
    .X(net1464));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer870 (.A(_09450_),
    .X(net1465));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer871 (.A(_10902_),
    .X(net1466));
 sky130_fd_sc_hd__buf_2 rebuffer872 (.A(net1466),
    .X(net1467));
 sky130_fd_sc_hd__buf_2 rebuffer873 (.A(net1466),
    .X(net1468));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer874 (.A(net1468),
    .X(net1469));
 sky130_fd_sc_hd__buf_12 rebuffer880 (.A(_04390_),
    .X(net1475));
 sky130_fd_sc_hd__clkbuf_16 clone881 (.A(net654),
    .X(net1476));
 sky130_fd_sc_hd__buf_2 rebuffer882 (.A(_05268_),
    .X(net1477));
 sky130_fd_sc_hd__buf_4 rebuffer883 (.A(net1477),
    .X(net1478));
 sky130_fd_sc_hd__buf_6 rebuffer884 (.A(net1477),
    .X(net1479));
 sky130_fd_sc_hd__nand3_4 clone885 (.A(_05847_),
    .B(_05796_),
    .C(net447),
    .Y(net1480));
 sky130_fd_sc_hd__nand3_4 clone886 (.A(_05847_),
    .B(_01919_),
    .C(net447),
    .Y(net1481));
 sky130_fd_sc_hd__nand3_4 clone887 (.A(_05847_),
    .B(_05955_),
    .C(net446),
    .Y(net1482));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer888 (.A(_01665_),
    .X(net1483));
 sky130_fd_sc_hd__buf_2 rebuffer889 (.A(net1483),
    .X(net1484));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer890 (.A(net1484),
    .X(net1485));
 sky130_fd_sc_hd__clkbuf_16 clone909 (.A(_04390_),
    .X(net1504));
 sky130_fd_sc_hd__buf_12 rebuffer910 (.A(_05059_),
    .X(net1505));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer911 (.A(_09111_),
    .X(net1506));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer915 (.A(_02917_),
    .X(net1510));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer916 (.A(_03584_),
    .X(net1511));
 sky130_fd_sc_hd__clkbuf_16 clone919 (.A(net1516),
    .X(net1514));
 sky130_fd_sc_hd__clkbuf_16 clone920 (.A(net1516),
    .X(net1515));
 sky130_fd_sc_hd__buf_12 rebuffer921 (.A(_04763_),
    .X(net1516));
 sky130_fd_sc_hd__o31a_4 clone922 (.A1(_11641_),
    .A2(_02646_),
    .A3(_04248_),
    .B1(_04251_),
    .X(net1517));
 sky130_fd_sc_hd__buf_2 rebuffer927 (.A(_03963_),
    .X(net1522));
 sky130_fd_sc_hd__buf_6 clone928 (.A(net1288),
    .X(net1523));
 sky130_fd_sc_hd__buf_2 rebuffer929 (.A(_08269_),
    .X(net1524));
 sky130_fd_sc_hd__buf_12 rebuffer930 (.A(net174),
    .X(net1525));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer931 (.A(net1525),
    .X(net1526));
 sky130_fd_sc_hd__or2_4 clone934 (.A(_04864_),
    .B(net1530),
    .X(net1529));
 sky130_fd_sc_hd__buf_12 rebuffer935 (.A(_04863_),
    .X(net1530));
 sky130_fd_sc_hd__or2_4 clone938 (.A(_04864_),
    .B(net1534),
    .X(net1533));
 sky130_fd_sc_hd__clkbuf_16 rebuffer939 (.A(_04863_),
    .X(net1534));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer940 (.A(net165),
    .X(net1535));
 sky130_fd_sc_hd__buf_12 clone941 (.A(net1516),
    .X(net1536));
 sky130_fd_sc_hd__a31oi_4 clone942 (.A1(_02646_),
    .A2(_03478_),
    .A3(_03871_),
    .B1(net1538),
    .Y(net1537));
 sky130_fd_sc_hd__buf_8 rebuffer943 (.A(_03981_),
    .X(net1538));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer944 (.A(net1533),
    .X(net1539));
 sky130_fd_sc_hd__buf_12 rebuffer945 (.A(net1533),
    .X(net1540));
 sky130_fd_sc_hd__buf_6 clone946 (.A(net1550),
    .X(net1541));
 sky130_fd_sc_hd__or2_4 clone947 (.A(_04864_),
    .B(net1530),
    .X(net1542));
 sky130_fd_sc_hd__buf_2 rebuffer948 (.A(net1024),
    .X(net1543));
 sky130_fd_sc_hd__a31oi_4 clone949 (.A1(_02646_),
    .A2(_03478_),
    .A3(_03871_),
    .B1(net1538),
    .Y(net1544));
 sky130_fd_sc_hd__buf_12 rebuffer952 (.A(net163),
    .X(net1547));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer953 (.A(net1547),
    .X(net1548));
 sky130_fd_sc_hd__clkbuf_2 rebuffer955 (.A(net874),
    .X(net1550));
 sky130_fd_sc_hd__a31oi_2 clone956 (.A1(_02646_),
    .A2(_03478_),
    .A3(_03744_),
    .B1(net1552),
    .Y(net1551));
 sky130_fd_sc_hd__buf_12 rebuffer957 (.A(_03865_),
    .X(net1552));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer958 (.A(_03865_),
    .X(net1553));
 sky130_fd_sc_hd__a2111o_2 clone959 (.A1(_10996_),
    .A2(_11004_),
    .B1(_11042_),
    .C1(_11034_),
    .D1(_11011_),
    .X(net1554));
 sky130_fd_sc_hd__buf_1 rebuffer960 (.A(_09871_),
    .X(net1555));
 sky130_fd_sc_hd__clkbuf_16 clone961 (.A(net430),
    .X(net1556));
 sky130_fd_sc_hd__buf_12 rebuffer962 (.A(net153),
    .X(net1557));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer963 (.A(net1557),
    .X(net1558));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer964 (.A(net1557),
    .X(net1559));
 sky130_fd_sc_hd__buf_12 rebuffer965 (.A(net158),
    .X(net1560));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer966 (.A(net1560),
    .X(net1561));
 sky130_fd_sc_hd__buf_16 clone969 (.A(net1565),
    .X(net1564));
 sky130_fd_sc_hd__buf_12 rebuffer970 (.A(_04661_),
    .X(net1565));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer974 (.A(net154),
    .X(net1569));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer975 (.A(net1569),
    .X(net1570));
 sky130_fd_sc_hd__buf_12 rebuffer976 (.A(net154),
    .X(net1571));
 sky130_fd_sc_hd__a31oi_4 clone980 (.A1(_02646_),
    .A2(_03478_),
    .A3(_03486_),
    .B1(_03613_),
    .Y(net1575));
 sky130_fd_sc_hd__buf_2 rebuffer984 (.A(net1578),
    .X(net1579));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer985 (.A(\id_stage_i.controller_i.instr_i[2] ),
    .X(net1580));
 sky130_fd_sc_hd__buf_12 rebuffer986 (.A(net157),
    .X(net1581));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer987 (.A(net1581),
    .X(net1582));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer988 (.A(net155),
    .X(net1583));
 sky130_fd_sc_hd__clkbuf_16 clone989 (.A(net1585),
    .X(net1584));
 sky130_fd_sc_hd__buf_12 rebuffer990 (.A(_04119_),
    .X(net1585));
 sky130_fd_sc_hd__clkbuf_16 clone991 (.A(net1565),
    .X(net1586));
 sky130_fd_sc_hd__buf_12 rebuffer992 (.A(net180),
    .X(net1587));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer993 (.A(net1587),
    .X(net1588));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer994 (.A(net1587),
    .X(net1589));
 sky130_fd_sc_hd__buf_12 rebuffer995 (.A(_09427_),
    .X(net1590));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_02113_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_02503_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_03343_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_03378_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_04865_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_04865_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_05305_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(_06990_));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(_07330_));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(_07330_));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(_08152_));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(_08547_));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(net1577));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(_09380_));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(_09524_));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(_09524_));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(_09632_));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(_09821_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(_09821_));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(_09969_));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(_10061_));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(_10061_));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(_10061_));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(_10130_));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(_10130_));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(_10130_));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(_10168_));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(_10168_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(_10168_));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(_10168_));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(_10259_));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(_10437_));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(_10437_));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(_10457_));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(_10457_));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(_10644_));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(_10644_));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(_10789_));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(_10789_));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(_10971_));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(_10974_));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(_11465_));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(_11486_));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(_11641_));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(_11641_));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(_11971_));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(_12739_));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[35] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(\gen_regfile_ff.register_file_i.waddr_a_i[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(net1273));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(net1526));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(net1530));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(net1543));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(net1552));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(net1581));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(_03738_));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(_09380_));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(_10040_));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(_10232_));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(_10232_));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(_10493_));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(_11864_));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(_11864_));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(_11971_));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(net1543));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(_10493_));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(_02301_));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(_02646_));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(_06006_));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(_08237_));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(_08269_));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(_08359_));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(_08359_));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(_08585_));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(_08658_));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(_09380_));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(_09524_));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(_09524_));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(_09606_));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(_09632_));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(_10365_));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(_10365_));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(_11273_));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(_11815_));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(_13357_));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(_13440_));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[58] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(\ex_block_i.alu_i.g_no_alu_rvb.unused_imd_val_q[58] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(net1255));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(net1259));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(net1310));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(net1534));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(net1571));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(net1571));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(net1584));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(_09283_));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_741 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_760 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_526 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_567 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_346 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_466 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_544 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_710 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_726 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_734 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_410 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_493 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_623 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_745 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_750 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_354 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_540 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_660 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_668 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_701 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_774 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_790 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_452 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_456 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_498 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_276 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_381 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_547 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_566 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_828 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_498 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_230 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_458 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_494 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_559 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_380 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_387 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_452 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_567 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_693 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_810 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_547 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_594 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_204 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_672 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_788 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_282 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_420 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_473 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_768 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_246 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_380 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_702 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_272 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_503 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_770 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_284 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_410 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_590 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_715 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_727 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_764 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_800 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_212 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_434 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_772 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_664 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_770 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_783 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_804 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_753 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_831 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_486 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_771 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_785 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_813 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_173 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_405 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_410 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_422 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_544 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_589 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_711 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_828 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_212 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_350 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_454 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_550 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_643 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_724 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_745 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_586 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_591 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_610 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_758 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_770 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_750 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_803 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_354 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_216 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_426 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_456 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_656 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_807 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_828 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_364 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_404 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_444 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_124 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_264 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_800 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_842 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_134 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_366 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_500 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_532 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_683 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_750 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_300 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_414 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_422 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_430 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_442 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_602 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_830 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_846 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_310 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_441 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_495 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_503 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_790 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_873 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_260 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_500 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_546 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_828 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_430 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_442 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_548 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_555 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_638 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_927 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_400 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_441 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_520 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_640 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_668 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_761 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_790 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_851 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_940 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_986 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_204 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_332 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_344 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_649 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_673 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_753 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_946 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_974 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_990 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_998 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1006 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_471 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_663 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_794 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_911 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_447 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_471 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_674 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_878 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_411 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_590 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_820 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_967 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1011 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_210 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_447 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_790 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_422 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_522 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_547 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_565 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_802 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_815 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_868 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1014 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1022 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1030 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_162 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_440 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_490 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_590 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_996 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1024 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1032 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1040 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1056 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1072 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_653 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_782 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_846 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_919 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_986 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1024 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1032 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_621 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_763 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_817 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_859 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_945 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1000 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1008 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_770 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_834 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_703 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_872 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_940 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1060 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1068 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_488 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_614 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_770 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_821 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_904 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_962 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1000 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1026 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1131 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1147 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_804 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_816 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_832 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_852 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_905 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_919 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1000 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1033 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1050 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1096 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1126 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_344 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_633 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_950 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_979 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_531 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_620 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_652 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_684 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_763 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_771 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_823 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_846 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_984 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_996 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1058 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1068 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1076 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1116 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1124 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1132 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_602 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1077 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_1085 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1146 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_771 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1009 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1034 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1136 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_420 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_766 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_777 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_875 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_964 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1014 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1096 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1030 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1046 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1058 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1144 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1170 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1186 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_194 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_878 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_988 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1039 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1130 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1148 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1156 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_390 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_552 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_702 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1056 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1115 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1129 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1155 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1163 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_574 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_803 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1011 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1030 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1058 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1137 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1156 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_710 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1069 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_1091 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1159 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1167 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1175 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1072 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1118 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1143 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1158 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1186 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_147 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1028 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1041 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1129 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1182 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_170 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_760 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1012 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1128 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_1166 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1186 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_564 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1002 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1050 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1054 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1071 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1098 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1120 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1159 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1176 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1184 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1002 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1010 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1026 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1048 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1086 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1132 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1161 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1175 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_518 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_704 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_958 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1028 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1056 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1175 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_646 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_650 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1027 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1035 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1074 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1096 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1131 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1173 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1200 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_170 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_556 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_986 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1053 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_170 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_979 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1023 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1035 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1054 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1083 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1099 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1146 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_477 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_976 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_986 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1088 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1120 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1129 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1137 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1161 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1177 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1185 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1200 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_958 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_980 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1012 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1078 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1107 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1138 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1147 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_411 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_974 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1010 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1073 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1128 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1159 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1184 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1200 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_974 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1012 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1033 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1053 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1116 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1125 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_982 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1094 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1119 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1131 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1161 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1200 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_636 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_652 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_964 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_984 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1002 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1182 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_653 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_724 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1108 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1131 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1140 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_700 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_963 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_980 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1028 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1036 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1044 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1060 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1076 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1160 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_650 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_727 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_964 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1080 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1159 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_652 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_676 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_684 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_770 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1023 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1034 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1132 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_776 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_988 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1035 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1072 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1113 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1133 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_968 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1028 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1048 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1072 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_960 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1006 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1014 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1131 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1146 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1189 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_523 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_644 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1023 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1096 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1104 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_1112 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_715 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_728 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_776 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_800 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1002 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1061 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1077 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1101 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1158 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1197 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_574 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_702 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_854 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1002 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1131 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1158 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_186 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_190 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_740 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_830 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_955 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1118 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1134 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1146 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1177 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_484 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_590 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1039 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1046 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1131 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_482 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_651 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_888 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_904 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_942 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1068 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1075 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1114 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1126 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1161 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1186 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_565 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_672 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_790 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_817 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_918 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_993 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1012 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1100 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1116 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1130 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1138 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1167 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_697 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_833 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_895 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1044 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1179 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_414 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_466 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_572 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_630 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_670 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_872 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_922 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_980 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1088 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1100 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1160 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_522 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_728 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_905 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_924 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_936 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_944 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_975 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1014 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1114 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1200 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_813 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_845 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_986 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1010 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1075 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1167 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_546 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_738 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_794 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_816 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_942 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_970 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1002 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1010 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1053 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1091 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1200 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_471 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_536 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_772 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_926 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1002 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1094 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1125 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_483 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_782 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_803 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_835 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1086 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1124 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1132 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_499 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_586 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_733 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_860 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_889 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_988 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1069 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1121 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1184 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_649 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_831 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_840 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1134 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1158 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1162 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1175 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_570 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_972 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1120 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1166 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_866 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_911 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1074 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1088 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1113 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1144 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1182 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_544 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_590 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_646 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_674 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1031 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1168 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_873 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1114 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1136 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1172 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1182 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_524 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_994 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1118 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1131 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1168 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1189 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1123 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1147 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_300 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_334 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_441 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_537 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_894 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1058 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1078 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1102 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1117 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1186 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_214 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_692 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_709 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1015 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1071 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1160 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1166 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_432 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_554 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_963 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1012 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1122 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1182 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_676 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1013 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1052 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1102 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1128 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1156 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1164 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1176 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_967 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_996 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1094 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1185 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_753 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_761 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_816 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_967 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_405 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_774 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_780 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1102 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1132 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1136 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1154 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1166 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_390 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_800 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1052 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1072 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1167 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_514 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_582 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_823 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_925 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_942 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_995 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1186 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_380 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_822 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_967 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1124 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1132 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1166 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_346 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_697 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_837 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_944 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1008 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1140 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1148 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1164 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_462 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_922 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_964 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_346 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_676 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_830 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_920 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_949 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_970 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_982 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1124 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1175 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_850 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_976 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_984 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_992 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_432 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_796 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_884 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_941 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_966 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1006 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1175 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_763 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_821 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_829 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_880 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_968 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1128 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1161 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1177 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1185 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_760 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_768 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_800 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_862 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_967 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_998 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1012 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1068 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1137 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1175 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_783 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_872 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1069 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1121 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1129 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1161 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1177 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1185 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_357 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_875 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_904 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1008 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1025 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1096 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1104 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1124 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1175 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1180 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1200 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_930 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1031 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1042 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1047 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1161 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1185 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_432 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1088 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1119 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1136 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_387 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_394 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_890 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1094 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1121 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1136 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1161 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1177 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1185 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_813 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1131 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_383 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_747 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_865 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_911 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1064 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1112 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_360 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1043 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1147 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_690 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_870 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1070 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1099 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_182 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_194 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_660 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_861 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_891 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_276 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_833 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1008 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1016 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1110 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1118 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1126 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1165 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_770 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_826 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_842 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1086 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_578 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_678 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_744 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_790 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_816 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_824 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_832 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_861 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1125 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_173 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_252 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_712 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_765 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_784 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_792 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_850 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_903 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_962 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1017 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1042 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1058 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1114 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1130 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1146 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_734 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_798 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_867 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1116 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1124 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1132 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1165 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1177 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1182 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_733 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_788 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_820 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_832 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_836 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1000 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1066 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1070 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_252 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_260 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_770 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_816 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_975 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1068 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1096 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_192 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_324 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_332 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_762 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_833 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_845 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_874 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_890 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1010 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1084 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1098 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1114 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_5 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_366 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_770 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_780 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_912 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_926 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1086 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1094 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_194 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_204 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_270 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_310 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_336 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_822 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_890 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_938 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_972 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1041 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1065 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_822 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1022 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1074 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_42 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_198 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_224 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_374 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_741 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_754 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_861 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_876 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_906 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_914 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1110 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1118 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1126 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_760 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_772 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_784 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_793 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_882 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_894 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1054 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1062 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1070 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1086 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1094 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_280 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_366 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_760 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_979 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1000 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1066 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_120 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_891 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_904 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_943 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_957 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1003 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1072 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_207 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_394 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_750 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_880 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_884 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_904 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_912 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_920 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_174 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_186 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_823 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_840 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_884 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_907 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_986 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1096 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_144 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_252 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_410 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_739 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_754 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_821 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_864 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_944 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1096 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1101 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1117 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1125 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_890 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_906 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_976 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1057 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1131 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1147 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_147 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_234 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_260 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_372 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_880 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_924 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1054 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1098 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_720 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_760 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_868 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_883 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1082 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1114 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1126 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1134 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1142 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1150 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1158 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1166 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_310 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_834 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1009 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1033 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1063 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1087 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_710 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_774 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_783 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1026 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1131 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1147 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_845 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_954 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1016 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1027 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1071 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1130 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_282 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_360 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_816 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_852 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_926 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_982 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1071 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1095 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1130 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_102 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_204 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_486 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_778 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_785 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_883 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_996 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1144 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1152 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1160 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1176 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1184 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_216 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_832 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_844 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_964 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1025 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1071 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1147 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_500 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_913 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_925 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1042 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1120 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_184 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_398 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_410 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_860 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_868 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_940 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_945 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1134 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1142 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1150 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1158 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1166 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_753 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1078 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1091 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1101 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1116 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_240 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_308 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_320 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_440 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_540 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_548 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_784 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_958 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1116 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1129 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1137 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_452 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_664 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_703 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_804 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_856 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_877 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_918 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1128 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1132 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_473 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_861 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_874 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_890 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_951 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1101 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1132 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1140 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1148 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1156 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_332 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_381 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_406 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_426 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_494 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_642 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_783 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_801 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_858 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_942 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_968 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_980 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1043 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_574 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_652 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_664 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_815 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1070 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1104 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_310 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_772 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_810 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_856 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_864 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_992 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1042 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1161 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1177 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1185 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_482 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_676 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_868 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_900 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_916 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_922 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_966 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_986 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_493 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_860 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_924 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_956 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1034 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1068 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_834 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_861 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_866 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_951 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1068 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1084 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1096 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1106 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_402 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_536 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_967 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_993 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1056 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1117 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1170 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1186 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_520 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_544 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_623 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_642 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_711 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_852 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_918 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_976 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1105 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1147 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_450 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_923 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1065 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_297 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_700 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_708 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_796 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_835 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_998 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1003 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1035 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1063 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1132 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1137 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_470 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_490 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_591 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_747 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_775 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_856 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_970 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_990 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_353 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_430 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_486 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_560 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_581 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_697 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_799 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_916 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_936 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_1034 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1144 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1152 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_490 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_502 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_567 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_623 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_674 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_774 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_796 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1006 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1063 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1072 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1096 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1112 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1161 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1177 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1185 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_380 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_594 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_663 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_771 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_919 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_944 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_972 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1072 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1084 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1144 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1152 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_441 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_578 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_852 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_905 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_967 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_992 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1047 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1065 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_1091 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_410 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_434 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_764 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_788 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_828 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_912 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_957 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1083 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1103 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1130 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1152 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_500 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_644 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_690 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_785 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_872 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_896 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_907 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_986 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_992 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1000 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1008 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1016 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1028 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1072 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1085 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1118 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_642 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_660 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_710 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_786 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_941 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1011 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1074 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1096 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1137 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_364 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_753 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_824 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_861 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_974 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_984 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1027 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1035 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1103 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_357 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_471 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_492 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_554 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_591 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_852 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_933 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_950 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1000 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1096 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1144 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1152 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_438 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_556 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_741 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_921 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_956 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1124 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_338 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_350 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_402 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_474 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_482 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_540 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_676 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_859 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_892 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_925 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1027 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1035 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_276 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_380 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_570 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_620 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_679 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_698 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_765 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_861 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_882 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_484 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_621 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_660 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_664 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_727 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_763 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_837 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_851 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_907 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_942 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_967 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1064 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1101 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1131 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1147 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_396 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_788 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_796 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_804 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_861 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_905 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_952 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1038 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1055 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_640 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_660 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_773 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_949 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1000 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1030 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_381 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_704 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_804 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_830 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_912 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_920 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_942 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_958 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1014 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_302 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_346 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_600 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_614 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_830 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_846 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_865 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_875 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_995 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1074 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_652 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1056 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1084 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1100 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1116 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1124 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1132 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_700 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_891 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_949 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_975 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1000 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1013 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1028 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1094 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_390 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_973 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_444 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_634 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_875 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_891 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_910 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_942 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1048 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_1054 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1065 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1073 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1201 ();
 assign alert_major_o = net470;
endmodule
