module clock_domain_crossing_fifo (rd_almost_empty,
    rd_clk,
    rd_empty,
    rd_en,
    rd_rst_n,
    wr_almost_full,
    wr_clk,
    wr_en,
    wr_full,
    wr_rst_n,
    rd_count,
    rd_data,
    wr_count,
    wr_data);
 output rd_almost_empty;
 input rd_clk;
 output rd_empty;
 input rd_en;
 input rd_rst_n;
 output wr_almost_full;
 input wr_clk;
 input wr_en;
 output wr_full;
 input wr_rst_n;
 output [4:0] rd_count;
 output [31:0] rd_data;
 output [4:0] wr_count;
 input [31:0] wr_data;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire \mem[0][0] ;
 wire \mem[0][10] ;
 wire \mem[0][11] ;
 wire \mem[0][12] ;
 wire \mem[0][13] ;
 wire \mem[0][14] ;
 wire \mem[0][15] ;
 wire \mem[0][16] ;
 wire \mem[0][17] ;
 wire \mem[0][18] ;
 wire \mem[0][19] ;
 wire \mem[0][1] ;
 wire \mem[0][20] ;
 wire \mem[0][21] ;
 wire \mem[0][22] ;
 wire \mem[0][23] ;
 wire \mem[0][24] ;
 wire \mem[0][25] ;
 wire \mem[0][26] ;
 wire \mem[0][27] ;
 wire \mem[0][28] ;
 wire \mem[0][29] ;
 wire \mem[0][2] ;
 wire \mem[0][30] ;
 wire \mem[0][31] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[0][8] ;
 wire \mem[0][9] ;
 wire \mem[10][0] ;
 wire \mem[10][10] ;
 wire \mem[10][11] ;
 wire \mem[10][12] ;
 wire \mem[10][13] ;
 wire \mem[10][14] ;
 wire \mem[10][15] ;
 wire \mem[10][16] ;
 wire \mem[10][17] ;
 wire \mem[10][18] ;
 wire \mem[10][19] ;
 wire \mem[10][1] ;
 wire \mem[10][20] ;
 wire \mem[10][21] ;
 wire \mem[10][22] ;
 wire \mem[10][23] ;
 wire \mem[10][24] ;
 wire \mem[10][25] ;
 wire \mem[10][26] ;
 wire \mem[10][27] ;
 wire \mem[10][28] ;
 wire \mem[10][29] ;
 wire \mem[10][2] ;
 wire \mem[10][30] ;
 wire \mem[10][31] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[10][8] ;
 wire \mem[10][9] ;
 wire \mem[11][0] ;
 wire \mem[11][10] ;
 wire \mem[11][11] ;
 wire \mem[11][12] ;
 wire \mem[11][13] ;
 wire \mem[11][14] ;
 wire \mem[11][15] ;
 wire \mem[11][16] ;
 wire \mem[11][17] ;
 wire \mem[11][18] ;
 wire \mem[11][19] ;
 wire \mem[11][1] ;
 wire \mem[11][20] ;
 wire \mem[11][21] ;
 wire \mem[11][22] ;
 wire \mem[11][23] ;
 wire \mem[11][24] ;
 wire \mem[11][25] ;
 wire \mem[11][26] ;
 wire \mem[11][27] ;
 wire \mem[11][28] ;
 wire \mem[11][29] ;
 wire \mem[11][2] ;
 wire \mem[11][30] ;
 wire \mem[11][31] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[11][8] ;
 wire \mem[11][9] ;
 wire \mem[12][0] ;
 wire \mem[12][10] ;
 wire \mem[12][11] ;
 wire \mem[12][12] ;
 wire \mem[12][13] ;
 wire \mem[12][14] ;
 wire \mem[12][15] ;
 wire \mem[12][16] ;
 wire \mem[12][17] ;
 wire \mem[12][18] ;
 wire \mem[12][19] ;
 wire \mem[12][1] ;
 wire \mem[12][20] ;
 wire \mem[12][21] ;
 wire \mem[12][22] ;
 wire \mem[12][23] ;
 wire \mem[12][24] ;
 wire \mem[12][25] ;
 wire \mem[12][26] ;
 wire \mem[12][27] ;
 wire \mem[12][28] ;
 wire \mem[12][29] ;
 wire \mem[12][2] ;
 wire \mem[12][30] ;
 wire \mem[12][31] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[12][8] ;
 wire \mem[12][9] ;
 wire \mem[13][0] ;
 wire \mem[13][10] ;
 wire \mem[13][11] ;
 wire \mem[13][12] ;
 wire \mem[13][13] ;
 wire \mem[13][14] ;
 wire \mem[13][15] ;
 wire \mem[13][16] ;
 wire \mem[13][17] ;
 wire \mem[13][18] ;
 wire \mem[13][19] ;
 wire \mem[13][1] ;
 wire \mem[13][20] ;
 wire \mem[13][21] ;
 wire \mem[13][22] ;
 wire \mem[13][23] ;
 wire \mem[13][24] ;
 wire \mem[13][25] ;
 wire \mem[13][26] ;
 wire \mem[13][27] ;
 wire \mem[13][28] ;
 wire \mem[13][29] ;
 wire \mem[13][2] ;
 wire \mem[13][30] ;
 wire \mem[13][31] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[13][8] ;
 wire \mem[13][9] ;
 wire \mem[14][0] ;
 wire \mem[14][10] ;
 wire \mem[14][11] ;
 wire \mem[14][12] ;
 wire \mem[14][13] ;
 wire \mem[14][14] ;
 wire \mem[14][15] ;
 wire \mem[14][16] ;
 wire \mem[14][17] ;
 wire \mem[14][18] ;
 wire \mem[14][19] ;
 wire \mem[14][1] ;
 wire \mem[14][20] ;
 wire \mem[14][21] ;
 wire \mem[14][22] ;
 wire \mem[14][23] ;
 wire \mem[14][24] ;
 wire \mem[14][25] ;
 wire \mem[14][26] ;
 wire \mem[14][27] ;
 wire \mem[14][28] ;
 wire \mem[14][29] ;
 wire \mem[14][2] ;
 wire \mem[14][30] ;
 wire \mem[14][31] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[14][8] ;
 wire \mem[14][9] ;
 wire \mem[15][0] ;
 wire \mem[15][10] ;
 wire \mem[15][11] ;
 wire \mem[15][12] ;
 wire \mem[15][13] ;
 wire \mem[15][14] ;
 wire \mem[15][15] ;
 wire \mem[15][16] ;
 wire \mem[15][17] ;
 wire \mem[15][18] ;
 wire \mem[15][19] ;
 wire \mem[15][1] ;
 wire \mem[15][20] ;
 wire \mem[15][21] ;
 wire \mem[15][22] ;
 wire \mem[15][23] ;
 wire \mem[15][24] ;
 wire \mem[15][25] ;
 wire \mem[15][26] ;
 wire \mem[15][27] ;
 wire \mem[15][28] ;
 wire \mem[15][29] ;
 wire \mem[15][2] ;
 wire \mem[15][30] ;
 wire \mem[15][31] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[15][8] ;
 wire \mem[15][9] ;
 wire \mem[1][0] ;
 wire \mem[1][10] ;
 wire \mem[1][11] ;
 wire \mem[1][12] ;
 wire \mem[1][13] ;
 wire \mem[1][14] ;
 wire \mem[1][15] ;
 wire \mem[1][16] ;
 wire \mem[1][17] ;
 wire \mem[1][18] ;
 wire \mem[1][19] ;
 wire \mem[1][1] ;
 wire \mem[1][20] ;
 wire \mem[1][21] ;
 wire \mem[1][22] ;
 wire \mem[1][23] ;
 wire \mem[1][24] ;
 wire \mem[1][25] ;
 wire \mem[1][26] ;
 wire \mem[1][27] ;
 wire \mem[1][28] ;
 wire \mem[1][29] ;
 wire \mem[1][2] ;
 wire \mem[1][30] ;
 wire \mem[1][31] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[1][8] ;
 wire \mem[1][9] ;
 wire \mem[2][0] ;
 wire \mem[2][10] ;
 wire \mem[2][11] ;
 wire \mem[2][12] ;
 wire \mem[2][13] ;
 wire \mem[2][14] ;
 wire \mem[2][15] ;
 wire \mem[2][16] ;
 wire \mem[2][17] ;
 wire \mem[2][18] ;
 wire \mem[2][19] ;
 wire \mem[2][1] ;
 wire \mem[2][20] ;
 wire \mem[2][21] ;
 wire \mem[2][22] ;
 wire \mem[2][23] ;
 wire \mem[2][24] ;
 wire \mem[2][25] ;
 wire \mem[2][26] ;
 wire \mem[2][27] ;
 wire \mem[2][28] ;
 wire \mem[2][29] ;
 wire \mem[2][2] ;
 wire \mem[2][30] ;
 wire \mem[2][31] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[2][8] ;
 wire \mem[2][9] ;
 wire \mem[3][0] ;
 wire \mem[3][10] ;
 wire \mem[3][11] ;
 wire \mem[3][12] ;
 wire \mem[3][13] ;
 wire \mem[3][14] ;
 wire \mem[3][15] ;
 wire \mem[3][16] ;
 wire \mem[3][17] ;
 wire \mem[3][18] ;
 wire \mem[3][19] ;
 wire \mem[3][1] ;
 wire \mem[3][20] ;
 wire \mem[3][21] ;
 wire \mem[3][22] ;
 wire \mem[3][23] ;
 wire \mem[3][24] ;
 wire \mem[3][25] ;
 wire \mem[3][26] ;
 wire \mem[3][27] ;
 wire \mem[3][28] ;
 wire \mem[3][29] ;
 wire \mem[3][2] ;
 wire \mem[3][30] ;
 wire \mem[3][31] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[3][8] ;
 wire \mem[3][9] ;
 wire \mem[4][0] ;
 wire \mem[4][10] ;
 wire \mem[4][11] ;
 wire \mem[4][12] ;
 wire \mem[4][13] ;
 wire \mem[4][14] ;
 wire \mem[4][15] ;
 wire \mem[4][16] ;
 wire \mem[4][17] ;
 wire \mem[4][18] ;
 wire \mem[4][19] ;
 wire \mem[4][1] ;
 wire \mem[4][20] ;
 wire \mem[4][21] ;
 wire \mem[4][22] ;
 wire \mem[4][23] ;
 wire \mem[4][24] ;
 wire \mem[4][25] ;
 wire \mem[4][26] ;
 wire \mem[4][27] ;
 wire \mem[4][28] ;
 wire \mem[4][29] ;
 wire \mem[4][2] ;
 wire \mem[4][30] ;
 wire \mem[4][31] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[4][8] ;
 wire \mem[4][9] ;
 wire \mem[5][0] ;
 wire \mem[5][10] ;
 wire \mem[5][11] ;
 wire \mem[5][12] ;
 wire \mem[5][13] ;
 wire \mem[5][14] ;
 wire \mem[5][15] ;
 wire \mem[5][16] ;
 wire \mem[5][17] ;
 wire \mem[5][18] ;
 wire \mem[5][19] ;
 wire \mem[5][1] ;
 wire \mem[5][20] ;
 wire \mem[5][21] ;
 wire \mem[5][22] ;
 wire \mem[5][23] ;
 wire \mem[5][24] ;
 wire \mem[5][25] ;
 wire \mem[5][26] ;
 wire \mem[5][27] ;
 wire \mem[5][28] ;
 wire \mem[5][29] ;
 wire \mem[5][2] ;
 wire \mem[5][30] ;
 wire \mem[5][31] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[5][8] ;
 wire \mem[5][9] ;
 wire \mem[6][0] ;
 wire \mem[6][10] ;
 wire \mem[6][11] ;
 wire \mem[6][12] ;
 wire \mem[6][13] ;
 wire \mem[6][14] ;
 wire \mem[6][15] ;
 wire \mem[6][16] ;
 wire \mem[6][17] ;
 wire \mem[6][18] ;
 wire \mem[6][19] ;
 wire \mem[6][1] ;
 wire \mem[6][20] ;
 wire \mem[6][21] ;
 wire \mem[6][22] ;
 wire \mem[6][23] ;
 wire \mem[6][24] ;
 wire \mem[6][25] ;
 wire \mem[6][26] ;
 wire \mem[6][27] ;
 wire \mem[6][28] ;
 wire \mem[6][29] ;
 wire \mem[6][2] ;
 wire \mem[6][30] ;
 wire \mem[6][31] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[6][8] ;
 wire \mem[6][9] ;
 wire \mem[7][0] ;
 wire \mem[7][10] ;
 wire \mem[7][11] ;
 wire \mem[7][12] ;
 wire \mem[7][13] ;
 wire \mem[7][14] ;
 wire \mem[7][15] ;
 wire \mem[7][16] ;
 wire \mem[7][17] ;
 wire \mem[7][18] ;
 wire \mem[7][19] ;
 wire \mem[7][1] ;
 wire \mem[7][20] ;
 wire \mem[7][21] ;
 wire \mem[7][22] ;
 wire \mem[7][23] ;
 wire \mem[7][24] ;
 wire \mem[7][25] ;
 wire \mem[7][26] ;
 wire \mem[7][27] ;
 wire \mem[7][28] ;
 wire \mem[7][29] ;
 wire \mem[7][2] ;
 wire \mem[7][30] ;
 wire \mem[7][31] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[7][8] ;
 wire \mem[7][9] ;
 wire \mem[8][0] ;
 wire \mem[8][10] ;
 wire \mem[8][11] ;
 wire \mem[8][12] ;
 wire \mem[8][13] ;
 wire \mem[8][14] ;
 wire \mem[8][15] ;
 wire \mem[8][16] ;
 wire \mem[8][17] ;
 wire \mem[8][18] ;
 wire \mem[8][19] ;
 wire \mem[8][1] ;
 wire \mem[8][20] ;
 wire \mem[8][21] ;
 wire \mem[8][22] ;
 wire \mem[8][23] ;
 wire \mem[8][24] ;
 wire \mem[8][25] ;
 wire \mem[8][26] ;
 wire \mem[8][27] ;
 wire \mem[8][28] ;
 wire \mem[8][29] ;
 wire \mem[8][2] ;
 wire \mem[8][30] ;
 wire \mem[8][31] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[8][8] ;
 wire \mem[8][9] ;
 wire \mem[9][0] ;
 wire \mem[9][10] ;
 wire \mem[9][11] ;
 wire \mem[9][12] ;
 wire \mem[9][13] ;
 wire \mem[9][14] ;
 wire \mem[9][15] ;
 wire \mem[9][16] ;
 wire \mem[9][17] ;
 wire \mem[9][18] ;
 wire \mem[9][19] ;
 wire \mem[9][1] ;
 wire \mem[9][20] ;
 wire \mem[9][21] ;
 wire \mem[9][22] ;
 wire \mem[9][23] ;
 wire \mem[9][24] ;
 wire \mem[9][25] ;
 wire \mem[9][26] ;
 wire \mem[9][27] ;
 wire \mem[9][28] ;
 wire \mem[9][29] ;
 wire \mem[9][2] ;
 wire \mem[9][30] ;
 wire \mem[9][31] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \mem[9][8] ;
 wire \mem[9][9] ;
 wire \rd_ptr_bin[0] ;
 wire \rd_ptr_bin[1] ;
 wire \rd_ptr_bin[2] ;
 wire \rd_ptr_bin[3] ;
 wire \rd_ptr_bin[4] ;
 wire \rd_ptr_gray[0] ;
 wire \rd_ptr_gray[1] ;
 wire \rd_ptr_gray[2] ;
 wire \rd_ptr_gray[3] ;
 wire \rd_ptr_gray_sync1[0] ;
 wire \rd_ptr_gray_sync1[1] ;
 wire \rd_ptr_gray_sync1[2] ;
 wire \rd_ptr_gray_sync1[3] ;
 wire \rd_ptr_gray_sync1[4] ;
 wire \rd_ptr_gray_sync2[0] ;
 wire \rd_ptr_gray_sync2[1] ;
 wire \rd_ptr_gray_sync2[2] ;
 wire \rd_ptr_gray_sync2[3] ;
 wire \rd_ptr_gray_sync2[4] ;
 wire \wr_ptr_bin[0] ;
 wire \wr_ptr_bin[1] ;
 wire \wr_ptr_bin[2] ;
 wire \wr_ptr_bin[3] ;
 wire \wr_ptr_bin[4] ;
 wire \wr_ptr_gray[0] ;
 wire \wr_ptr_gray[1] ;
 wire \wr_ptr_gray[2] ;
 wire \wr_ptr_gray[3] ;
 wire \wr_ptr_gray_sync1[0] ;
 wire \wr_ptr_gray_sync1[1] ;
 wire \wr_ptr_gray_sync1[2] ;
 wire \wr_ptr_gray_sync1[3] ;
 wire \wr_ptr_gray_sync1[4] ;
 wire \wr_ptr_gray_sync2[0] ;
 wire \wr_ptr_gray_sync2[1] ;
 wire \wr_ptr_gray_sync2[2] ;
 wire \wr_ptr_gray_sync2[3] ;
 wire \wr_ptr_gray_sync2[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire clknet_leaf_0_wr_clk;
 wire clknet_leaf_1_wr_clk;
 wire clknet_leaf_2_wr_clk;
 wire clknet_leaf_3_wr_clk;
 wire clknet_leaf_4_wr_clk;
 wire clknet_leaf_5_wr_clk;
 wire clknet_leaf_6_wr_clk;
 wire clknet_leaf_7_wr_clk;
 wire clknet_leaf_8_wr_clk;
 wire clknet_leaf_9_wr_clk;
 wire clknet_leaf_10_wr_clk;
 wire clknet_leaf_11_wr_clk;
 wire clknet_leaf_12_wr_clk;
 wire clknet_leaf_13_wr_clk;
 wire clknet_leaf_14_wr_clk;
 wire clknet_leaf_15_wr_clk;
 wire clknet_leaf_16_wr_clk;
 wire clknet_leaf_17_wr_clk;
 wire clknet_leaf_18_wr_clk;
 wire clknet_leaf_19_wr_clk;
 wire clknet_0_wr_clk;
 wire clknet_1_0__leaf_wr_clk;
 wire clknet_1_1__leaf_wr_clk;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;

 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1525_ (.A1(\rd_ptr_gray_sync2[3] ),
    .A2(\rd_ptr_gray_sync2[4] ),
    .ZN(_1492_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1526_ (.A1(\rd_ptr_gray_sync2[2] ),
    .A2(_1492_),
    .Z(_1489_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1527_ (.A1(\rd_ptr_gray_sync2[1] ),
    .A2(_1489_),
    .Z(_1482_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1528_ (.I(_1524_),
    .ZN(net79));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1529_ (.A1(\rd_ptr_gray_sync2[4] ),
    .A2(\wr_ptr_bin[4] ),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _1530_ (.A1(_1494_),
    .A2(_1491_),
    .A3(_1488_),
    .A4(_1524_),
    .Z(_0567_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _1531_ (.A1(_0566_),
    .A2(_0567_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1532_ (.I(_0568_),
    .ZN(net84));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1533_ (.I(_1478_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1534_ (.A1(_0569_),
    .A2(_1488_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1535_ (.A1(_1487_),
    .A2(_0570_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1536_ (.A1(_1491_),
    .A2(_0571_),
    .B(_1490_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1537_ (.A1(_1494_),
    .A2(_0572_),
    .Z(_0573_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1538_ (.I(_0573_),
    .ZN(net82));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1539_ (.I(_1480_),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1540_ (.A1(_0574_),
    .A2(_1491_),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1541_ (.A1(_1490_),
    .A2(_0575_),
    .Z(_0576_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1542_ (.A1(_1494_),
    .A2(_0576_),
    .B(_1493_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1543_ (.A1(_0566_),
    .A2(_0577_),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1544_ (.I(_0578_),
    .ZN(net83));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1545_ (.A1(\wr_ptr_gray_sync2[3] ),
    .A2(\wr_ptr_gray_sync2[4] ),
    .Z(_1500_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1546_ (.A1(\wr_ptr_gray_sync2[2] ),
    .A2(_1500_),
    .Z(_1504_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1547_ (.A1(\wr_ptr_gray_sync2[1] ),
    .A2(_1504_),
    .ZN(_1484_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1548_ (.I(_1486_),
    .ZN(net41));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1549_ (.A1(_1485_),
    .A2(_1506_),
    .ZN(net42));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1550_ (.I(_1483_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1551_ (.A1(_1498_),
    .A2(_0579_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1552_ (.A1(_1497_),
    .A2(_0580_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1553_ (.A1(_1506_),
    .A2(_0581_),
    .B(_1505_),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1554_ (.A1(_1502_),
    .A2(_0582_),
    .ZN(net43));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1555_ (.A1(\wr_ptr_gray_sync2[4] ),
    .A2(\rd_ptr_bin[4] ),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1556_ (.I(_1485_),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1557_ (.A1(_0584_),
    .A2(_1506_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1558_ (.A1(_1505_),
    .A2(_0585_),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _1559_ (.A1(_1502_),
    .A2(_0586_),
    .B(_1501_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1560_ (.A1(_0583_),
    .A2(_0587_),
    .Z(net44));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1561_ (.A1(\wr_ptr_gray_sync2[3] ),
    .A2(\rd_ptr_gray[3] ),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1562_ (.A1(\wr_ptr_gray_sync2[0] ),
    .A2(\rd_ptr_gray[0] ),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _1563_ (.A1(_0588_),
    .A2(_0589_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1564_ (.A1(\wr_ptr_gray_sync2[1] ),
    .A2(\rd_ptr_gray[1] ),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1565_ (.A1(\wr_ptr_gray_sync2[2] ),
    .A2(\rd_ptr_gray[2] ),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _1566_ (.A1(_0583_),
    .A2(_0590_),
    .A3(_0591_),
    .A4(_0592_),
    .Z(_0593_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1567_ (.I(_0593_),
    .ZN(net77));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _1568_ (.I(\rd_ptr_bin[2] ),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _1569_ (.I(_0594_),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1570_ (.I(_0595_),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _1571_ (.I(_0596_),
    .Z(_1503_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _1572_ (.I(\rd_ptr_bin[3] ),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1573_ (.I(_0597_),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1574_ (.I(_0598_),
    .Z(_1499_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1575_ (.I(_1482_),
    .ZN(_1479_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1576_ (.I(\wr_ptr_bin[0] ),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1577_ (.I(\rd_ptr_bin[0] ),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1578_ (.I(_1484_),
    .ZN(_1496_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1579_ (.I(\wr_ptr_bin[1] ),
    .ZN(_1477_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _1580_ (.I(\rd_ptr_bin[1] ),
    .ZN(_1495_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _1581_ (.A1(\wr_ptr_gray_sync2[0] ),
    .A2(_1484_),
    .Z(_1521_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _1582_ (.A1(\rd_ptr_gray_sync2[0] ),
    .A2(_1482_),
    .ZN(_1523_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1583_ (.I(_1522_),
    .ZN(net40));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _1584_ (.I(net5),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1585_ (.I(\wr_ptr_bin[2] ),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _1586_ (.I(\wr_ptr_bin[3] ),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1587_ (.A1(_0600_),
    .A2(_0601_),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1588_ (.A1(net37),
    .A2(net38),
    .A3(_1507_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1589_ (.A1(_0568_),
    .A2(_0603_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _1590_ (.A1(_0602_),
    .A2(_0604_),
    .Z(_0605_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _1591_ (.I(_0605_),
    .Z(_0606_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1592_ (.I0(\mem[0][0] ),
    .I1(_0599_),
    .S(_0606_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _1593_ (.I(net6),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1594_ (.I0(\mem[0][10] ),
    .I1(_0607_),
    .S(_0606_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _1595_ (.I(net7),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1596_ (.I0(\mem[0][11] ),
    .I1(_0608_),
    .S(_0606_),
    .Z(_0006_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _1597_ (.I(net8),
    .Z(_0609_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1598_ (.I0(\mem[0][12] ),
    .I1(_0609_),
    .S(_0606_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _1599_ (.I(net9),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1600_ (.I0(\mem[0][13] ),
    .I1(_0610_),
    .S(_0606_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _1601_ (.I(net10),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1602_ (.I0(\mem[0][14] ),
    .I1(_0611_),
    .S(_0606_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _1603_ (.I(net11),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1604_ (.I0(\mem[0][15] ),
    .I1(_0612_),
    .S(_0606_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _1605_ (.I(net12),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1606_ (.I0(\mem[0][16] ),
    .I1(_0613_),
    .S(_0606_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _1607_ (.I(net13),
    .Z(_0614_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1608_ (.I0(\mem[0][17] ),
    .I1(_0614_),
    .S(_0606_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _1609_ (.I(net14),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1610_ (.I0(\mem[0][18] ),
    .I1(_0615_),
    .S(_0606_),
    .Z(_0013_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _1611_ (.I(net15),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _1612_ (.I(_0605_),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1613_ (.I0(\mem[0][19] ),
    .I1(_0616_),
    .S(_0617_),
    .Z(_0014_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _1614_ (.I(net16),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1615_ (.I0(\mem[0][1] ),
    .I1(_0618_),
    .S(_0617_),
    .Z(_0015_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _1616_ (.I(net17),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1617_ (.I0(\mem[0][20] ),
    .I1(_0619_),
    .S(_0617_),
    .Z(_0016_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _1618_ (.I(net18),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1619_ (.I0(\mem[0][21] ),
    .I1(_0620_),
    .S(_0617_),
    .Z(_0017_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _1620_ (.I(net19),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1621_ (.I0(\mem[0][22] ),
    .I1(_0621_),
    .S(_0617_),
    .Z(_0018_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _1622_ (.I(net20),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1623_ (.I0(\mem[0][23] ),
    .I1(_0622_),
    .S(_0617_),
    .Z(_0019_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _1624_ (.I(net21),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1625_ (.I0(\mem[0][24] ),
    .I1(_0623_),
    .S(_0617_),
    .Z(_0020_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _1626_ (.I(net22),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1627_ (.I0(\mem[0][25] ),
    .I1(_0624_),
    .S(_0617_),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _1628_ (.I(net23),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1629_ (.I0(\mem[0][26] ),
    .I1(_0625_),
    .S(_0617_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _1630_ (.I(net24),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1631_ (.I0(\mem[0][27] ),
    .I1(_0626_),
    .S(_0617_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 _1632_ (.I(net25),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1633_ (.I(_0605_),
    .Z(_0628_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1634_ (.I0(\mem[0][28] ),
    .I1(_0627_),
    .S(_0628_),
    .Z(_0024_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _1635_ (.I(net26),
    .Z(_0629_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1636_ (.I0(\mem[0][29] ),
    .I1(_0629_),
    .S(_0628_),
    .Z(_0025_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _1637_ (.I(net27),
    .Z(_0630_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1638_ (.I0(\mem[0][2] ),
    .I1(_0630_),
    .S(_0628_),
    .Z(_0026_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _1639_ (.I(net28),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1640_ (.I0(\mem[0][30] ),
    .I1(_0631_),
    .S(_0628_),
    .Z(_0027_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _1641_ (.I(net29),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1642_ (.I0(\mem[0][31] ),
    .I1(_0632_),
    .S(_0628_),
    .Z(_0028_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 _1643_ (.I(net30),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1644_ (.I0(\mem[0][3] ),
    .I1(_0633_),
    .S(_0628_),
    .Z(_0029_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _1645_ (.I(net31),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1646_ (.I0(\mem[0][4] ),
    .I1(_0634_),
    .S(_0628_),
    .Z(_0030_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _1647_ (.I(net32),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1648_ (.I0(\mem[0][5] ),
    .I1(_0635_),
    .S(_0628_),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _1649_ (.I(net33),
    .Z(_0636_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1650_ (.I0(\mem[0][6] ),
    .I1(_0636_),
    .S(_0628_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _1651_ (.I(net34),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1652_ (.I0(\mem[0][7] ),
    .I1(_0637_),
    .S(_0628_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _1653_ (.I(net35),
    .Z(_0638_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1654_ (.I0(\mem[0][8] ),
    .I1(_0638_),
    .S(_0605_),
    .Z(_0034_));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 _1655_ (.I(net36),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1656_ (.I0(\mem[0][9] ),
    .I1(_0639_),
    .S(_0605_),
    .Z(_0035_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1657_ (.A1(net37),
    .A2(net38),
    .A3(_1508_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1658_ (.A1(_0600_),
    .A2(\wr_ptr_bin[3] ),
    .A3(_0568_),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _1659_ (.A1(_0640_),
    .A2(_0641_),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1660_ (.I(_0642_),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1661_ (.I0(\mem[10][0] ),
    .I1(_0599_),
    .S(_0643_),
    .Z(_0036_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1662_ (.I0(\mem[10][10] ),
    .I1(_0607_),
    .S(_0643_),
    .Z(_0037_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1663_ (.I0(\mem[10][11] ),
    .I1(_0608_),
    .S(_0643_),
    .Z(_0038_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1664_ (.I0(\mem[10][12] ),
    .I1(_0609_),
    .S(_0643_),
    .Z(_0039_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1665_ (.I0(\mem[10][13] ),
    .I1(_0610_),
    .S(_0643_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1666_ (.I0(\mem[10][14] ),
    .I1(_0611_),
    .S(_0643_),
    .Z(_0041_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1667_ (.I0(\mem[10][15] ),
    .I1(_0612_),
    .S(_0643_),
    .Z(_0042_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1668_ (.I0(\mem[10][16] ),
    .I1(_0613_),
    .S(_0643_),
    .Z(_0043_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1669_ (.I0(\mem[10][17] ),
    .I1(_0614_),
    .S(_0643_),
    .Z(_0044_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1670_ (.I0(\mem[10][18] ),
    .I1(_0615_),
    .S(_0643_),
    .Z(_0045_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _1671_ (.I(_0642_),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1672_ (.I0(\mem[10][19] ),
    .I1(_0616_),
    .S(_0644_),
    .Z(_0046_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1673_ (.I0(\mem[10][1] ),
    .I1(_0618_),
    .S(_0644_),
    .Z(_0047_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1674_ (.I0(\mem[10][20] ),
    .I1(_0619_),
    .S(_0644_),
    .Z(_0048_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1675_ (.I0(\mem[10][21] ),
    .I1(_0620_),
    .S(_0644_),
    .Z(_0049_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1676_ (.I0(\mem[10][22] ),
    .I1(_0621_),
    .S(_0644_),
    .Z(_0050_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1677_ (.I0(\mem[10][23] ),
    .I1(_0622_),
    .S(_0644_),
    .Z(_0051_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1678_ (.I0(\mem[10][24] ),
    .I1(_0623_),
    .S(_0644_),
    .Z(_0052_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1679_ (.I0(\mem[10][25] ),
    .I1(_0624_),
    .S(_0644_),
    .Z(_0053_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1680_ (.I0(\mem[10][26] ),
    .I1(_0625_),
    .S(_0644_),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1681_ (.I0(\mem[10][27] ),
    .I1(_0626_),
    .S(_0644_),
    .Z(_0055_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _1682_ (.I(_0642_),
    .Z(_0645_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1683_ (.I0(\mem[10][28] ),
    .I1(_0627_),
    .S(_0645_),
    .Z(_0056_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1684_ (.I0(\mem[10][29] ),
    .I1(_0629_),
    .S(_0645_),
    .Z(_0057_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1685_ (.I0(\mem[10][2] ),
    .I1(_0630_),
    .S(_0645_),
    .Z(_0058_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1686_ (.I0(\mem[10][30] ),
    .I1(_0631_),
    .S(_0645_),
    .Z(_0059_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1687_ (.I0(\mem[10][31] ),
    .I1(_0632_),
    .S(_0645_),
    .Z(_0060_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1688_ (.I0(\mem[10][3] ),
    .I1(_0633_),
    .S(_0645_),
    .Z(_0061_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1689_ (.I0(\mem[10][4] ),
    .I1(_0634_),
    .S(_0645_),
    .Z(_0062_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1690_ (.I0(\mem[10][5] ),
    .I1(_0635_),
    .S(_0645_),
    .Z(_0063_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1691_ (.I0(\mem[10][6] ),
    .I1(_0636_),
    .S(_0645_),
    .Z(_0064_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1692_ (.I0(\mem[10][7] ),
    .I1(_0637_),
    .S(_0645_),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1693_ (.I0(\mem[10][8] ),
    .I1(_0638_),
    .S(_0642_),
    .Z(_0066_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1694_ (.I0(\mem[10][9] ),
    .I1(_0639_),
    .S(_0642_),
    .Z(_0067_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1695_ (.A1(net37),
    .A2(net38),
    .A3(_1512_),
    .Z(_0646_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _1696_ (.A1(_0641_),
    .A2(_0646_),
    .Z(_0647_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1697_ (.I(_0647_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1698_ (.I0(\mem[11][0] ),
    .I1(_0599_),
    .S(_0648_),
    .Z(_0068_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1699_ (.I0(\mem[11][10] ),
    .I1(_0607_),
    .S(_0648_),
    .Z(_0069_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1700_ (.I0(\mem[11][11] ),
    .I1(_0608_),
    .S(_0648_),
    .Z(_0070_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1701_ (.I0(\mem[11][12] ),
    .I1(_0609_),
    .S(_0648_),
    .Z(_0071_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1702_ (.I0(\mem[11][13] ),
    .I1(_0610_),
    .S(_0648_),
    .Z(_0072_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1703_ (.I0(\mem[11][14] ),
    .I1(_0611_),
    .S(_0648_),
    .Z(_0073_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1704_ (.I0(\mem[11][15] ),
    .I1(_0612_),
    .S(_0648_),
    .Z(_0074_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1705_ (.I0(\mem[11][16] ),
    .I1(_0613_),
    .S(_0648_),
    .Z(_0075_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1706_ (.I0(\mem[11][17] ),
    .I1(_0614_),
    .S(_0648_),
    .Z(_0076_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1707_ (.I0(\mem[11][18] ),
    .I1(_0615_),
    .S(_0648_),
    .Z(_0077_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1708_ (.I(_0647_),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1709_ (.I0(\mem[11][19] ),
    .I1(_0616_),
    .S(_0649_),
    .Z(_0078_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1710_ (.I0(\mem[11][1] ),
    .I1(_0618_),
    .S(_0649_),
    .Z(_0079_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1711_ (.I0(\mem[11][20] ),
    .I1(_0619_),
    .S(_0649_),
    .Z(_0080_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1712_ (.I0(\mem[11][21] ),
    .I1(_0620_),
    .S(_0649_),
    .Z(_0081_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1713_ (.I0(\mem[11][22] ),
    .I1(_0621_),
    .S(_0649_),
    .Z(_0082_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1714_ (.I0(\mem[11][23] ),
    .I1(_0622_),
    .S(_0649_),
    .Z(_0083_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1715_ (.I0(\mem[11][24] ),
    .I1(_0623_),
    .S(_0649_),
    .Z(_0084_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1716_ (.I0(\mem[11][25] ),
    .I1(_0624_),
    .S(_0649_),
    .Z(_0085_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1717_ (.I0(\mem[11][26] ),
    .I1(_0625_),
    .S(_0649_),
    .Z(_0086_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1718_ (.I0(\mem[11][27] ),
    .I1(_0626_),
    .S(_0649_),
    .Z(_0087_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1719_ (.I(_0647_),
    .Z(_0650_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1720_ (.I0(\mem[11][28] ),
    .I1(_0627_),
    .S(_0650_),
    .Z(_0088_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1721_ (.I0(\mem[11][29] ),
    .I1(_0629_),
    .S(_0650_),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1722_ (.I0(\mem[11][2] ),
    .I1(_0630_),
    .S(_0650_),
    .Z(_0090_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1723_ (.I0(\mem[11][30] ),
    .I1(_0631_),
    .S(_0650_),
    .Z(_0091_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1724_ (.I0(\mem[11][31] ),
    .I1(_0632_),
    .S(_0650_),
    .Z(_0092_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1725_ (.I0(\mem[11][3] ),
    .I1(_0633_),
    .S(_0650_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1726_ (.I0(\mem[11][4] ),
    .I1(_0634_),
    .S(_0650_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1727_ (.I0(\mem[11][5] ),
    .I1(_0635_),
    .S(_0650_),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1728_ (.I0(\mem[11][6] ),
    .I1(_0636_),
    .S(_0650_),
    .Z(_0096_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1729_ (.I0(\mem[11][7] ),
    .I1(_0637_),
    .S(_0650_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1730_ (.I0(\mem[11][8] ),
    .I1(_0638_),
    .S(_0647_),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1731_ (.I0(\mem[11][9] ),
    .I1(_0639_),
    .S(_0647_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1732_ (.A1(\wr_ptr_bin[2] ),
    .A2(\wr_ptr_bin[3] ),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _1733_ (.A1(_0604_),
    .A2(_0651_),
    .Z(_0652_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _1734_ (.I(_0652_),
    .Z(_0653_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1735_ (.I0(\mem[12][0] ),
    .I1(_0599_),
    .S(_0653_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1736_ (.I0(\mem[12][10] ),
    .I1(_0607_),
    .S(_0653_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1737_ (.I0(\mem[12][11] ),
    .I1(_0608_),
    .S(_0653_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1738_ (.I0(\mem[12][12] ),
    .I1(_0609_),
    .S(_0653_),
    .Z(_0103_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1739_ (.I0(\mem[12][13] ),
    .I1(_0610_),
    .S(_0653_),
    .Z(_0104_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1740_ (.I0(\mem[12][14] ),
    .I1(_0611_),
    .S(_0653_),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1741_ (.I0(\mem[12][15] ),
    .I1(_0612_),
    .S(_0653_),
    .Z(_0106_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1742_ (.I0(\mem[12][16] ),
    .I1(_0613_),
    .S(_0653_),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1743_ (.I0(\mem[12][17] ),
    .I1(_0614_),
    .S(_0653_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1744_ (.I0(\mem[12][18] ),
    .I1(_0615_),
    .S(_0653_),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _1745_ (.I(_0652_),
    .Z(_0654_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1746_ (.I0(\mem[12][19] ),
    .I1(_0616_),
    .S(_0654_),
    .Z(_0110_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1747_ (.I0(\mem[12][1] ),
    .I1(_0618_),
    .S(_0654_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1748_ (.I0(\mem[12][20] ),
    .I1(_0619_),
    .S(_0654_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1749_ (.I0(\mem[12][21] ),
    .I1(_0620_),
    .S(_0654_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1750_ (.I0(\mem[12][22] ),
    .I1(_0621_),
    .S(_0654_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1751_ (.I0(\mem[12][23] ),
    .I1(_0622_),
    .S(_0654_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1752_ (.I0(\mem[12][24] ),
    .I1(_0623_),
    .S(_0654_),
    .Z(_0116_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1753_ (.I0(\mem[12][25] ),
    .I1(_0624_),
    .S(_0654_),
    .Z(_0117_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1754_ (.I0(\mem[12][26] ),
    .I1(_0625_),
    .S(_0654_),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1755_ (.I0(\mem[12][27] ),
    .I1(_0626_),
    .S(_0654_),
    .Z(_0119_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1756_ (.I(_0652_),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1757_ (.I0(\mem[12][28] ),
    .I1(_0627_),
    .S(_0655_),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1758_ (.I0(\mem[12][29] ),
    .I1(_0629_),
    .S(_0655_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1759_ (.I0(\mem[12][2] ),
    .I1(_0630_),
    .S(_0655_),
    .Z(_0122_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1760_ (.I0(\mem[12][30] ),
    .I1(_0631_),
    .S(_0655_),
    .Z(_0123_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1761_ (.I0(\mem[12][31] ),
    .I1(_0632_),
    .S(_0655_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1762_ (.I0(\mem[12][3] ),
    .I1(_0633_),
    .S(_0655_),
    .Z(_0125_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1763_ (.I0(\mem[12][4] ),
    .I1(_0634_),
    .S(_0655_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1764_ (.I0(\mem[12][5] ),
    .I1(_0635_),
    .S(_0655_),
    .Z(_0127_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1765_ (.I0(\mem[12][6] ),
    .I1(_0636_),
    .S(_0655_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1766_ (.I0(\mem[12][7] ),
    .I1(_0637_),
    .S(_0655_),
    .Z(_0129_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1767_ (.I0(\mem[12][8] ),
    .I1(_0638_),
    .S(_0652_),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1768_ (.I0(\mem[12][9] ),
    .I1(_0639_),
    .S(_0652_),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1769_ (.A1(net37),
    .A2(net38),
    .A3(_1510_),
    .Z(_0656_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1770_ (.A1(_0568_),
    .A2(_0656_),
    .Z(_0657_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _1771_ (.A1(_0651_),
    .A2(_0657_),
    .Z(_0658_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _1772_ (.I(_0658_),
    .Z(_0659_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1773_ (.I0(\mem[13][0] ),
    .I1(_0599_),
    .S(_0659_),
    .Z(_0132_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1774_ (.I0(\mem[13][10] ),
    .I1(_0607_),
    .S(_0659_),
    .Z(_0133_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1775_ (.I0(\mem[13][11] ),
    .I1(_0608_),
    .S(_0659_),
    .Z(_0134_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1776_ (.I0(\mem[13][12] ),
    .I1(_0609_),
    .S(_0659_),
    .Z(_0135_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1777_ (.I0(\mem[13][13] ),
    .I1(_0610_),
    .S(_0659_),
    .Z(_0136_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1778_ (.I0(\mem[13][14] ),
    .I1(_0611_),
    .S(_0659_),
    .Z(_0137_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1779_ (.I0(\mem[13][15] ),
    .I1(_0612_),
    .S(_0659_),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1780_ (.I0(\mem[13][16] ),
    .I1(_0613_),
    .S(_0659_),
    .Z(_0139_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1781_ (.I0(\mem[13][17] ),
    .I1(_0614_),
    .S(_0659_),
    .Z(_0140_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1782_ (.I0(\mem[13][18] ),
    .I1(_0615_),
    .S(_0659_),
    .Z(_0141_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _1783_ (.I(_0658_),
    .Z(_0660_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1784_ (.I0(\mem[13][19] ),
    .I1(_0616_),
    .S(_0660_),
    .Z(_0142_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1785_ (.I0(\mem[13][1] ),
    .I1(_0618_),
    .S(_0660_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1786_ (.I0(\mem[13][20] ),
    .I1(_0619_),
    .S(_0660_),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1787_ (.I0(\mem[13][21] ),
    .I1(_0620_),
    .S(_0660_),
    .Z(_0145_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1788_ (.I0(\mem[13][22] ),
    .I1(_0621_),
    .S(_0660_),
    .Z(_0146_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1789_ (.I0(\mem[13][23] ),
    .I1(_0622_),
    .S(_0660_),
    .Z(_0147_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1790_ (.I0(\mem[13][24] ),
    .I1(_0623_),
    .S(_0660_),
    .Z(_0148_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1791_ (.I0(\mem[13][25] ),
    .I1(_0624_),
    .S(_0660_),
    .Z(_0149_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1792_ (.I0(\mem[13][26] ),
    .I1(_0625_),
    .S(_0660_),
    .Z(_0150_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1793_ (.I0(\mem[13][27] ),
    .I1(_0626_),
    .S(_0660_),
    .Z(_0151_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _1794_ (.I(_0658_),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1795_ (.I0(\mem[13][28] ),
    .I1(_0627_),
    .S(_0661_),
    .Z(_0152_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1796_ (.I0(\mem[13][29] ),
    .I1(_0629_),
    .S(_0661_),
    .Z(_0153_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1797_ (.I0(\mem[13][2] ),
    .I1(_0630_),
    .S(_0661_),
    .Z(_0154_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1798_ (.I0(\mem[13][30] ),
    .I1(_0631_),
    .S(_0661_),
    .Z(_0155_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1799_ (.I0(\mem[13][31] ),
    .I1(_0632_),
    .S(_0661_),
    .Z(_0156_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1800_ (.I0(\mem[13][3] ),
    .I1(_0633_),
    .S(_0661_),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1801_ (.I0(\mem[13][4] ),
    .I1(_0634_),
    .S(_0661_),
    .Z(_0158_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1802_ (.I0(\mem[13][5] ),
    .I1(_0635_),
    .S(_0661_),
    .Z(_0159_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1803_ (.I0(\mem[13][6] ),
    .I1(_0636_),
    .S(_0661_),
    .Z(_0160_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1804_ (.I0(\mem[13][7] ),
    .I1(_0637_),
    .S(_0661_),
    .Z(_0161_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1805_ (.I0(\mem[13][8] ),
    .I1(_0638_),
    .S(_0658_),
    .Z(_0162_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1806_ (.I0(\mem[13][9] ),
    .I1(_0639_),
    .S(_0658_),
    .Z(_0163_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1807_ (.A1(_0568_),
    .A2(_0640_),
    .Z(_0662_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _1808_ (.A1(_0662_),
    .A2(_0651_),
    .Z(_0663_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _1809_ (.I(_0663_),
    .Z(_0664_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1810_ (.I0(\mem[14][0] ),
    .I1(_0599_),
    .S(_0664_),
    .Z(_0164_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1811_ (.I0(\mem[14][10] ),
    .I1(_0607_),
    .S(_0664_),
    .Z(_0165_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1812_ (.I0(\mem[14][11] ),
    .I1(_0608_),
    .S(_0664_),
    .Z(_0166_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1813_ (.I0(\mem[14][12] ),
    .I1(_0609_),
    .S(_0664_),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1814_ (.I0(\mem[14][13] ),
    .I1(_0610_),
    .S(_0664_),
    .Z(_0168_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1815_ (.I0(\mem[14][14] ),
    .I1(_0611_),
    .S(_0664_),
    .Z(_0169_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1816_ (.I0(\mem[14][15] ),
    .I1(_0612_),
    .S(_0664_),
    .Z(_0170_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1817_ (.I0(\mem[14][16] ),
    .I1(_0613_),
    .S(_0664_),
    .Z(_0171_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1818_ (.I0(\mem[14][17] ),
    .I1(_0614_),
    .S(_0664_),
    .Z(_0172_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1819_ (.I0(\mem[14][18] ),
    .I1(_0615_),
    .S(_0664_),
    .Z(_0173_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _1820_ (.I(_0663_),
    .Z(_0665_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1821_ (.I0(\mem[14][19] ),
    .I1(_0616_),
    .S(_0665_),
    .Z(_0174_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1822_ (.I0(\mem[14][1] ),
    .I1(_0618_),
    .S(_0665_),
    .Z(_0175_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1823_ (.I0(\mem[14][20] ),
    .I1(_0619_),
    .S(_0665_),
    .Z(_0176_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1824_ (.I0(\mem[14][21] ),
    .I1(_0620_),
    .S(_0665_),
    .Z(_0177_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1825_ (.I0(\mem[14][22] ),
    .I1(_0621_),
    .S(_0665_),
    .Z(_0178_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1826_ (.I0(\mem[14][23] ),
    .I1(_0622_),
    .S(_0665_),
    .Z(_0179_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1827_ (.I0(\mem[14][24] ),
    .I1(_0623_),
    .S(_0665_),
    .Z(_0180_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1828_ (.I0(\mem[14][25] ),
    .I1(_0624_),
    .S(_0665_),
    .Z(_0181_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1829_ (.I0(\mem[14][26] ),
    .I1(_0625_),
    .S(_0665_),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1830_ (.I0(\mem[14][27] ),
    .I1(_0626_),
    .S(_0665_),
    .Z(_0183_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1831_ (.I(_0663_),
    .Z(_0666_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1832_ (.I0(\mem[14][28] ),
    .I1(_0627_),
    .S(_0666_),
    .Z(_0184_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1833_ (.I0(\mem[14][29] ),
    .I1(_0629_),
    .S(_0666_),
    .Z(_0185_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1834_ (.I0(\mem[14][2] ),
    .I1(_0630_),
    .S(_0666_),
    .Z(_0186_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1835_ (.I0(\mem[14][30] ),
    .I1(_0631_),
    .S(_0666_),
    .Z(_0187_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1836_ (.I0(\mem[14][31] ),
    .I1(_0632_),
    .S(_0666_),
    .Z(_0188_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1837_ (.I0(\mem[14][3] ),
    .I1(_0633_),
    .S(_0666_),
    .Z(_0189_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1838_ (.I0(\mem[14][4] ),
    .I1(_0634_),
    .S(_0666_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1839_ (.I0(\mem[14][5] ),
    .I1(_0635_),
    .S(_0666_),
    .Z(_0191_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1840_ (.I0(\mem[14][6] ),
    .I1(_0636_),
    .S(_0666_),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1841_ (.I0(\mem[14][7] ),
    .I1(_0637_),
    .S(_0666_),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1842_ (.I0(\mem[14][8] ),
    .I1(_0638_),
    .S(_0663_),
    .Z(_0194_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1843_ (.I0(\mem[14][9] ),
    .I1(_0639_),
    .S(_0663_),
    .Z(_0195_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _1844_ (.A1(_0568_),
    .A2(_0646_),
    .Z(_0667_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _1845_ (.A1(_0667_),
    .A2(_0651_),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _1846_ (.I(_0668_),
    .Z(_0669_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1847_ (.I0(\mem[15][0] ),
    .I1(_0599_),
    .S(_0669_),
    .Z(_0196_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1848_ (.I0(\mem[15][10] ),
    .I1(_0607_),
    .S(_0669_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1849_ (.I0(\mem[15][11] ),
    .I1(_0608_),
    .S(_0669_),
    .Z(_0198_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1850_ (.I0(\mem[15][12] ),
    .I1(_0609_),
    .S(_0669_),
    .Z(_0199_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1851_ (.I0(\mem[15][13] ),
    .I1(_0610_),
    .S(_0669_),
    .Z(_0200_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1852_ (.I0(\mem[15][14] ),
    .I1(_0611_),
    .S(_0669_),
    .Z(_0201_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1853_ (.I0(\mem[15][15] ),
    .I1(_0612_),
    .S(_0669_),
    .Z(_0202_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1854_ (.I0(\mem[15][16] ),
    .I1(_0613_),
    .S(_0669_),
    .Z(_0203_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1855_ (.I0(\mem[15][17] ),
    .I1(_0614_),
    .S(_0669_),
    .Z(_0204_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1856_ (.I0(\mem[15][18] ),
    .I1(_0615_),
    .S(_0669_),
    .Z(_0205_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _1857_ (.I(_0668_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1858_ (.I0(\mem[15][19] ),
    .I1(_0616_),
    .S(_0670_),
    .Z(_0206_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1859_ (.I0(\mem[15][1] ),
    .I1(_0618_),
    .S(_0670_),
    .Z(_0207_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1860_ (.I0(\mem[15][20] ),
    .I1(_0619_),
    .S(_0670_),
    .Z(_0208_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1861_ (.I0(\mem[15][21] ),
    .I1(_0620_),
    .S(_0670_),
    .Z(_0209_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1862_ (.I0(\mem[15][22] ),
    .I1(_0621_),
    .S(_0670_),
    .Z(_0210_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1863_ (.I0(\mem[15][23] ),
    .I1(_0622_),
    .S(_0670_),
    .Z(_0211_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1864_ (.I0(\mem[15][24] ),
    .I1(_0623_),
    .S(_0670_),
    .Z(_0212_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1865_ (.I0(\mem[15][25] ),
    .I1(_0624_),
    .S(_0670_),
    .Z(_0213_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1866_ (.I0(\mem[15][26] ),
    .I1(_0625_),
    .S(_0670_),
    .Z(_0214_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1867_ (.I0(\mem[15][27] ),
    .I1(_0626_),
    .S(_0670_),
    .Z(_0215_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1868_ (.I(_0668_),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1869_ (.I0(\mem[15][28] ),
    .I1(_0627_),
    .S(_0671_),
    .Z(_0216_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1870_ (.I0(\mem[15][29] ),
    .I1(_0629_),
    .S(_0671_),
    .Z(_0217_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1871_ (.I0(\mem[15][2] ),
    .I1(_0630_),
    .S(_0671_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1872_ (.I0(\mem[15][30] ),
    .I1(_0631_),
    .S(_0671_),
    .Z(_0219_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1873_ (.I0(\mem[15][31] ),
    .I1(_0632_),
    .S(_0671_),
    .Z(_0220_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1874_ (.I0(\mem[15][3] ),
    .I1(_0633_),
    .S(_0671_),
    .Z(_0221_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1875_ (.I0(\mem[15][4] ),
    .I1(_0634_),
    .S(_0671_),
    .Z(_0222_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1876_ (.I0(\mem[15][5] ),
    .I1(_0635_),
    .S(_0671_),
    .Z(_0223_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1877_ (.I0(\mem[15][6] ),
    .I1(_0636_),
    .S(_0671_),
    .Z(_0224_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1878_ (.I0(\mem[15][7] ),
    .I1(_0637_),
    .S(_0671_),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1879_ (.I0(\mem[15][8] ),
    .I1(_0638_),
    .S(_0668_),
    .Z(_0226_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1880_ (.I0(\mem[15][9] ),
    .I1(_0639_),
    .S(_0668_),
    .Z(_0227_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _1881_ (.A1(_0602_),
    .A2(_0657_),
    .Z(_0672_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1882_ (.I(_0672_),
    .Z(_0673_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1883_ (.I0(\mem[1][0] ),
    .I1(_0599_),
    .S(_0673_),
    .Z(_0228_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1884_ (.I0(\mem[1][10] ),
    .I1(_0607_),
    .S(_0673_),
    .Z(_0229_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1885_ (.I0(\mem[1][11] ),
    .I1(_0608_),
    .S(_0673_),
    .Z(_0230_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1886_ (.I0(\mem[1][12] ),
    .I1(_0609_),
    .S(_0673_),
    .Z(_0231_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1887_ (.I0(\mem[1][13] ),
    .I1(_0610_),
    .S(_0673_),
    .Z(_0232_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1888_ (.I0(\mem[1][14] ),
    .I1(_0611_),
    .S(_0673_),
    .Z(_0233_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1889_ (.I0(\mem[1][15] ),
    .I1(_0612_),
    .S(_0673_),
    .Z(_0234_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1890_ (.I0(\mem[1][16] ),
    .I1(_0613_),
    .S(_0673_),
    .Z(_0235_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1891_ (.I0(\mem[1][17] ),
    .I1(_0614_),
    .S(_0673_),
    .Z(_0236_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1892_ (.I0(\mem[1][18] ),
    .I1(_0615_),
    .S(_0673_),
    .Z(_0237_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1893_ (.I(_0672_),
    .Z(_0674_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1894_ (.I0(\mem[1][19] ),
    .I1(_0616_),
    .S(_0674_),
    .Z(_0238_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1895_ (.I0(\mem[1][1] ),
    .I1(_0618_),
    .S(_0674_),
    .Z(_0239_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1896_ (.I0(\mem[1][20] ),
    .I1(_0619_),
    .S(_0674_),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1897_ (.I0(\mem[1][21] ),
    .I1(_0620_),
    .S(_0674_),
    .Z(_0241_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1898_ (.I0(\mem[1][22] ),
    .I1(_0621_),
    .S(_0674_),
    .Z(_0242_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1899_ (.I0(\mem[1][23] ),
    .I1(_0622_),
    .S(_0674_),
    .Z(_0243_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1900_ (.I0(\mem[1][24] ),
    .I1(_0623_),
    .S(_0674_),
    .Z(_0244_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1901_ (.I0(\mem[1][25] ),
    .I1(_0624_),
    .S(_0674_),
    .Z(_0245_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1902_ (.I0(\mem[1][26] ),
    .I1(_0625_),
    .S(_0674_),
    .Z(_0246_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1903_ (.I0(\mem[1][27] ),
    .I1(_0626_),
    .S(_0674_),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1904_ (.I(_0672_),
    .Z(_0675_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1905_ (.I0(\mem[1][28] ),
    .I1(_0627_),
    .S(_0675_),
    .Z(_0248_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1906_ (.I0(\mem[1][29] ),
    .I1(_0629_),
    .S(_0675_),
    .Z(_0249_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1907_ (.I0(\mem[1][2] ),
    .I1(_0630_),
    .S(_0675_),
    .Z(_0250_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1908_ (.I0(\mem[1][30] ),
    .I1(_0631_),
    .S(_0675_),
    .Z(_0251_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1909_ (.I0(\mem[1][31] ),
    .I1(_0632_),
    .S(_0675_),
    .Z(_0252_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1910_ (.I0(\mem[1][3] ),
    .I1(_0633_),
    .S(_0675_),
    .Z(_0253_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1911_ (.I0(\mem[1][4] ),
    .I1(_0634_),
    .S(_0675_),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1912_ (.I0(\mem[1][5] ),
    .I1(_0635_),
    .S(_0675_),
    .Z(_0255_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1913_ (.I0(\mem[1][6] ),
    .I1(_0636_),
    .S(_0675_),
    .Z(_0256_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1914_ (.I0(\mem[1][7] ),
    .I1(_0637_),
    .S(_0675_),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1915_ (.I0(\mem[1][8] ),
    .I1(_0638_),
    .S(_0672_),
    .Z(_0258_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1916_ (.I0(\mem[1][9] ),
    .I1(_0639_),
    .S(_0672_),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _1917_ (.A1(_0602_),
    .A2(_0662_),
    .Z(_0676_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1918_ (.I(_0676_),
    .Z(_0677_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1919_ (.I0(\mem[2][0] ),
    .I1(_0599_),
    .S(_0677_),
    .Z(_0260_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1920_ (.I0(\mem[2][10] ),
    .I1(_0607_),
    .S(_0677_),
    .Z(_0261_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1921_ (.I0(\mem[2][11] ),
    .I1(_0608_),
    .S(_0677_),
    .Z(_0262_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1922_ (.I0(\mem[2][12] ),
    .I1(_0609_),
    .S(_0677_),
    .Z(_0263_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1923_ (.I0(\mem[2][13] ),
    .I1(_0610_),
    .S(_0677_),
    .Z(_0264_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1924_ (.I0(\mem[2][14] ),
    .I1(_0611_),
    .S(_0677_),
    .Z(_0265_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1925_ (.I0(\mem[2][15] ),
    .I1(_0612_),
    .S(_0677_),
    .Z(_0266_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1926_ (.I0(\mem[2][16] ),
    .I1(_0613_),
    .S(_0677_),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1927_ (.I0(\mem[2][17] ),
    .I1(_0614_),
    .S(_0677_),
    .Z(_0268_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1928_ (.I0(\mem[2][18] ),
    .I1(_0615_),
    .S(_0677_),
    .Z(_0269_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _1929_ (.I(_0676_),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1930_ (.I0(\mem[2][19] ),
    .I1(_0616_),
    .S(_0678_),
    .Z(_0270_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1931_ (.I0(\mem[2][1] ),
    .I1(_0618_),
    .S(_0678_),
    .Z(_0271_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1932_ (.I0(\mem[2][20] ),
    .I1(_0619_),
    .S(_0678_),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1933_ (.I0(\mem[2][21] ),
    .I1(_0620_),
    .S(_0678_),
    .Z(_0273_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1934_ (.I0(\mem[2][22] ),
    .I1(_0621_),
    .S(_0678_),
    .Z(_0274_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1935_ (.I0(\mem[2][23] ),
    .I1(_0622_),
    .S(_0678_),
    .Z(_0275_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1936_ (.I0(\mem[2][24] ),
    .I1(_0623_),
    .S(_0678_),
    .Z(_0276_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1937_ (.I0(\mem[2][25] ),
    .I1(_0624_),
    .S(_0678_),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1938_ (.I0(\mem[2][26] ),
    .I1(_0625_),
    .S(_0678_),
    .Z(_0278_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1939_ (.I0(\mem[2][27] ),
    .I1(_0626_),
    .S(_0678_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1940_ (.I(_0676_),
    .Z(_0679_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1941_ (.I0(\mem[2][28] ),
    .I1(_0627_),
    .S(_0679_),
    .Z(_0280_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1942_ (.I0(\mem[2][29] ),
    .I1(_0629_),
    .S(_0679_),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1943_ (.I0(\mem[2][2] ),
    .I1(_0630_),
    .S(_0679_),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1944_ (.I0(\mem[2][30] ),
    .I1(_0631_),
    .S(_0679_),
    .Z(_0283_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1945_ (.I0(\mem[2][31] ),
    .I1(_0632_),
    .S(_0679_),
    .Z(_0284_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1946_ (.I0(\mem[2][3] ),
    .I1(_0633_),
    .S(_0679_),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1947_ (.I0(\mem[2][4] ),
    .I1(_0634_),
    .S(_0679_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1948_ (.I0(\mem[2][5] ),
    .I1(_0635_),
    .S(_0679_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1949_ (.I0(\mem[2][6] ),
    .I1(_0636_),
    .S(_0679_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1950_ (.I0(\mem[2][7] ),
    .I1(_0637_),
    .S(_0679_),
    .Z(_0289_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1951_ (.I0(\mem[2][8] ),
    .I1(_0638_),
    .S(_0676_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1952_ (.I0(\mem[2][9] ),
    .I1(_0639_),
    .S(_0676_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _1953_ (.A1(_0602_),
    .A2(_0667_),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1954_ (.I(_0680_),
    .Z(_0681_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1955_ (.I0(\mem[3][0] ),
    .I1(_0599_),
    .S(_0681_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1956_ (.I0(\mem[3][10] ),
    .I1(_0607_),
    .S(_0681_),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1957_ (.I0(\mem[3][11] ),
    .I1(_0608_),
    .S(_0681_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1958_ (.I0(\mem[3][12] ),
    .I1(_0609_),
    .S(_0681_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1959_ (.I0(\mem[3][13] ),
    .I1(_0610_),
    .S(_0681_),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1960_ (.I0(\mem[3][14] ),
    .I1(_0611_),
    .S(_0681_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1961_ (.I0(\mem[3][15] ),
    .I1(_0612_),
    .S(_0681_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1962_ (.I0(\mem[3][16] ),
    .I1(_0613_),
    .S(_0681_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1963_ (.I0(\mem[3][17] ),
    .I1(_0614_),
    .S(_0681_),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1964_ (.I0(\mem[3][18] ),
    .I1(_0615_),
    .S(_0681_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _1965_ (.I(_0680_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1966_ (.I0(\mem[3][19] ),
    .I1(_0616_),
    .S(_0682_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1967_ (.I0(\mem[3][1] ),
    .I1(_0618_),
    .S(_0682_),
    .Z(_0303_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1968_ (.I0(\mem[3][20] ),
    .I1(_0619_),
    .S(_0682_),
    .Z(_0304_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1969_ (.I0(\mem[3][21] ),
    .I1(_0620_),
    .S(_0682_),
    .Z(_0305_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1970_ (.I0(\mem[3][22] ),
    .I1(_0621_),
    .S(_0682_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1971_ (.I0(\mem[3][23] ),
    .I1(_0622_),
    .S(_0682_),
    .Z(_0307_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1972_ (.I0(\mem[3][24] ),
    .I1(_0623_),
    .S(_0682_),
    .Z(_0308_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1973_ (.I0(\mem[3][25] ),
    .I1(_0624_),
    .S(_0682_),
    .Z(_0309_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1974_ (.I0(\mem[3][26] ),
    .I1(_0625_),
    .S(_0682_),
    .Z(_0310_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1975_ (.I0(\mem[3][27] ),
    .I1(_0626_),
    .S(_0682_),
    .Z(_0311_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1976_ (.I(_0680_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1977_ (.I0(\mem[3][28] ),
    .I1(_0627_),
    .S(_0683_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1978_ (.I0(\mem[3][29] ),
    .I1(_0629_),
    .S(_0683_),
    .Z(_0313_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1979_ (.I0(\mem[3][2] ),
    .I1(_0630_),
    .S(_0683_),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1980_ (.I0(\mem[3][30] ),
    .I1(_0631_),
    .S(_0683_),
    .Z(_0315_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1981_ (.I0(\mem[3][31] ),
    .I1(_0632_),
    .S(_0683_),
    .Z(_0316_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1982_ (.I0(\mem[3][3] ),
    .I1(_0633_),
    .S(_0683_),
    .Z(_0317_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1983_ (.I0(\mem[3][4] ),
    .I1(_0634_),
    .S(_0683_),
    .Z(_0318_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1984_ (.I0(\mem[3][5] ),
    .I1(_0635_),
    .S(_0683_),
    .Z(_0319_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1985_ (.I0(\mem[3][6] ),
    .I1(_0636_),
    .S(_0683_),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1986_ (.I0(\mem[3][7] ),
    .I1(_0637_),
    .S(_0683_),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1987_ (.I0(\mem[3][8] ),
    .I1(_0638_),
    .S(_0680_),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1988_ (.I0(\mem[3][9] ),
    .I1(_0639_),
    .S(_0680_),
    .Z(_0323_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _1989_ (.A1(\wr_ptr_bin[2] ),
    .A2(_0601_),
    .A3(_0568_),
    .Z(_0684_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _1990_ (.A1(_0603_),
    .A2(_0684_),
    .Z(_0685_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _1991_ (.I(_0685_),
    .Z(_0686_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1992_ (.I0(\mem[4][0] ),
    .I1(net5),
    .S(_0686_),
    .Z(_0324_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1993_ (.I0(\mem[4][10] ),
    .I1(net6),
    .S(_0686_),
    .Z(_0325_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1994_ (.I0(\mem[4][11] ),
    .I1(net7),
    .S(_0686_),
    .Z(_0326_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1995_ (.I0(\mem[4][12] ),
    .I1(net8),
    .S(_0686_),
    .Z(_0327_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1996_ (.I0(\mem[4][13] ),
    .I1(net9),
    .S(_0686_),
    .Z(_0328_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1997_ (.I0(\mem[4][14] ),
    .I1(net10),
    .S(_0686_),
    .Z(_0329_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1998_ (.I0(\mem[4][15] ),
    .I1(net11),
    .S(_0686_),
    .Z(_0330_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _1999_ (.I0(\mem[4][16] ),
    .I1(net12),
    .S(_0686_),
    .Z(_0331_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2000_ (.I0(\mem[4][17] ),
    .I1(net13),
    .S(_0686_),
    .Z(_0332_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2001_ (.I0(\mem[4][18] ),
    .I1(net14),
    .S(_0686_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2002_ (.I(_0685_),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2003_ (.I0(\mem[4][19] ),
    .I1(net15),
    .S(_0687_),
    .Z(_0334_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2004_ (.I0(\mem[4][1] ),
    .I1(net16),
    .S(_0687_),
    .Z(_0335_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2005_ (.I0(\mem[4][20] ),
    .I1(net17),
    .S(_0687_),
    .Z(_0336_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2006_ (.I0(\mem[4][21] ),
    .I1(net18),
    .S(_0687_),
    .Z(_0337_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2007_ (.I0(\mem[4][22] ),
    .I1(net19),
    .S(_0687_),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2008_ (.I0(\mem[4][23] ),
    .I1(net20),
    .S(_0687_),
    .Z(_0339_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2009_ (.I0(\mem[4][24] ),
    .I1(net21),
    .S(_0687_),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2010_ (.I0(\mem[4][25] ),
    .I1(net22),
    .S(_0687_),
    .Z(_0341_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2011_ (.I0(\mem[4][26] ),
    .I1(net23),
    .S(_0687_),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2012_ (.I0(\mem[4][27] ),
    .I1(net24),
    .S(_0687_),
    .Z(_0343_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2013_ (.I(_0685_),
    .Z(_0688_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2014_ (.I0(\mem[4][28] ),
    .I1(net25),
    .S(_0688_),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2015_ (.I0(\mem[4][29] ),
    .I1(net26),
    .S(_0688_),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2016_ (.I0(\mem[4][2] ),
    .I1(net27),
    .S(_0688_),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2017_ (.I0(\mem[4][30] ),
    .I1(net28),
    .S(_0688_),
    .Z(_0347_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2018_ (.I0(\mem[4][31] ),
    .I1(net29),
    .S(_0688_),
    .Z(_0348_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2019_ (.I0(\mem[4][3] ),
    .I1(net30),
    .S(_0688_),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2020_ (.I0(\mem[4][4] ),
    .I1(net31),
    .S(_0688_),
    .Z(_0350_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2021_ (.I0(\mem[4][5] ),
    .I1(net32),
    .S(_0688_),
    .Z(_0351_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2022_ (.I0(\mem[4][6] ),
    .I1(net33),
    .S(_0688_),
    .Z(_0352_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2023_ (.I0(\mem[4][7] ),
    .I1(net34),
    .S(_0688_),
    .Z(_0353_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2024_ (.I0(\mem[4][8] ),
    .I1(net35),
    .S(_0685_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2025_ (.I0(\mem[4][9] ),
    .I1(net36),
    .S(_0685_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _2026_ (.A1(_0656_),
    .A2(_0684_),
    .Z(_0689_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2027_ (.I(_0689_),
    .Z(_0690_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2028_ (.I0(\mem[5][0] ),
    .I1(net5),
    .S(_0690_),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2029_ (.I0(\mem[5][10] ),
    .I1(net6),
    .S(_0690_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2030_ (.I0(\mem[5][11] ),
    .I1(net7),
    .S(_0690_),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2031_ (.I0(\mem[5][12] ),
    .I1(net8),
    .S(_0690_),
    .Z(_0359_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2032_ (.I0(\mem[5][13] ),
    .I1(net9),
    .S(_0690_),
    .Z(_0360_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2033_ (.I0(\mem[5][14] ),
    .I1(net10),
    .S(_0690_),
    .Z(_0361_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2034_ (.I0(\mem[5][15] ),
    .I1(net11),
    .S(_0690_),
    .Z(_0362_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2035_ (.I0(\mem[5][16] ),
    .I1(net12),
    .S(_0690_),
    .Z(_0363_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2036_ (.I0(\mem[5][17] ),
    .I1(net13),
    .S(_0690_),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2037_ (.I0(\mem[5][18] ),
    .I1(net14),
    .S(_0690_),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2038_ (.I(_0689_),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2039_ (.I0(\mem[5][19] ),
    .I1(net15),
    .S(_0691_),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2040_ (.I0(\mem[5][1] ),
    .I1(net16),
    .S(_0691_),
    .Z(_0367_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2041_ (.I0(\mem[5][20] ),
    .I1(net17),
    .S(_0691_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2042_ (.I0(\mem[5][21] ),
    .I1(net18),
    .S(_0691_),
    .Z(_0369_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2043_ (.I0(\mem[5][22] ),
    .I1(net19),
    .S(_0691_),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2044_ (.I0(\mem[5][23] ),
    .I1(net20),
    .S(_0691_),
    .Z(_0371_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2045_ (.I0(\mem[5][24] ),
    .I1(net21),
    .S(_0691_),
    .Z(_0372_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2046_ (.I0(\mem[5][25] ),
    .I1(net22),
    .S(_0691_),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2047_ (.I0(\mem[5][26] ),
    .I1(net23),
    .S(_0691_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2048_ (.I0(\mem[5][27] ),
    .I1(net24),
    .S(_0691_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2049_ (.I(_0689_),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2050_ (.I0(\mem[5][28] ),
    .I1(net25),
    .S(_0692_),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2051_ (.I0(\mem[5][29] ),
    .I1(net26),
    .S(_0692_),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2052_ (.I0(\mem[5][2] ),
    .I1(net27),
    .S(_0692_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2053_ (.I0(\mem[5][30] ),
    .I1(net28),
    .S(_0692_),
    .Z(_0379_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2054_ (.I0(\mem[5][31] ),
    .I1(net29),
    .S(_0692_),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2055_ (.I0(\mem[5][3] ),
    .I1(net30),
    .S(_0692_),
    .Z(_0381_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2056_ (.I0(\mem[5][4] ),
    .I1(net31),
    .S(_0692_),
    .Z(_0382_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2057_ (.I0(\mem[5][5] ),
    .I1(net32),
    .S(_0692_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2058_ (.I0(\mem[5][6] ),
    .I1(net33),
    .S(_0692_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2059_ (.I0(\mem[5][7] ),
    .I1(net34),
    .S(_0692_),
    .Z(_0385_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2060_ (.I0(\mem[5][8] ),
    .I1(net35),
    .S(_0689_),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2061_ (.I0(\mem[5][9] ),
    .I1(net36),
    .S(_0689_),
    .Z(_0387_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _2062_ (.A1(_0640_),
    .A2(_0684_),
    .Z(_0693_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2063_ (.I(_0693_),
    .Z(_0694_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2064_ (.I0(\mem[6][0] ),
    .I1(net5),
    .S(_0694_),
    .Z(_0388_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2065_ (.I0(\mem[6][10] ),
    .I1(net6),
    .S(_0694_),
    .Z(_0389_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2066_ (.I0(\mem[6][11] ),
    .I1(net7),
    .S(_0694_),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2067_ (.I0(\mem[6][12] ),
    .I1(net8),
    .S(_0694_),
    .Z(_0391_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2068_ (.I0(\mem[6][13] ),
    .I1(net9),
    .S(_0694_),
    .Z(_0392_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2069_ (.I0(\mem[6][14] ),
    .I1(net10),
    .S(_0694_),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2070_ (.I0(\mem[6][15] ),
    .I1(net11),
    .S(_0694_),
    .Z(_0394_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2071_ (.I0(\mem[6][16] ),
    .I1(net12),
    .S(_0694_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2072_ (.I0(\mem[6][17] ),
    .I1(net13),
    .S(_0694_),
    .Z(_0396_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2073_ (.I0(\mem[6][18] ),
    .I1(net14),
    .S(_0694_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2074_ (.I(_0693_),
    .Z(_0695_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2075_ (.I0(\mem[6][19] ),
    .I1(net15),
    .S(_0695_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2076_ (.I0(\mem[6][1] ),
    .I1(net16),
    .S(_0695_),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2077_ (.I0(\mem[6][20] ),
    .I1(net17),
    .S(_0695_),
    .Z(_0400_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2078_ (.I0(\mem[6][21] ),
    .I1(net18),
    .S(_0695_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2079_ (.I0(\mem[6][22] ),
    .I1(net19),
    .S(_0695_),
    .Z(_0402_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2080_ (.I0(\mem[6][23] ),
    .I1(net20),
    .S(_0695_),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2081_ (.I0(\mem[6][24] ),
    .I1(net21),
    .S(_0695_),
    .Z(_0404_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2082_ (.I0(\mem[6][25] ),
    .I1(net22),
    .S(_0695_),
    .Z(_0405_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2083_ (.I0(\mem[6][26] ),
    .I1(net23),
    .S(_0695_),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2084_ (.I0(\mem[6][27] ),
    .I1(net24),
    .S(_0695_),
    .Z(_0407_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2085_ (.I(_0693_),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2086_ (.I0(\mem[6][28] ),
    .I1(net25),
    .S(_0696_),
    .Z(_0408_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2087_ (.I0(\mem[6][29] ),
    .I1(net26),
    .S(_0696_),
    .Z(_0409_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2088_ (.I0(\mem[6][2] ),
    .I1(net27),
    .S(_0696_),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2089_ (.I0(\mem[6][30] ),
    .I1(net28),
    .S(_0696_),
    .Z(_0411_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2090_ (.I0(\mem[6][31] ),
    .I1(net29),
    .S(_0696_),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2091_ (.I0(\mem[6][3] ),
    .I1(net30),
    .S(_0696_),
    .Z(_0413_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2092_ (.I0(\mem[6][4] ),
    .I1(net31),
    .S(_0696_),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2093_ (.I0(\mem[6][5] ),
    .I1(net32),
    .S(_0696_),
    .Z(_0415_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2094_ (.I0(\mem[6][6] ),
    .I1(net33),
    .S(_0696_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2095_ (.I0(\mem[6][7] ),
    .I1(net34),
    .S(_0696_),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2096_ (.I0(\mem[6][8] ),
    .I1(net35),
    .S(_0693_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2097_ (.I0(\mem[6][9] ),
    .I1(net36),
    .S(_0693_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _2098_ (.A1(_0646_),
    .A2(_0684_),
    .Z(_0697_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2099_ (.I(_0697_),
    .Z(_0698_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2100_ (.I0(\mem[7][0] ),
    .I1(net5),
    .S(_0698_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2101_ (.I0(\mem[7][10] ),
    .I1(net6),
    .S(_0698_),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2102_ (.I0(\mem[7][11] ),
    .I1(net7),
    .S(_0698_),
    .Z(_0422_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2103_ (.I0(\mem[7][12] ),
    .I1(net8),
    .S(_0698_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2104_ (.I0(\mem[7][13] ),
    .I1(net9),
    .S(_0698_),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2105_ (.I0(\mem[7][14] ),
    .I1(net10),
    .S(_0698_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2106_ (.I0(\mem[7][15] ),
    .I1(net11),
    .S(_0698_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2107_ (.I0(\mem[7][16] ),
    .I1(net12),
    .S(_0698_),
    .Z(_0427_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2108_ (.I0(\mem[7][17] ),
    .I1(net13),
    .S(_0698_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2109_ (.I0(\mem[7][18] ),
    .I1(net14),
    .S(_0698_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2110_ (.I(_0697_),
    .Z(_0699_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2111_ (.I0(\mem[7][19] ),
    .I1(net15),
    .S(_0699_),
    .Z(_0430_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2112_ (.I0(\mem[7][1] ),
    .I1(net16),
    .S(_0699_),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2113_ (.I0(\mem[7][20] ),
    .I1(net17),
    .S(_0699_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2114_ (.I0(\mem[7][21] ),
    .I1(net18),
    .S(_0699_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2115_ (.I0(\mem[7][22] ),
    .I1(net19),
    .S(_0699_),
    .Z(_0434_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2116_ (.I0(\mem[7][23] ),
    .I1(net20),
    .S(_0699_),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2117_ (.I0(\mem[7][24] ),
    .I1(net21),
    .S(_0699_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2118_ (.I0(\mem[7][25] ),
    .I1(net22),
    .S(_0699_),
    .Z(_0437_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2119_ (.I0(\mem[7][26] ),
    .I1(net23),
    .S(_0699_),
    .Z(_0438_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2120_ (.I0(\mem[7][27] ),
    .I1(net24),
    .S(_0699_),
    .Z(_0439_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2121_ (.I(_0697_),
    .Z(_0700_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2122_ (.I0(\mem[7][28] ),
    .I1(net25),
    .S(_0700_),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2123_ (.I0(\mem[7][29] ),
    .I1(net26),
    .S(_0700_),
    .Z(_0441_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2124_ (.I0(\mem[7][2] ),
    .I1(net27),
    .S(_0700_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2125_ (.I0(\mem[7][30] ),
    .I1(net28),
    .S(_0700_),
    .Z(_0443_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2126_ (.I0(\mem[7][31] ),
    .I1(net29),
    .S(_0700_),
    .Z(_0444_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2127_ (.I0(\mem[7][3] ),
    .I1(net30),
    .S(_0700_),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2128_ (.I0(\mem[7][4] ),
    .I1(net31),
    .S(_0700_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2129_ (.I0(\mem[7][5] ),
    .I1(net32),
    .S(_0700_),
    .Z(_0447_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2130_ (.I0(\mem[7][6] ),
    .I1(net33),
    .S(_0700_),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2131_ (.I0(\mem[7][7] ),
    .I1(net34),
    .S(_0700_),
    .Z(_0449_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2132_ (.I0(\mem[7][8] ),
    .I1(net35),
    .S(_0697_),
    .Z(_0450_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2133_ (.I0(\mem[7][9] ),
    .I1(net36),
    .S(_0697_),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _2134_ (.A1(_0603_),
    .A2(_0641_),
    .Z(_0701_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2135_ (.I(_0701_),
    .Z(_0702_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2136_ (.I0(\mem[8][0] ),
    .I1(net5),
    .S(_0702_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2137_ (.I0(\mem[8][10] ),
    .I1(net6),
    .S(_0702_),
    .Z(_0453_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2138_ (.I0(\mem[8][11] ),
    .I1(net7),
    .S(_0702_),
    .Z(_0454_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2139_ (.I0(\mem[8][12] ),
    .I1(net8),
    .S(_0702_),
    .Z(_0455_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2140_ (.I0(\mem[8][13] ),
    .I1(net9),
    .S(_0702_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2141_ (.I0(\mem[8][14] ),
    .I1(net10),
    .S(_0702_),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2142_ (.I0(\mem[8][15] ),
    .I1(net11),
    .S(_0702_),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2143_ (.I0(\mem[8][16] ),
    .I1(net12),
    .S(_0702_),
    .Z(_0459_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2144_ (.I0(\mem[8][17] ),
    .I1(net13),
    .S(_0702_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2145_ (.I0(\mem[8][18] ),
    .I1(net14),
    .S(_0702_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2146_ (.I(_0701_),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2147_ (.I0(\mem[8][19] ),
    .I1(net15),
    .S(_0703_),
    .Z(_0462_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2148_ (.I0(\mem[8][1] ),
    .I1(net16),
    .S(_0703_),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2149_ (.I0(\mem[8][20] ),
    .I1(net17),
    .S(_0703_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2150_ (.I0(\mem[8][21] ),
    .I1(net18),
    .S(_0703_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2151_ (.I0(\mem[8][22] ),
    .I1(net19),
    .S(_0703_),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2152_ (.I0(\mem[8][23] ),
    .I1(net20),
    .S(_0703_),
    .Z(_0467_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2153_ (.I0(\mem[8][24] ),
    .I1(net21),
    .S(_0703_),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2154_ (.I0(\mem[8][25] ),
    .I1(net22),
    .S(_0703_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2155_ (.I0(\mem[8][26] ),
    .I1(net23),
    .S(_0703_),
    .Z(_0470_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2156_ (.I0(\mem[8][27] ),
    .I1(net24),
    .S(_0703_),
    .Z(_0471_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2157_ (.I(_0701_),
    .Z(_0704_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2158_ (.I0(\mem[8][28] ),
    .I1(net25),
    .S(_0704_),
    .Z(_0472_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2159_ (.I0(\mem[8][29] ),
    .I1(net26),
    .S(_0704_),
    .Z(_0473_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2160_ (.I0(\mem[8][2] ),
    .I1(net27),
    .S(_0704_),
    .Z(_0474_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2161_ (.I0(\mem[8][30] ),
    .I1(net28),
    .S(_0704_),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2162_ (.I0(\mem[8][31] ),
    .I1(net29),
    .S(_0704_),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2163_ (.I0(\mem[8][3] ),
    .I1(net30),
    .S(_0704_),
    .Z(_0477_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2164_ (.I0(\mem[8][4] ),
    .I1(net31),
    .S(_0704_),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2165_ (.I0(\mem[8][5] ),
    .I1(net32),
    .S(_0704_),
    .Z(_0479_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2166_ (.I0(\mem[8][6] ),
    .I1(net33),
    .S(_0704_),
    .Z(_0480_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2167_ (.I0(\mem[8][7] ),
    .I1(net34),
    .S(_0704_),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2168_ (.I0(\mem[8][8] ),
    .I1(net35),
    .S(_0701_),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2169_ (.I0(\mem[8][9] ),
    .I1(net36),
    .S(_0701_),
    .Z(_0483_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _2170_ (.A1(_0641_),
    .A2(_0656_),
    .Z(_0705_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2171_ (.I(_0705_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2172_ (.I0(\mem[9][0] ),
    .I1(net5),
    .S(_0706_),
    .Z(_0484_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2173_ (.I0(\mem[9][10] ),
    .I1(net6),
    .S(_0706_),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2174_ (.I0(\mem[9][11] ),
    .I1(net7),
    .S(_0706_),
    .Z(_0486_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2175_ (.I0(\mem[9][12] ),
    .I1(net8),
    .S(_0706_),
    .Z(_0487_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2176_ (.I0(\mem[9][13] ),
    .I1(net9),
    .S(_0706_),
    .Z(_0488_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2177_ (.I0(\mem[9][14] ),
    .I1(net10),
    .S(_0706_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2178_ (.I0(\mem[9][15] ),
    .I1(net11),
    .S(_0706_),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2179_ (.I0(\mem[9][16] ),
    .I1(net12),
    .S(_0706_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2180_ (.I0(\mem[9][17] ),
    .I1(net13),
    .S(_0706_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2181_ (.I0(\mem[9][18] ),
    .I1(net14),
    .S(_0706_),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2182_ (.I(_0705_),
    .Z(_0707_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2183_ (.I0(\mem[9][19] ),
    .I1(net15),
    .S(_0707_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2184_ (.I0(\mem[9][1] ),
    .I1(net16),
    .S(_0707_),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2185_ (.I0(\mem[9][20] ),
    .I1(net17),
    .S(_0707_),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2186_ (.I0(\mem[9][21] ),
    .I1(net18),
    .S(_0707_),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2187_ (.I0(\mem[9][22] ),
    .I1(net19),
    .S(_0707_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2188_ (.I0(\mem[9][23] ),
    .I1(net20),
    .S(_0707_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2189_ (.I0(\mem[9][24] ),
    .I1(net21),
    .S(_0707_),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2190_ (.I0(\mem[9][25] ),
    .I1(net22),
    .S(_0707_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2191_ (.I0(\mem[9][26] ),
    .I1(net23),
    .S(_0707_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2192_ (.I0(\mem[9][27] ),
    .I1(net24),
    .S(_0707_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2193_ (.I(_0705_),
    .Z(_0708_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2194_ (.I0(\mem[9][28] ),
    .I1(net25),
    .S(_0708_),
    .Z(_0504_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2195_ (.I0(\mem[9][29] ),
    .I1(net26),
    .S(_0708_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2196_ (.I0(\mem[9][2] ),
    .I1(net27),
    .S(_0708_),
    .Z(_0506_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2197_ (.I0(\mem[9][30] ),
    .I1(net28),
    .S(_0708_),
    .Z(_0507_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2198_ (.I0(\mem[9][31] ),
    .I1(net29),
    .S(_0708_),
    .Z(_0508_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2199_ (.I0(\mem[9][3] ),
    .I1(net30),
    .S(_0708_),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2200_ (.I0(\mem[9][4] ),
    .I1(net31),
    .S(_0708_),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2201_ (.I0(\mem[9][5] ),
    .I1(net32),
    .S(_0708_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2202_ (.I0(\mem[9][6] ),
    .I1(net33),
    .S(_0708_),
    .Z(_0512_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2203_ (.I0(\mem[9][7] ),
    .I1(net34),
    .S(_0708_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2204_ (.I0(\mem[9][8] ),
    .I1(net35),
    .S(_0705_),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2205_ (.I0(\mem[9][9] ),
    .I1(net36),
    .S(_0705_),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2206_ (.I(_0595_),
    .Z(_0709_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2207_ (.I(_1519_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2208_ (.I(_1514_),
    .Z(_0711_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2209_ (.I(_1517_),
    .Z(_0712_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2210_ (.A1(_0710_),
    .A2(\mem[15][0] ),
    .B1(\mem[12][0] ),
    .B2(_0711_),
    .C1(_0712_),
    .C2(\mem[13][0] ),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2211_ (.I(_1515_),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2212_ (.A1(\mem[6][0] ),
    .A2(_0714_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2213_ (.I(_0597_),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2214_ (.I0(_0713_),
    .I1(_0715_),
    .S(_0716_),
    .Z(_0717_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2215_ (.A1(_0709_),
    .A2(_0717_),
    .Z(_0718_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2216_ (.I(\rd_ptr_bin[3] ),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2217_ (.I(_0719_),
    .Z(_0720_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2218_ (.I(_1514_),
    .Z(_0721_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2219_ (.I(_0721_),
    .Z(_0722_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2220_ (.I(_1515_),
    .Z(_0723_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2221_ (.I(_0723_),
    .Z(_0724_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2222_ (.A1(\mem[8][0] ),
    .A2(_0722_),
    .B1(_0724_),
    .B2(\mem[10][0] ),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2223_ (.I(_1517_),
    .Z(_0726_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2224_ (.I(_0726_),
    .Z(_0727_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2225_ (.I(\rd_ptr_bin[2] ),
    .Z(_0728_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2226_ (.I(_0728_),
    .Z(_0729_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2227_ (.A1(\mem[9][0] ),
    .A2(_0727_),
    .B(_0729_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2228_ (.I(_0723_),
    .Z(_0731_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2229_ (.A1(\mem[14][0] ),
    .A2(_0731_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2230_ (.I(_0728_),
    .Z(_0733_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2231_ (.I(_0733_),
    .Z(_0734_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2232_ (.A1(_0725_),
    .A2(_0730_),
    .B1(_0732_),
    .B2(_0734_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2233_ (.I(\mem[7][0] ),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _2234_ (.A1(_0597_),
    .A2(_0728_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2235_ (.I(_0737_),
    .Z(_0738_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _2236_ (.A1(\rd_ptr_bin[3] ),
    .A2(_0594_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2237_ (.I(_0739_),
    .Z(_0740_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2238_ (.I(\mem[11][0] ),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2239_ (.A1(_0736_),
    .A2(_0738_),
    .B1(_0740_),
    .B2(_0741_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2240_ (.I(_0710_),
    .Z(_0743_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2241_ (.I(_0743_),
    .Z(_0744_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2242_ (.A1(_0720_),
    .A2(_0735_),
    .B1(_0742_),
    .B2(_0744_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2243_ (.I(_1519_),
    .Z(_0746_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2244_ (.I(_1517_),
    .Z(_0747_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2245_ (.A1(_0746_),
    .A2(\mem[3][0] ),
    .B1(\mem[1][0] ),
    .B2(_0747_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2246_ (.A1(\mem[2][0] ),
    .A2(_0724_),
    .B(_0729_),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2247_ (.A1(\mem[4][0] ),
    .A2(_0722_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2248_ (.A1(_0748_),
    .A2(_0749_),
    .B1(_0750_),
    .B2(_0729_),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2249_ (.A1(_0597_),
    .A2(_0728_),
    .A3(_1517_),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2250_ (.I(_0752_),
    .Z(_0753_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2251_ (.I(_1514_),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _2252_ (.A1(\rd_ptr_bin[3] ),
    .A2(\rd_ptr_bin[2] ),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2253_ (.A1(_0754_),
    .A2(_0755_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _2254_ (.A1(_1519_),
    .A2(_1515_),
    .A3(_1517_),
    .A4(_0756_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2255_ (.I(_0757_),
    .Z(_0758_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2256_ (.A1(_1499_),
    .A2(_0751_),
    .B1(_0753_),
    .B2(\mem[5][0] ),
    .C(_0758_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2257_ (.A1(_0718_),
    .A2(_0745_),
    .A3(_0759_),
    .Z(_0760_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _2258_ (.A1(net3),
    .A2(_0593_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2259_ (.I(_0761_),
    .Z(_0762_));
 gf180mcu_fd_sc_mcu9t5v0__or4_4 _2260_ (.A1(_0710_),
    .A2(_0723_),
    .A3(_1517_),
    .A4(_0756_),
    .Z(_0763_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2261_ (.I(_0763_),
    .Z(_0764_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2262_ (.I(_0764_),
    .Z(_0765_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2263_ (.A1(\mem[0][0] ),
    .A2(_0765_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2264_ (.A1(net45),
    .A2(_0762_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2265_ (.A1(_0760_),
    .A2(_0762_),
    .A3(_0766_),
    .B(_0767_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2266_ (.I(_0761_),
    .Z(_0768_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2267_ (.A1(_0743_),
    .A2(\mem[15][10] ),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2268_ (.A1(\mem[6][10] ),
    .A2(_0731_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2269_ (.I(_0711_),
    .Z(_0771_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2270_ (.A1(\mem[8][10] ),
    .A2(_0771_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2271_ (.A1(\mem[1][10] ),
    .A2(_0727_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2272_ (.I(_0598_),
    .Z(_0774_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2273_ (.I0(_0769_),
    .I1(_0770_),
    .I2(_0772_),
    .I3(_0773_),
    .S0(_0774_),
    .S1(_0709_),
    .Z(_0775_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2274_ (.I(_0712_),
    .Z(_0776_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2275_ (.A1(\mem[13][10] ),
    .A2(_0776_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2276_ (.I(_0723_),
    .Z(_0778_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2277_ (.A1(\mem[10][10] ),
    .A2(_0778_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2278_ (.I(_1514_),
    .Z(_0780_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2279_ (.A1(\mem[4][10] ),
    .A2(_0780_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2280_ (.I(_0710_),
    .Z(_0782_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2281_ (.A1(_0782_),
    .A2(\mem[3][10] ),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2282_ (.I(_0595_),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2283_ (.I0(_0777_),
    .I1(_0779_),
    .I2(_0781_),
    .I3(_0783_),
    .S0(_0784_),
    .S1(_1499_),
    .Z(_0785_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2284_ (.I(\mem[7][10] ),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2285_ (.I(_0739_),
    .Z(_0787_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2286_ (.I(\mem[11][10] ),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2287_ (.A1(_0786_),
    .A2(_0738_),
    .B1(_0787_),
    .B2(_0788_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2288_ (.I(_0755_),
    .Z(_0790_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2289_ (.A1(\rd_ptr_bin[3] ),
    .A2(\rd_ptr_bin[2] ),
    .Z(_0791_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2290_ (.I(_0791_),
    .Z(_0792_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2291_ (.A1(\mem[2][10] ),
    .A2(_0790_),
    .B1(_0792_),
    .B2(\mem[14][10] ),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2292_ (.I(_0793_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2293_ (.I(_0731_),
    .Z(_0795_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2294_ (.A1(_0744_),
    .A2(_0789_),
    .B1(_0794_),
    .B2(_0795_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2295_ (.A1(_0733_),
    .A2(\mem[12][10] ),
    .A3(_0721_),
    .Z(_0797_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2296_ (.A1(_0595_),
    .A2(\mem[9][10] ),
    .A3(_0726_),
    .Z(_0798_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2297_ (.A1(_0797_),
    .A2(_0798_),
    .Z(_0799_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2298_ (.I(_0719_),
    .Z(_0800_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2299_ (.A1(\mem[5][10] ),
    .A2(_0753_),
    .B1(_0799_),
    .B2(_0800_),
    .C(_0758_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2300_ (.A1(_0775_),
    .A2(_0785_),
    .A3(_0796_),
    .A4(_0801_),
    .Z(_0802_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2301_ (.A1(\mem[0][10] ),
    .A2(_0765_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2302_ (.A1(net46),
    .A2(_0762_),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2303_ (.A1(_0768_),
    .A2(_0802_),
    .A3(_0803_),
    .B(_0804_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _2304_ (.A1(_0594_),
    .A2(_1519_),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2305_ (.I(_0805_),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2306_ (.I(_0719_),
    .Z(_0807_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2307_ (.A1(\mem[3][11] ),
    .A2(_0806_),
    .B(_0807_),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2308_ (.I(_0746_),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2309_ (.I(_0721_),
    .Z(_0810_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2310_ (.I(_0714_),
    .Z(_0811_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2311_ (.A1(_0809_),
    .A2(\mem[7][11] ),
    .B1(\mem[4][11] ),
    .B2(_0810_),
    .C1(_0811_),
    .C2(\mem[6][11] ),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _2312_ (.A1(_0594_),
    .A2(_0723_),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2313_ (.I(_0813_),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2314_ (.I(_0598_),
    .Z(_0815_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2315_ (.A1(\mem[10][11] ),
    .A2(_0814_),
    .B(_0815_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2316_ (.I(_0714_),
    .Z(_0817_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2317_ (.I(_1517_),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2318_ (.I(_0818_),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2319_ (.I(_0721_),
    .Z(_0820_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2320_ (.A1(\mem[14][11] ),
    .A2(_0817_),
    .B1(_0819_),
    .B2(\mem[13][11] ),
    .C1(\mem[12][11] ),
    .C2(_0820_),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2321_ (.A1(_0808_),
    .A2(_0812_),
    .B1(_0816_),
    .B2(_0821_),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2322_ (.A1(_0808_),
    .A2(_0816_),
    .B(_1503_),
    .ZN(_0823_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2323_ (.I(_0729_),
    .Z(_0824_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2324_ (.A1(\rd_ptr_bin[3] ),
    .A2(_1519_),
    .Z(_0825_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2325_ (.I(_0825_),
    .Z(_0826_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2326_ (.I(_1517_),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2327_ (.A1(_0716_),
    .A2(\mem[1][11] ),
    .A3(_0827_),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2328_ (.A1(\mem[11][11] ),
    .A2(_0826_),
    .B(_0828_),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2329_ (.A1(_0729_),
    .A2(\mem[5][11] ),
    .A3(_0747_),
    .Z(_0830_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2330_ (.I(_0594_),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2331_ (.I(_0723_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2332_ (.A1(_0831_),
    .A2(\mem[2][11] ),
    .A3(_0832_),
    .Z(_0833_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2333_ (.A1(_0830_),
    .A2(_0833_),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2334_ (.A1(_0824_),
    .A2(_0829_),
    .B1(_0834_),
    .B2(_0720_),
    .ZN(_0835_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2335_ (.I(_0787_),
    .Z(_0836_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2336_ (.I(_1514_),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2337_ (.I(_0837_),
    .Z(_0838_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2338_ (.I(_0818_),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2339_ (.A1(\mem[8][11] ),
    .A2(_0838_),
    .B1(_0839_),
    .B2(\mem[9][11] ),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2340_ (.A1(_1519_),
    .A2(_0791_),
    .Z(_0841_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2341_ (.I(_0841_),
    .Z(_0842_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2342_ (.I(_0842_),
    .Z(_0843_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2343_ (.A1(\mem[15][11] ),
    .A2(_0843_),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2344_ (.A1(_0836_),
    .A2(_0840_),
    .B(_0844_),
    .C(_0764_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2345_ (.A1(_0822_),
    .A2(_0823_),
    .B(_0835_),
    .C(_0845_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2346_ (.A1(\mem[0][11] ),
    .A2(_0765_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2347_ (.A1(net47),
    .A2(_0762_),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2348_ (.A1(_0768_),
    .A2(_0846_),
    .A3(_0847_),
    .B(_0848_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2349_ (.I(_0825_),
    .Z(_0849_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2350_ (.A1(_0598_),
    .A2(\mem[6][12] ),
    .A3(_0723_),
    .Z(_0850_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2351_ (.A1(\mem[15][12] ),
    .A2(_0849_),
    .B(_0850_),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2352_ (.A1(_0598_),
    .A2(\mem[1][12] ),
    .A3(_0726_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2353_ (.A1(\mem[11][12] ),
    .A2(_0849_),
    .B(_0852_),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2354_ (.I0(_0851_),
    .I1(_0853_),
    .S(_0784_),
    .Z(_0854_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2355_ (.A1(\mem[12][12] ),
    .A2(_0780_),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2356_ (.A1(\mem[9][12] ),
    .A2(_0776_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2357_ (.I(_1517_),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2358_ (.A1(\mem[5][12] ),
    .A2(_0857_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2359_ (.A1(\mem[2][12] ),
    .A2(_0832_),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2360_ (.I0(_0855_),
    .I1(_0856_),
    .I2(_0858_),
    .I3(_0859_),
    .S0(_0784_),
    .S1(_1499_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2361_ (.A1(\mem[13][12] ),
    .A2(_0747_),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2362_ (.A1(\mem[10][12] ),
    .A2(_0832_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2363_ (.A1(\mem[4][12] ),
    .A2(_0837_),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2364_ (.A1(_0746_),
    .A2(\mem[3][12] ),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2365_ (.I(_0594_),
    .Z(_0865_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2366_ (.I0(_0861_),
    .I1(_0862_),
    .I2(_0863_),
    .I3(_0864_),
    .S0(_0865_),
    .S1(_0774_),
    .Z(_0866_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2367_ (.A1(_0754_),
    .A2(_0739_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2368_ (.A1(\rd_ptr_bin[3] ),
    .A2(\mem[14][12] ),
    .A3(_0714_),
    .Z(_0868_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2369_ (.A1(_0597_),
    .A2(_0710_),
    .A3(\mem[7][12] ),
    .Z(_0869_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2370_ (.A1(_0868_),
    .A2(_0869_),
    .Z(_0870_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2371_ (.A1(\mem[8][12] ),
    .A2(_0867_),
    .B1(_0870_),
    .B2(_0734_),
    .C(_0758_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2372_ (.A1(_0854_),
    .A2(_0860_),
    .A3(_0866_),
    .A4(_0871_),
    .Z(_0872_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2373_ (.A1(\mem[0][12] ),
    .A2(_0765_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2374_ (.A1(net48),
    .A2(_0762_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2375_ (.A1(_0768_),
    .A2(_0872_),
    .A3(_0873_),
    .B(_0874_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2376_ (.A1(\mem[3][13] ),
    .A2(_0806_),
    .B(_0807_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2377_ (.I(_0714_),
    .Z(_0876_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2378_ (.A1(_0809_),
    .A2(\mem[7][13] ),
    .B1(\mem[4][13] ),
    .B2(_0810_),
    .C1(_0876_),
    .C2(\mem[6][13] ),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2379_ (.A1(\mem[10][13] ),
    .A2(_0814_),
    .B(_0815_),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2380_ (.A1(\mem[14][13] ),
    .A2(_0817_),
    .B1(_0819_),
    .B2(\mem[13][13] ),
    .C1(\mem[12][13] ),
    .C2(_0820_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2381_ (.A1(_0875_),
    .A2(_0877_),
    .B1(_0878_),
    .B2(_0879_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2382_ (.A1(_0875_),
    .A2(_0878_),
    .B(_1503_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2383_ (.A1(_0716_),
    .A2(\mem[1][13] ),
    .A3(_0827_),
    .Z(_0882_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2384_ (.A1(\mem[11][13] ),
    .A2(_0826_),
    .B(_0882_),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2385_ (.A1(_0729_),
    .A2(\mem[5][13] ),
    .A3(_0747_),
    .Z(_0884_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2386_ (.A1(_0831_),
    .A2(\mem[2][13] ),
    .A3(_0832_),
    .Z(_0885_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2387_ (.A1(_0884_),
    .A2(_0885_),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2388_ (.A1(_0824_),
    .A2(_0883_),
    .B1(_0886_),
    .B2(_0720_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2389_ (.A1(\mem[8][13] ),
    .A2(_0838_),
    .B1(_0839_),
    .B2(\mem[9][13] ),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2390_ (.A1(\mem[15][13] ),
    .A2(_0843_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2391_ (.A1(_0836_),
    .A2(_0888_),
    .B(_0889_),
    .C(_0764_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2392_ (.A1(_0880_),
    .A2(_0881_),
    .B(_0887_),
    .C(_0890_),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2393_ (.A1(\mem[0][13] ),
    .A2(_0765_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2394_ (.A1(net49),
    .A2(_0762_),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2395_ (.A1(_0768_),
    .A2(_0891_),
    .A3(_0892_),
    .B(_0893_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2396_ (.A1(_0598_),
    .A2(\mem[6][14] ),
    .A3(_0723_),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2397_ (.A1(\mem[15][14] ),
    .A2(_0849_),
    .B(_0894_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2398_ (.A1(_0597_),
    .A2(\mem[1][14] ),
    .A3(_0726_),
    .Z(_0896_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2399_ (.A1(\mem[11][14] ),
    .A2(_0849_),
    .B(_0896_),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2400_ (.I0(_0895_),
    .I1(_0897_),
    .S(_0784_),
    .Z(_0898_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2401_ (.A1(\mem[12][14] ),
    .A2(_0780_),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2402_ (.A1(\mem[9][14] ),
    .A2(_0776_),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2403_ (.A1(\mem[5][14] ),
    .A2(_0857_),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2404_ (.A1(\mem[2][14] ),
    .A2(_0832_),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2405_ (.I0(_0899_),
    .I1(_0900_),
    .I2(_0901_),
    .I3(_0902_),
    .S0(_0784_),
    .S1(_1499_),
    .Z(_0903_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2406_ (.A1(\mem[13][14] ),
    .A2(_0747_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2407_ (.A1(\mem[10][14] ),
    .A2(_0832_),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2408_ (.A1(\mem[4][14] ),
    .A2(_0837_),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2409_ (.A1(_0746_),
    .A2(\mem[3][14] ),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2410_ (.I0(_0904_),
    .I1(_0905_),
    .I2(_0906_),
    .I3(_0907_),
    .S0(_0865_),
    .S1(_0774_),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2411_ (.A1(\rd_ptr_bin[3] ),
    .A2(\mem[14][14] ),
    .A3(_0723_),
    .Z(_0909_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2412_ (.A1(_0597_),
    .A2(_0710_),
    .A3(\mem[7][14] ),
    .Z(_0910_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2413_ (.A1(_0909_),
    .A2(_0910_),
    .Z(_0911_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2414_ (.A1(\mem[8][14] ),
    .A2(_0867_),
    .B1(_0911_),
    .B2(_0734_),
    .C(_0758_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2415_ (.A1(_0898_),
    .A2(_0903_),
    .A3(_0908_),
    .A4(_0912_),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2416_ (.A1(\mem[0][14] ),
    .A2(_0765_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2417_ (.A1(net50),
    .A2(_0762_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2418_ (.A1(_0768_),
    .A2(_0913_),
    .A3(_0914_),
    .B(_0915_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2419_ (.I(_0719_),
    .Z(_0916_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2420_ (.A1(\mem[3][15] ),
    .A2(_0806_),
    .B(_0916_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2421_ (.A1(_0809_),
    .A2(\mem[7][15] ),
    .B1(\mem[4][15] ),
    .B2(_0810_),
    .C1(_0876_),
    .C2(\mem[6][15] ),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2422_ (.A1(\mem[10][15] ),
    .A2(_0814_),
    .B(_0815_),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2423_ (.A1(\mem[14][15] ),
    .A2(_0817_),
    .B1(_0819_),
    .B2(\mem[13][15] ),
    .C1(\mem[12][15] ),
    .C2(_0820_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2424_ (.A1(_0917_),
    .A2(_0918_),
    .B1(_0919_),
    .B2(_0920_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2425_ (.A1(_0917_),
    .A2(_0919_),
    .B(_1503_),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2426_ (.A1(_0716_),
    .A2(\mem[1][15] ),
    .A3(_0827_),
    .Z(_0923_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2427_ (.A1(\mem[11][15] ),
    .A2(_0826_),
    .B(_0923_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2428_ (.A1(_0729_),
    .A2(\mem[5][15] ),
    .A3(_0747_),
    .Z(_0925_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2429_ (.A1(_0831_),
    .A2(\mem[2][15] ),
    .A3(_0832_),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2430_ (.A1(_0925_),
    .A2(_0926_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2431_ (.A1(_0824_),
    .A2(_0924_),
    .B1(_0927_),
    .B2(_0720_),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2432_ (.A1(\mem[8][15] ),
    .A2(_0838_),
    .B1(_0839_),
    .B2(\mem[9][15] ),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2433_ (.A1(\mem[15][15] ),
    .A2(_0843_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2434_ (.A1(_0836_),
    .A2(_0929_),
    .B(_0930_),
    .C(_0764_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2435_ (.A1(_0921_),
    .A2(_0922_),
    .B(_0928_),
    .C(_0931_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2436_ (.A1(\mem[0][15] ),
    .A2(_0765_),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2437_ (.A1(net51),
    .A2(_0762_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2438_ (.A1(_0768_),
    .A2(_0932_),
    .A3(_0933_),
    .B(_0934_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2439_ (.I(\mem[7][16] ),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2440_ (.I(\mem[11][16] ),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2441_ (.A1(_0935_),
    .A2(_0738_),
    .B1(_0740_),
    .B2(_0936_),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2442_ (.A1(\mem[2][16] ),
    .A2(_0790_),
    .B1(_0792_),
    .B2(\mem[14][16] ),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2443_ (.I(_0938_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2444_ (.A1(_0744_),
    .A2(_0937_),
    .B1(_0939_),
    .B2(_0795_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2445_ (.A1(_0716_),
    .A2(_0865_),
    .A3(_0727_),
    .Z(_0941_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2446_ (.A1(\mem[8][16] ),
    .A2(_0771_),
    .B1(_0747_),
    .B2(\mem[9][16] ),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2447_ (.A1(_0740_),
    .A2(_0942_),
    .ZN(_0943_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2448_ (.A1(\mem[1][16] ),
    .A2(_0941_),
    .B(_0943_),
    .ZN(_0944_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2449_ (.A1(\mem[6][16] ),
    .A2(_0714_),
    .B1(_0726_),
    .B2(\mem[5][16] ),
    .C1(\mem[4][16] ),
    .C2(_0721_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2450_ (.A1(_0746_),
    .A2(\mem[3][16] ),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2451_ (.A1(_0710_),
    .A2(\mem[15][16] ),
    .B1(\mem[12][16] ),
    .B2(_0721_),
    .C1(_0726_),
    .C2(\mem[13][16] ),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2452_ (.A1(\mem[10][16] ),
    .A2(_0832_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2453_ (.I0(_0945_),
    .I1(_0946_),
    .I2(_0947_),
    .I3(_0948_),
    .S0(_0865_),
    .S1(_0719_),
    .Z(_0949_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2454_ (.A1(_0764_),
    .A2(_0940_),
    .A3(_0944_),
    .A4(_0949_),
    .Z(_0950_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2455_ (.A1(\mem[0][16] ),
    .A2(_0765_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2456_ (.A1(net52),
    .A2(_0762_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2457_ (.A1(_0768_),
    .A2(_0950_),
    .A3(_0951_),
    .B(_0952_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2458_ (.A1(\mem[3][17] ),
    .A2(_0806_),
    .B(_0916_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2459_ (.A1(_0809_),
    .A2(\mem[7][17] ),
    .B1(\mem[4][17] ),
    .B2(_0810_),
    .C1(_0876_),
    .C2(\mem[6][17] ),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2460_ (.A1(\mem[10][17] ),
    .A2(_0814_),
    .B(_0815_),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2461_ (.A1(\mem[14][17] ),
    .A2(_0817_),
    .B1(_0819_),
    .B2(\mem[13][17] ),
    .C1(\mem[12][17] ),
    .C2(_0820_),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2462_ (.A1(_0953_),
    .A2(_0954_),
    .B1(_0955_),
    .B2(_0956_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2463_ (.A1(_0953_),
    .A2(_0955_),
    .B(_1503_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2464_ (.I(_0597_),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2465_ (.A1(_0959_),
    .A2(\mem[1][17] ),
    .A3(_0827_),
    .Z(_0960_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2466_ (.A1(\mem[11][17] ),
    .A2(_0826_),
    .B(_0960_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2467_ (.A1(_0729_),
    .A2(\mem[5][17] ),
    .A3(_0747_),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2468_ (.I(_0723_),
    .Z(_0963_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2469_ (.A1(_0831_),
    .A2(\mem[2][17] ),
    .A3(_0963_),
    .Z(_0964_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2470_ (.A1(_0962_),
    .A2(_0964_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2471_ (.A1(_0824_),
    .A2(_0961_),
    .B1(_0965_),
    .B2(_0720_),
    .ZN(_0966_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2472_ (.A1(\mem[8][17] ),
    .A2(_0838_),
    .B1(_0839_),
    .B2(\mem[9][17] ),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2473_ (.A1(\mem[15][17] ),
    .A2(_0843_),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2474_ (.I(_0763_),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2475_ (.A1(_0836_),
    .A2(_0967_),
    .B(_0968_),
    .C(_0969_),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2476_ (.A1(_0957_),
    .A2(_0958_),
    .B(_0966_),
    .C(_0970_),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2477_ (.A1(\mem[0][17] ),
    .A2(_0765_),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2478_ (.I(_0761_),
    .Z(_0973_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2479_ (.A1(net53),
    .A2(_0973_),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2480_ (.A1(_0768_),
    .A2(_0971_),
    .A3(_0972_),
    .B(_0974_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2481_ (.A1(_0743_),
    .A2(\mem[15][18] ),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2482_ (.A1(\mem[6][18] ),
    .A2(_0731_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2483_ (.A1(\mem[8][18] ),
    .A2(_0771_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2484_ (.A1(\mem[1][18] ),
    .A2(_0727_),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2485_ (.I0(_0975_),
    .I1(_0976_),
    .I2(_0977_),
    .I3(_0978_),
    .S0(_0774_),
    .S1(_0709_),
    .Z(_0979_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2486_ (.A1(\mem[13][18] ),
    .A2(_0776_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2487_ (.A1(\mem[10][18] ),
    .A2(_0778_),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2488_ (.A1(\mem[4][18] ),
    .A2(_0780_),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2489_ (.A1(_0782_),
    .A2(\mem[3][18] ),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2490_ (.I0(_0980_),
    .I1(_0981_),
    .I2(_0982_),
    .I3(_0983_),
    .S0(_0784_),
    .S1(_1499_),
    .Z(_0984_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2491_ (.I(\mem[7][18] ),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2492_ (.I(\mem[11][18] ),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2493_ (.A1(_0985_),
    .A2(_0738_),
    .B1(_0787_),
    .B2(_0986_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2494_ (.A1(\mem[2][18] ),
    .A2(_0790_),
    .B1(_0792_),
    .B2(\mem[14][18] ),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2495_ (.I(_0988_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2496_ (.A1(_0744_),
    .A2(_0987_),
    .B1(_0989_),
    .B2(_0795_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2497_ (.A1(_0733_),
    .A2(\mem[12][18] ),
    .A3(_0721_),
    .Z(_0991_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2498_ (.I(_0594_),
    .Z(_0992_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2499_ (.A1(_0992_),
    .A2(\mem[9][18] ),
    .A3(_0726_),
    .Z(_0993_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2500_ (.A1(_0991_),
    .A2(_0993_),
    .Z(_0994_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2501_ (.A1(\mem[5][18] ),
    .A2(_0753_),
    .B1(_0994_),
    .B2(_0800_),
    .C(_0758_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2502_ (.A1(_0979_),
    .A2(_0984_),
    .A3(_0990_),
    .A4(_0995_),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2503_ (.A1(\mem[0][18] ),
    .A2(_0765_),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2504_ (.A1(net54),
    .A2(_0973_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2505_ (.A1(_0768_),
    .A2(_0996_),
    .A3(_0997_),
    .B(_0998_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2506_ (.A1(\mem[3][19] ),
    .A2(_0806_),
    .B(_0916_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2507_ (.I(_0837_),
    .Z(_1000_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2508_ (.A1(_0809_),
    .A2(\mem[7][19] ),
    .B1(\mem[4][19] ),
    .B2(_1000_),
    .C1(_0876_),
    .C2(\mem[6][19] ),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2509_ (.I(_0598_),
    .Z(_1002_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2510_ (.A1(\mem[10][19] ),
    .A2(_0814_),
    .B(_1002_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2511_ (.I(_0818_),
    .Z(_1004_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2512_ (.A1(\mem[14][19] ),
    .A2(_0817_),
    .B1(_1004_),
    .B2(\mem[13][19] ),
    .C1(\mem[12][19] ),
    .C2(_0820_),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2513_ (.A1(_0999_),
    .A2(_1001_),
    .B1(_1003_),
    .B2(_1005_),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2514_ (.A1(_0999_),
    .A2(_1003_),
    .B(_1503_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2515_ (.A1(_0959_),
    .A2(\mem[1][19] ),
    .A3(_0827_),
    .Z(_1008_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2516_ (.A1(\mem[11][19] ),
    .A2(_0826_),
    .B(_1008_),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2517_ (.A1(_0729_),
    .A2(\mem[5][19] ),
    .A3(_0747_),
    .Z(_1010_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2518_ (.A1(_0831_),
    .A2(\mem[2][19] ),
    .A3(_0963_),
    .Z(_1011_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2519_ (.A1(_1010_),
    .A2(_1011_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2520_ (.A1(_0824_),
    .A2(_1009_),
    .B1(_1012_),
    .B2(_0720_),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2521_ (.A1(\mem[8][19] ),
    .A2(_0838_),
    .B1(_0839_),
    .B2(\mem[9][19] ),
    .ZN(_1014_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2522_ (.A1(\mem[15][19] ),
    .A2(_0843_),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2523_ (.A1(_0836_),
    .A2(_1014_),
    .B(_1015_),
    .C(_0969_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2524_ (.A1(_1006_),
    .A2(_1007_),
    .B(_1013_),
    .C(_1016_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2525_ (.I(_0764_),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2526_ (.A1(\mem[0][19] ),
    .A2(_1018_),
    .ZN(_1019_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2527_ (.A1(net55),
    .A2(_0973_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2528_ (.A1(_0768_),
    .A2(_1017_),
    .A3(_1019_),
    .B(_1020_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 _2529_ (.I(_0761_),
    .Z(_1021_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2530_ (.A1(\mem[3][1] ),
    .A2(_0806_),
    .B(_0916_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 _2531_ (.I(_0710_),
    .Z(_1023_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2532_ (.A1(_1023_),
    .A2(\mem[7][1] ),
    .B1(\mem[4][1] ),
    .B2(_1000_),
    .C1(_0876_),
    .C2(\mem[6][1] ),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2533_ (.A1(\mem[10][1] ),
    .A2(_0814_),
    .B(_1002_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2534_ (.A1(\mem[14][1] ),
    .A2(_0817_),
    .B1(_1004_),
    .B2(\mem[13][1] ),
    .C1(\mem[12][1] ),
    .C2(_0820_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2535_ (.A1(_1022_),
    .A2(_1024_),
    .B1(_1025_),
    .B2(_1026_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2536_ (.A1(_1022_),
    .A2(_1025_),
    .B(_1503_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2537_ (.A1(_0959_),
    .A2(\mem[1][1] ),
    .A3(_0827_),
    .Z(_1029_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2538_ (.A1(\mem[11][1] ),
    .A2(_0826_),
    .B(_1029_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2539_ (.I(_1517_),
    .Z(_1031_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2540_ (.A1(_0729_),
    .A2(\mem[5][1] ),
    .A3(_1031_),
    .Z(_1032_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2541_ (.A1(_0831_),
    .A2(\mem[2][1] ),
    .A3(_0963_),
    .Z(_1033_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2542_ (.A1(_1032_),
    .A2(_1033_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2543_ (.A1(_0824_),
    .A2(_1030_),
    .B1(_1034_),
    .B2(_0720_),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2544_ (.A1(\mem[8][1] ),
    .A2(_0838_),
    .B1(_0839_),
    .B2(\mem[9][1] ),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2545_ (.A1(\mem[15][1] ),
    .A2(_0843_),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2546_ (.A1(_0836_),
    .A2(_1036_),
    .B(_1037_),
    .C(_0969_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2547_ (.A1(_1027_),
    .A2(_1028_),
    .B(_1035_),
    .C(_1038_),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2548_ (.A1(\mem[0][1] ),
    .A2(_1018_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2549_ (.A1(net56),
    .A2(_0973_),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2550_ (.A1(_1021_),
    .A2(_1039_),
    .A3(_1040_),
    .B(_1041_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2551_ (.A1(_0743_),
    .A2(\mem[15][20] ),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2552_ (.A1(\mem[6][20] ),
    .A2(_0731_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2553_ (.A1(\mem[8][20] ),
    .A2(_0771_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2554_ (.A1(\mem[1][20] ),
    .A2(_0727_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2555_ (.I0(_1042_),
    .I1(_1043_),
    .I2(_1044_),
    .I3(_1045_),
    .S0(_0774_),
    .S1(_0596_),
    .Z(_1046_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2556_ (.A1(\mem[13][20] ),
    .A2(_0776_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2557_ (.A1(\mem[10][20] ),
    .A2(_0778_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2558_ (.A1(\mem[4][20] ),
    .A2(_0780_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2559_ (.A1(_0782_),
    .A2(\mem[3][20] ),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2560_ (.I0(_1047_),
    .I1(_1048_),
    .I2(_1049_),
    .I3(_1050_),
    .S0(_0784_),
    .S1(_1499_),
    .Z(_1051_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2561_ (.I(\mem[7][20] ),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2562_ (.I(\mem[11][20] ),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2563_ (.A1(_1052_),
    .A2(_0738_),
    .B1(_0787_),
    .B2(_1053_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2564_ (.A1(\mem[2][20] ),
    .A2(_0790_),
    .B1(_0792_),
    .B2(\mem[14][20] ),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2565_ (.I(_1055_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2566_ (.A1(_0744_),
    .A2(_1054_),
    .B1(_1056_),
    .B2(_0795_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2567_ (.A1(_0733_),
    .A2(\mem[12][20] ),
    .A3(_0721_),
    .Z(_1058_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2568_ (.A1(_0992_),
    .A2(\mem[9][20] ),
    .A3(_0726_),
    .Z(_1059_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2569_ (.A1(_1058_),
    .A2(_1059_),
    .Z(_1060_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2570_ (.A1(\mem[5][20] ),
    .A2(_0753_),
    .B1(_1060_),
    .B2(_0800_),
    .C(_0758_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2571_ (.A1(_1046_),
    .A2(_1051_),
    .A3(_1057_),
    .A4(_1061_),
    .Z(_1062_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2572_ (.A1(\mem[0][20] ),
    .A2(_1018_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2573_ (.A1(net57),
    .A2(_0973_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2574_ (.A1(_1021_),
    .A2(_1062_),
    .A3(_1063_),
    .B(_1064_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2575_ (.A1(\mem[3][21] ),
    .A2(_0806_),
    .B(_0916_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_4 _2576_ (.A1(_1023_),
    .A2(\mem[7][21] ),
    .B1(\mem[4][21] ),
    .B2(_1000_),
    .C1(_0876_),
    .C2(\mem[6][21] ),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2577_ (.A1(\mem[10][21] ),
    .A2(_0814_),
    .B(_1002_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2578_ (.A1(\mem[14][21] ),
    .A2(_0817_),
    .B1(_1004_),
    .B2(\mem[13][21] ),
    .C1(\mem[12][21] ),
    .C2(_0820_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2579_ (.A1(_1065_),
    .A2(_1066_),
    .B1(_1067_),
    .B2(_1068_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2580_ (.A1(_1065_),
    .A2(_1067_),
    .B(_1503_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2581_ (.A1(_0959_),
    .A2(\mem[1][21] ),
    .A3(_0827_),
    .Z(_1071_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2582_ (.A1(\mem[11][21] ),
    .A2(_0826_),
    .B(_1071_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _2583_ (.I(_0728_),
    .Z(_1073_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2584_ (.A1(_1073_),
    .A2(\mem[5][21] ),
    .A3(_1031_),
    .Z(_1074_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2585_ (.A1(_0831_),
    .A2(\mem[2][21] ),
    .A3(_0963_),
    .Z(_1075_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2586_ (.A1(_1074_),
    .A2(_1075_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2587_ (.A1(_0824_),
    .A2(_1072_),
    .B1(_1076_),
    .B2(_0720_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2588_ (.A1(\mem[8][21] ),
    .A2(_0838_),
    .B1(_0839_),
    .B2(\mem[9][21] ),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2589_ (.A1(\mem[15][21] ),
    .A2(_0843_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2590_ (.A1(_0836_),
    .A2(_1078_),
    .B(_1079_),
    .C(_0969_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2591_ (.A1(_1069_),
    .A2(_1070_),
    .B(_1077_),
    .C(_1080_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2592_ (.A1(\mem[0][21] ),
    .A2(_1018_),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2593_ (.A1(net58),
    .A2(_0973_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2594_ (.A1(_1021_),
    .A2(_1081_),
    .A3(_1082_),
    .B(_1083_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2595_ (.A1(_0743_),
    .A2(\mem[15][22] ),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2596_ (.A1(\mem[6][22] ),
    .A2(_0724_),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2597_ (.A1(\mem[8][22] ),
    .A2(_0771_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2598_ (.A1(\mem[1][22] ),
    .A2(_0727_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2599_ (.I0(_1084_),
    .I1(_1085_),
    .I2(_1086_),
    .I3(_1087_),
    .S0(_0774_),
    .S1(_0596_),
    .Z(_1088_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2600_ (.A1(\mem[13][22] ),
    .A2(_0857_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2601_ (.A1(\mem[10][22] ),
    .A2(_0778_),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2602_ (.A1(\mem[4][22] ),
    .A2(_0780_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2603_ (.A1(_0782_),
    .A2(\mem[3][22] ),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2604_ (.I0(_1089_),
    .I1(_1090_),
    .I2(_1091_),
    .I3(_1092_),
    .S0(_0784_),
    .S1(_1499_),
    .Z(_1093_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2605_ (.I(\mem[7][22] ),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2606_ (.I(\mem[11][22] ),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2607_ (.A1(_1094_),
    .A2(_0738_),
    .B1(_0787_),
    .B2(_1095_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2608_ (.A1(\mem[2][22] ),
    .A2(_0790_),
    .B1(_0792_),
    .B2(\mem[14][22] ),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2609_ (.I(_1097_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2610_ (.A1(_0744_),
    .A2(_1096_),
    .B1(_1098_),
    .B2(_0795_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2611_ (.A1(_0733_),
    .A2(\mem[12][22] ),
    .A3(_0711_),
    .Z(_1100_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2612_ (.A1(_0992_),
    .A2(\mem[9][22] ),
    .A3(_0712_),
    .Z(_1101_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2613_ (.A1(_1100_),
    .A2(_1101_),
    .Z(_1102_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2614_ (.A1(\mem[5][22] ),
    .A2(_0753_),
    .B1(_1102_),
    .B2(_0807_),
    .C(_0758_),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2615_ (.A1(_1088_),
    .A2(_1093_),
    .A3(_1099_),
    .A4(_1103_),
    .Z(_1104_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2616_ (.A1(\mem[0][22] ),
    .A2(_1018_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2617_ (.A1(net59),
    .A2(_0973_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2618_ (.A1(_1021_),
    .A2(_1104_),
    .A3(_1105_),
    .B(_1106_),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2619_ (.A1(\mem[3][23] ),
    .A2(_0806_),
    .B(_0916_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2620_ (.A1(_1023_),
    .A2(\mem[7][23] ),
    .B1(\mem[4][23] ),
    .B2(_1000_),
    .C1(_0876_),
    .C2(\mem[6][23] ),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2621_ (.A1(\mem[10][23] ),
    .A2(_0814_),
    .B(_1002_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2622_ (.A1(\mem[14][23] ),
    .A2(_0811_),
    .B1(_1004_),
    .B2(\mem[13][23] ),
    .C1(\mem[12][23] ),
    .C2(_0820_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2623_ (.A1(_1107_),
    .A2(_1108_),
    .B1(_1109_),
    .B2(_1110_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2624_ (.A1(_1107_),
    .A2(_1109_),
    .B(_1503_),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2625_ (.A1(_0959_),
    .A2(\mem[1][23] ),
    .A3(_0827_),
    .Z(_1113_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2626_ (.A1(\mem[11][23] ),
    .A2(_0826_),
    .B(_1113_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2627_ (.A1(_1073_),
    .A2(\mem[5][23] ),
    .A3(_1031_),
    .Z(_1115_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2628_ (.A1(_0831_),
    .A2(\mem[2][23] ),
    .A3(_0963_),
    .Z(_1116_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2629_ (.A1(_1115_),
    .A2(_1116_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2630_ (.A1(_0824_),
    .A2(_1114_),
    .B1(_1117_),
    .B2(_0720_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2631_ (.A1(\mem[8][23] ),
    .A2(_0838_),
    .B1(_0839_),
    .B2(\mem[9][23] ),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2632_ (.A1(\mem[15][23] ),
    .A2(_0843_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2633_ (.A1(_0836_),
    .A2(_1119_),
    .B(_1120_),
    .C(_0969_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2634_ (.A1(_1111_),
    .A2(_1112_),
    .B(_1118_),
    .C(_1121_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2635_ (.A1(\mem[0][23] ),
    .A2(_1018_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2636_ (.A1(net60),
    .A2(_0973_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2637_ (.A1(_1021_),
    .A2(_1122_),
    .A3(_1123_),
    .B(_1124_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2638_ (.A1(_0743_),
    .A2(\mem[15][24] ),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2639_ (.A1(\mem[6][24] ),
    .A2(_0724_),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2640_ (.A1(\mem[8][24] ),
    .A2(_0771_),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2641_ (.A1(\mem[1][24] ),
    .A2(_0727_),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2642_ (.I0(_1125_),
    .I1(_1126_),
    .I2(_1127_),
    .I3(_1128_),
    .S0(_0774_),
    .S1(_0596_),
    .Z(_1129_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2643_ (.A1(\mem[13][24] ),
    .A2(_0857_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2644_ (.A1(\mem[10][24] ),
    .A2(_0778_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2645_ (.A1(\mem[4][24] ),
    .A2(_0780_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2646_ (.A1(_0782_),
    .A2(\mem[3][24] ),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2647_ (.I0(_1130_),
    .I1(_1131_),
    .I2(_1132_),
    .I3(_1133_),
    .S0(_0784_),
    .S1(_1499_),
    .Z(_1134_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2648_ (.I(\mem[7][24] ),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2649_ (.I(\mem[11][24] ),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2650_ (.A1(_1135_),
    .A2(_0738_),
    .B1(_0787_),
    .B2(_1136_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2651_ (.A1(\mem[2][24] ),
    .A2(_0790_),
    .B1(_0792_),
    .B2(\mem[14][24] ),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2652_ (.I(_1138_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2653_ (.A1(_0744_),
    .A2(_1137_),
    .B1(_1139_),
    .B2(_0795_),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2654_ (.A1(_0733_),
    .A2(\mem[12][24] ),
    .A3(_0711_),
    .Z(_1141_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2655_ (.A1(_0992_),
    .A2(\mem[9][24] ),
    .A3(_0712_),
    .Z(_1142_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2656_ (.A1(_1141_),
    .A2(_1142_),
    .Z(_1143_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2657_ (.A1(\mem[5][24] ),
    .A2(_0753_),
    .B1(_1143_),
    .B2(_0807_),
    .C(_0758_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2658_ (.A1(_1129_),
    .A2(_1134_),
    .A3(_1140_),
    .A4(_1144_),
    .Z(_1145_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2659_ (.A1(\mem[0][24] ),
    .A2(_1018_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2660_ (.A1(net61),
    .A2(_0973_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2661_ (.A1(_1021_),
    .A2(_1145_),
    .A3(_1146_),
    .B(_1147_),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2662_ (.A1(\mem[3][25] ),
    .A2(_0806_),
    .B(_0916_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2663_ (.A1(_1023_),
    .A2(\mem[7][25] ),
    .B1(\mem[4][25] ),
    .B2(_1000_),
    .C1(_0876_),
    .C2(\mem[6][25] ),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2664_ (.A1(\mem[10][25] ),
    .A2(_0814_),
    .B(_1002_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2665_ (.A1(\mem[14][25] ),
    .A2(_0811_),
    .B1(_1004_),
    .B2(\mem[13][25] ),
    .C1(\mem[12][25] ),
    .C2(_0722_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2666_ (.A1(_1148_),
    .A2(_1149_),
    .B1(_1150_),
    .B2(_1151_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2667_ (.A1(_1148_),
    .A2(_1150_),
    .B(_1503_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2668_ (.A1(_0959_),
    .A2(\mem[1][25] ),
    .A3(_0827_),
    .Z(_1154_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2669_ (.A1(\mem[11][25] ),
    .A2(_0826_),
    .B(_1154_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2670_ (.A1(_1073_),
    .A2(\mem[5][25] ),
    .A3(_1031_),
    .Z(_1156_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2671_ (.A1(_0831_),
    .A2(\mem[2][25] ),
    .A3(_0963_),
    .Z(_1157_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2672_ (.A1(_1156_),
    .A2(_1157_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2673_ (.A1(_0824_),
    .A2(_1155_),
    .B1(_1158_),
    .B2(_0720_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2674_ (.A1(\mem[8][25] ),
    .A2(_0838_),
    .B1(_0839_),
    .B2(\mem[9][25] ),
    .ZN(_1160_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2675_ (.A1(\mem[15][25] ),
    .A2(_0843_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2676_ (.A1(_0836_),
    .A2(_1160_),
    .B(_1161_),
    .C(_0969_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2677_ (.A1(_1152_),
    .A2(_1153_),
    .B(_1159_),
    .C(_1162_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2678_ (.A1(\mem[0][25] ),
    .A2(_1018_),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2679_ (.A1(net62),
    .A2(_0973_),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2680_ (.A1(_1021_),
    .A2(_1163_),
    .A3(_1164_),
    .B(_1165_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2681_ (.A1(_0743_),
    .A2(\mem[15][26] ),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2682_ (.A1(\mem[6][26] ),
    .A2(_0724_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2683_ (.A1(\mem[8][26] ),
    .A2(_0771_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2684_ (.A1(\mem[1][26] ),
    .A2(_0727_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2685_ (.I0(_1166_),
    .I1(_1167_),
    .I2(_1168_),
    .I3(_1169_),
    .S0(_0774_),
    .S1(_0596_),
    .Z(_1170_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2686_ (.A1(\mem[13][26] ),
    .A2(_0857_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2687_ (.A1(\mem[10][26] ),
    .A2(_0778_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2688_ (.A1(\mem[4][26] ),
    .A2(_0837_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2689_ (.A1(_0782_),
    .A2(\mem[3][26] ),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2690_ (.I0(_1171_),
    .I1(_1172_),
    .I2(_1173_),
    .I3(_1174_),
    .S0(_0784_),
    .S1(_0815_),
    .Z(_1175_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2691_ (.I(\mem[7][26] ),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2692_ (.I(\mem[11][26] ),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2693_ (.A1(_1176_),
    .A2(_0738_),
    .B1(_0787_),
    .B2(_1177_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2694_ (.A1(\mem[2][26] ),
    .A2(_0790_),
    .B1(_0792_),
    .B2(\mem[14][26] ),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2695_ (.I(_1179_),
    .ZN(_1180_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2696_ (.A1(_0744_),
    .A2(_1178_),
    .B1(_1180_),
    .B2(_0795_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2697_ (.A1(_0733_),
    .A2(\mem[12][26] ),
    .A3(_0711_),
    .Z(_1182_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2698_ (.A1(_0992_),
    .A2(\mem[9][26] ),
    .A3(_0712_),
    .Z(_1183_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2699_ (.A1(_1182_),
    .A2(_1183_),
    .Z(_1184_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2700_ (.A1(\mem[5][26] ),
    .A2(_0753_),
    .B1(_1184_),
    .B2(_0807_),
    .C(_0758_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2701_ (.A1(_1170_),
    .A2(_1175_),
    .A3(_1181_),
    .A4(_1185_),
    .Z(_1186_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2702_ (.A1(\mem[0][26] ),
    .A2(_1018_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2703_ (.I(_0761_),
    .Z(_1188_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2704_ (.A1(net63),
    .A2(_1188_),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2705_ (.A1(_1021_),
    .A2(_1186_),
    .A3(_1187_),
    .B(_1189_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2706_ (.A1(\mem[3][27] ),
    .A2(_0806_),
    .B(_0916_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2707_ (.A1(_1023_),
    .A2(\mem[7][27] ),
    .B1(\mem[4][27] ),
    .B2(_1000_),
    .C1(_0876_),
    .C2(\mem[6][27] ),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2708_ (.A1(\mem[10][27] ),
    .A2(_0814_),
    .B(_1002_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2709_ (.A1(\mem[14][27] ),
    .A2(_0811_),
    .B1(_1004_),
    .B2(\mem[13][27] ),
    .C1(\mem[12][27] ),
    .C2(_0722_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2710_ (.A1(_1190_),
    .A2(_1191_),
    .B1(_1192_),
    .B2(_1193_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2711_ (.A1(_1190_),
    .A2(_1192_),
    .B(_0709_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2712_ (.A1(_0959_),
    .A2(\mem[1][27] ),
    .A3(_0818_),
    .Z(_1196_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2713_ (.A1(\mem[11][27] ),
    .A2(_0826_),
    .B(_1196_),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2714_ (.A1(_1073_),
    .A2(\mem[5][27] ),
    .A3(_1031_),
    .Z(_1198_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2715_ (.A1(_0831_),
    .A2(\mem[2][27] ),
    .A3(_0963_),
    .Z(_1199_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2716_ (.A1(_1198_),
    .A2(_1199_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2717_ (.A1(_0734_),
    .A2(_1197_),
    .B1(_1200_),
    .B2(_0800_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2718_ (.A1(\mem[8][27] ),
    .A2(_0838_),
    .B1(_0839_),
    .B2(\mem[9][27] ),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2719_ (.A1(\mem[15][27] ),
    .A2(_0842_),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2720_ (.A1(_0836_),
    .A2(_1202_),
    .B(_1203_),
    .C(_0969_),
    .ZN(_1204_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2721_ (.A1(_1194_),
    .A2(_1195_),
    .B(_1201_),
    .C(_1204_),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2722_ (.A1(\mem[0][27] ),
    .A2(_1018_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2723_ (.A1(net64),
    .A2(_1188_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2724_ (.A1(_1021_),
    .A2(_1205_),
    .A3(_1206_),
    .B(_1207_),
    .ZN(_0535_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2725_ (.A1(_0743_),
    .A2(\mem[15][28] ),
    .ZN(_1208_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2726_ (.A1(\mem[6][28] ),
    .A2(_0724_),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2727_ (.A1(\mem[8][28] ),
    .A2(_0771_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2728_ (.A1(\mem[1][28] ),
    .A2(_0776_),
    .ZN(_1211_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2729_ (.I0(_1208_),
    .I1(_1209_),
    .I2(_1210_),
    .I3(_1211_),
    .S0(_0716_),
    .S1(_0596_),
    .Z(_1212_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2730_ (.A1(\mem[13][28] ),
    .A2(_0857_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2731_ (.A1(\mem[10][28] ),
    .A2(_0778_),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2732_ (.A1(\mem[4][28] ),
    .A2(_0837_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2733_ (.A1(_0782_),
    .A2(\mem[3][28] ),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2734_ (.I0(_1213_),
    .I1(_1214_),
    .I2(_1215_),
    .I3(_1216_),
    .S0(_0865_),
    .S1(_0815_),
    .Z(_1217_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2735_ (.I(\mem[7][28] ),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2736_ (.I(\mem[11][28] ),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2737_ (.A1(_1218_),
    .A2(_0738_),
    .B1(_0787_),
    .B2(_1219_),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2738_ (.A1(\mem[2][28] ),
    .A2(_0790_),
    .B1(_0792_),
    .B2(\mem[14][28] ),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2739_ (.I(_1221_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2740_ (.A1(_0744_),
    .A2(_1220_),
    .B1(_1222_),
    .B2(_0795_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2741_ (.A1(_0733_),
    .A2(\mem[12][28] ),
    .A3(_0711_),
    .Z(_1224_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2742_ (.A1(_0992_),
    .A2(\mem[9][28] ),
    .A3(_0712_),
    .Z(_1225_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2743_ (.A1(_1224_),
    .A2(_1225_),
    .Z(_1226_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2744_ (.A1(\mem[5][28] ),
    .A2(_0753_),
    .B1(_1226_),
    .B2(_0807_),
    .C(_0758_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2745_ (.A1(_1212_),
    .A2(_1217_),
    .A3(_1223_),
    .A4(_1227_),
    .Z(_1228_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2746_ (.I(_0764_),
    .Z(_1229_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2747_ (.A1(\mem[0][28] ),
    .A2(_1229_),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2748_ (.A1(net65),
    .A2(_1188_),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2749_ (.A1(_1021_),
    .A2(_1228_),
    .A3(_1230_),
    .B(_1231_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 _2750_ (.I(_0761_),
    .Z(_1232_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2751_ (.A1(\mem[3][29] ),
    .A2(_0805_),
    .B(_0916_),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_4 _2752_ (.A1(_1023_),
    .A2(\mem[7][29] ),
    .B1(\mem[4][29] ),
    .B2(_1000_),
    .C1(_0876_),
    .C2(\mem[6][29] ),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2753_ (.A1(\mem[10][29] ),
    .A2(_0813_),
    .B(_1002_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_4 _2754_ (.A1(\mem[14][29] ),
    .A2(_0811_),
    .B1(_1004_),
    .B2(\mem[13][29] ),
    .C1(\mem[12][29] ),
    .C2(_0722_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2755_ (.A1(_1233_),
    .A2(_1234_),
    .B1(_1235_),
    .B2(_1236_),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2756_ (.A1(_1233_),
    .A2(_1235_),
    .B(_0709_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2757_ (.A1(_0959_),
    .A2(\mem[1][29] ),
    .A3(_0818_),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2758_ (.A1(\mem[11][29] ),
    .A2(_0849_),
    .B(_1239_),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2759_ (.A1(_1073_),
    .A2(\mem[5][29] ),
    .A3(_1031_),
    .Z(_1241_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2760_ (.A1(_0595_),
    .A2(\mem[2][29] ),
    .A3(_0963_),
    .Z(_1242_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2761_ (.A1(_1241_),
    .A2(_1242_),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2762_ (.A1(_0734_),
    .A2(_1240_),
    .B1(_1243_),
    .B2(_0800_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2763_ (.A1(\mem[8][29] ),
    .A2(_0810_),
    .B1(_0819_),
    .B2(\mem[9][29] ),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2764_ (.A1(\mem[15][29] ),
    .A2(_0842_),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2765_ (.A1(_0740_),
    .A2(_1245_),
    .B(_1246_),
    .C(_0969_),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _2766_ (.A1(_1237_),
    .A2(_1238_),
    .B(_1244_),
    .C(_1247_),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2767_ (.A1(\mem[0][29] ),
    .A2(_1229_),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2768_ (.A1(net66),
    .A2(_1188_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2769_ (.A1(_1232_),
    .A2(_1248_),
    .A3(_1249_),
    .B(_1250_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2770_ (.A1(_0743_),
    .A2(\mem[15][2] ),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2771_ (.A1(\mem[6][2] ),
    .A2(_0724_),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2772_ (.A1(\mem[8][2] ),
    .A2(_0771_),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2773_ (.A1(\mem[1][2] ),
    .A2(_0776_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2774_ (.I0(_1251_),
    .I1(_1252_),
    .I2(_1253_),
    .I3(_1254_),
    .S0(_0716_),
    .S1(_0596_),
    .Z(_1255_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2775_ (.A1(\mem[13][2] ),
    .A2(_0857_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2776_ (.A1(\mem[10][2] ),
    .A2(_0778_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2777_ (.A1(\mem[4][2] ),
    .A2(_0837_),
    .ZN(_1258_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2778_ (.A1(_0746_),
    .A2(\mem[3][2] ),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2779_ (.I0(_1256_),
    .I1(_1257_),
    .I2(_1258_),
    .I3(_1259_),
    .S0(_0865_),
    .S1(_0815_),
    .Z(_1260_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2780_ (.I(\mem[7][2] ),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2781_ (.I(\mem[11][2] ),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2782_ (.A1(_1261_),
    .A2(_0737_),
    .B1(_0787_),
    .B2(_1262_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2783_ (.A1(\mem[2][2] ),
    .A2(_0790_),
    .B1(_0792_),
    .B2(\mem[14][2] ),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2784_ (.I(_1264_),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2785_ (.A1(_0809_),
    .A2(_1263_),
    .B1(_1265_),
    .B2(_0795_),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2786_ (.A1(_0733_),
    .A2(\mem[12][2] ),
    .A3(_0711_),
    .Z(_1267_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2787_ (.A1(_0992_),
    .A2(\mem[9][2] ),
    .A3(_0712_),
    .Z(_1268_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2788_ (.A1(_1267_),
    .A2(_1268_),
    .Z(_1269_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2789_ (.A1(\mem[5][2] ),
    .A2(_0753_),
    .B1(_1269_),
    .B2(_0807_),
    .C(_0757_),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2790_ (.A1(_1255_),
    .A2(_1260_),
    .A3(_1266_),
    .A4(_1270_),
    .Z(_1271_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2791_ (.A1(\mem[0][2] ),
    .A2(_1229_),
    .ZN(_1272_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2792_ (.A1(net67),
    .A2(_1188_),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2793_ (.A1(_1232_),
    .A2(_1271_),
    .A3(_1272_),
    .B(_1273_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2794_ (.I(\mem[7][30] ),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2795_ (.I(\mem[11][30] ),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2796_ (.A1(_1274_),
    .A2(_0738_),
    .B1(_0787_),
    .B2(_1275_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2797_ (.A1(\mem[2][30] ),
    .A2(_0790_),
    .B1(_0792_),
    .B2(\mem[14][30] ),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2798_ (.I(_1277_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2799_ (.A1(_0744_),
    .A2(_1276_),
    .B1(_1278_),
    .B2(_0795_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2800_ (.A1(\mem[8][30] ),
    .A2(_0771_),
    .B1(_0747_),
    .B2(\mem[9][30] ),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2801_ (.A1(_0740_),
    .A2(_1280_),
    .ZN(_1281_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2802_ (.A1(\mem[1][30] ),
    .A2(_0941_),
    .B(_1281_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2803_ (.A1(\mem[6][30] ),
    .A2(_0714_),
    .B1(_0726_),
    .B2(\mem[5][30] ),
    .C1(\mem[4][30] ),
    .C2(_0721_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2804_ (.A1(_0746_),
    .A2(\mem[3][30] ),
    .ZN(_1284_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2805_ (.A1(_0710_),
    .A2(\mem[15][30] ),
    .B1(\mem[12][30] ),
    .B2(_0721_),
    .C1(_0726_),
    .C2(\mem[13][30] ),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2806_ (.A1(\mem[10][30] ),
    .A2(_0832_),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2807_ (.I0(_1283_),
    .I1(_1284_),
    .I2(_1285_),
    .I3(_1286_),
    .S0(_0865_),
    .S1(_0719_),
    .Z(_1287_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2808_ (.A1(_0764_),
    .A2(_1279_),
    .A3(_1282_),
    .A4(_1287_),
    .Z(_1288_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2809_ (.A1(\mem[0][30] ),
    .A2(_1229_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2810_ (.A1(net68),
    .A2(_1188_),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2811_ (.A1(_1232_),
    .A2(_1288_),
    .A3(_1289_),
    .B(_1290_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2812_ (.A1(\mem[3][31] ),
    .A2(_0805_),
    .B(_0916_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2813_ (.A1(_1023_),
    .A2(\mem[7][31] ),
    .B1(\mem[4][31] ),
    .B2(_1000_),
    .C1(_0731_),
    .C2(\mem[6][31] ),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2814_ (.A1(\mem[10][31] ),
    .A2(_0813_),
    .B(_1002_),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2815_ (.A1(\mem[14][31] ),
    .A2(_0811_),
    .B1(_1004_),
    .B2(\mem[13][31] ),
    .C1(\mem[12][31] ),
    .C2(_0722_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2816_ (.A1(_1291_),
    .A2(_1292_),
    .B1(_1293_),
    .B2(_1294_),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2817_ (.A1(_1291_),
    .A2(_1293_),
    .B(_0709_),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2818_ (.A1(_0959_),
    .A2(\mem[1][31] ),
    .A3(_0818_),
    .Z(_1297_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2819_ (.A1(\mem[11][31] ),
    .A2(_0849_),
    .B(_1297_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2820_ (.A1(_1073_),
    .A2(\mem[5][31] ),
    .A3(_1031_),
    .Z(_1299_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2821_ (.A1(_0595_),
    .A2(\mem[2][31] ),
    .A3(_0963_),
    .Z(_1300_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2822_ (.A1(_1299_),
    .A2(_1300_),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2823_ (.A1(_0734_),
    .A2(_1298_),
    .B1(_1301_),
    .B2(_0800_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2824_ (.A1(\mem[8][31] ),
    .A2(_0810_),
    .B1(_0819_),
    .B2(\mem[9][31] ),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2825_ (.A1(\mem[15][31] ),
    .A2(_0842_),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2826_ (.A1(_0740_),
    .A2(_1303_),
    .B(_1304_),
    .C(_0969_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2827_ (.A1(_1295_),
    .A2(_1296_),
    .B(_1302_),
    .C(_1305_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2828_ (.A1(\mem[0][31] ),
    .A2(_1229_),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2829_ (.A1(net69),
    .A2(_1188_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2830_ (.A1(_1232_),
    .A2(_1306_),
    .A3(_1307_),
    .B(_1308_),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2831_ (.A1(\mem[3][3] ),
    .A2(_0805_),
    .B(_0719_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2832_ (.A1(_1023_),
    .A2(\mem[7][3] ),
    .B1(\mem[4][3] ),
    .B2(_1000_),
    .C1(_0731_),
    .C2(\mem[6][3] ),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2833_ (.A1(\mem[10][3] ),
    .A2(_0813_),
    .B(_1002_),
    .ZN(_1311_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2834_ (.A1(\mem[14][3] ),
    .A2(_0811_),
    .B1(_1004_),
    .B2(\mem[13][3] ),
    .C1(\mem[12][3] ),
    .C2(_0722_),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2835_ (.A1(_1309_),
    .A2(_1310_),
    .B1(_1311_),
    .B2(_1312_),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2836_ (.A1(_1309_),
    .A2(_1311_),
    .B(_0709_),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2837_ (.A1(_0959_),
    .A2(\mem[1][3] ),
    .A3(_0818_),
    .Z(_1315_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2838_ (.A1(\mem[11][3] ),
    .A2(_0849_),
    .B(_1315_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2839_ (.A1(_1073_),
    .A2(\mem[5][3] ),
    .A3(_1031_),
    .Z(_1317_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2840_ (.A1(_0595_),
    .A2(\mem[2][3] ),
    .A3(_0963_),
    .Z(_1318_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2841_ (.A1(_1317_),
    .A2(_1318_),
    .ZN(_1319_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2842_ (.A1(_0734_),
    .A2(_1316_),
    .B1(_1319_),
    .B2(_0800_),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2843_ (.A1(\mem[8][3] ),
    .A2(_0810_),
    .B1(_0819_),
    .B2(\mem[9][3] ),
    .ZN(_1321_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2844_ (.A1(\mem[15][3] ),
    .A2(_0842_),
    .ZN(_1322_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2845_ (.A1(_0740_),
    .A2(_1321_),
    .B(_1322_),
    .C(_0969_),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _2846_ (.A1(_1313_),
    .A2(_1314_),
    .B(_1320_),
    .C(_1323_),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2847_ (.A1(\mem[0][3] ),
    .A2(_1229_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2848_ (.A1(net70),
    .A2(_1188_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2849_ (.A1(_1232_),
    .A2(_1324_),
    .A3(_1325_),
    .B(_1326_),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2850_ (.A1(_0782_),
    .A2(\mem[15][4] ),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2851_ (.A1(\mem[6][4] ),
    .A2(_0724_),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2852_ (.A1(\mem[8][4] ),
    .A2(_0780_),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2853_ (.A1(\mem[1][4] ),
    .A2(_0776_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2854_ (.I0(_1327_),
    .I1(_1328_),
    .I2(_1329_),
    .I3(_1330_),
    .S0(_0716_),
    .S1(_0596_),
    .Z(_1331_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2855_ (.A1(\mem[13][4] ),
    .A2(_0857_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2856_ (.A1(\mem[10][4] ),
    .A2(_0778_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2857_ (.A1(\mem[4][4] ),
    .A2(_0837_),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2858_ (.A1(_0746_),
    .A2(\mem[3][4] ),
    .ZN(_1335_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2859_ (.I0(_1332_),
    .I1(_1333_),
    .I2(_1334_),
    .I3(_1335_),
    .S0(_0865_),
    .S1(_0815_),
    .Z(_1336_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2860_ (.I(\mem[7][4] ),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2861_ (.I(\mem[11][4] ),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2862_ (.A1(_1337_),
    .A2(_0737_),
    .B1(_0739_),
    .B2(_1338_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2863_ (.A1(\mem[2][4] ),
    .A2(_0755_),
    .B1(_0791_),
    .B2(\mem[14][4] ),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2864_ (.I(_1340_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2865_ (.A1(_0809_),
    .A2(_1339_),
    .B1(_1341_),
    .B2(_0817_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2866_ (.A1(_0733_),
    .A2(\mem[12][4] ),
    .A3(_0711_),
    .Z(_1343_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2867_ (.A1(_0992_),
    .A2(\mem[9][4] ),
    .A3(_0712_),
    .Z(_1344_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2868_ (.A1(_1343_),
    .A2(_1344_),
    .Z(_1345_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2869_ (.A1(\mem[5][4] ),
    .A2(_0753_),
    .B1(_1345_),
    .B2(_0807_),
    .C(_0757_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2870_ (.A1(_1331_),
    .A2(_1336_),
    .A3(_1342_),
    .A4(_1346_),
    .Z(_1347_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2871_ (.A1(\mem[0][4] ),
    .A2(_1229_),
    .ZN(_1348_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2872_ (.A1(net71),
    .A2(_1188_),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2873_ (.A1(_1232_),
    .A2(_1347_),
    .A3(_1348_),
    .B(_1349_),
    .ZN(_0542_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2874_ (.A1(\mem[3][5] ),
    .A2(_0805_),
    .B(_0719_),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_4 _2875_ (.A1(_1023_),
    .A2(\mem[7][5] ),
    .B1(\mem[4][5] ),
    .B2(_1000_),
    .C1(_0731_),
    .C2(\mem[6][5] ),
    .ZN(_1351_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2876_ (.A1(\mem[10][5] ),
    .A2(_0813_),
    .B(_1002_),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2877_ (.A1(\mem[14][5] ),
    .A2(_0811_),
    .B1(_1004_),
    .B2(\mem[13][5] ),
    .C1(\mem[12][5] ),
    .C2(_0722_),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2878_ (.A1(_1350_),
    .A2(_1351_),
    .B1(_1352_),
    .B2(_1353_),
    .ZN(_1354_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2879_ (.A1(_1350_),
    .A2(_1352_),
    .B(_0709_),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2880_ (.A1(_0598_),
    .A2(\mem[1][5] ),
    .A3(_0818_),
    .Z(_1356_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2881_ (.A1(\mem[11][5] ),
    .A2(_0849_),
    .B(_1356_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2882_ (.A1(_1073_),
    .A2(\mem[5][5] ),
    .A3(_1031_),
    .Z(_1358_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2883_ (.A1(_0595_),
    .A2(\mem[2][5] ),
    .A3(_0714_),
    .Z(_1359_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2884_ (.A1(_1358_),
    .A2(_1359_),
    .ZN(_1360_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2885_ (.A1(_0734_),
    .A2(_1357_),
    .B1(_1360_),
    .B2(_0800_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2886_ (.A1(\mem[8][5] ),
    .A2(_0810_),
    .B1(_0819_),
    .B2(\mem[9][5] ),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2887_ (.A1(\mem[15][5] ),
    .A2(_0842_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2888_ (.A1(_0740_),
    .A2(_1362_),
    .B(_1363_),
    .C(_0763_),
    .ZN(_1364_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_4 _2889_ (.A1(_1354_),
    .A2(_1355_),
    .B(_1361_),
    .C(_1364_),
    .ZN(_1365_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2890_ (.A1(\mem[0][5] ),
    .A2(_1229_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2891_ (.A1(net72),
    .A2(_1188_),
    .ZN(_1367_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2892_ (.A1(_1232_),
    .A2(_1365_),
    .A3(_1366_),
    .B(_1367_),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2893_ (.A1(_0782_),
    .A2(\mem[15][6] ),
    .ZN(_1368_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2894_ (.A1(\mem[6][6] ),
    .A2(_0724_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2895_ (.A1(\mem[8][6] ),
    .A2(_0780_),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2896_ (.A1(\mem[1][6] ),
    .A2(_0776_),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2897_ (.I0(_1368_),
    .I1(_1369_),
    .I2(_1370_),
    .I3(_1371_),
    .S0(_0716_),
    .S1(_0596_),
    .Z(_1372_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2898_ (.A1(\mem[13][6] ),
    .A2(_0857_),
    .ZN(_1373_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2899_ (.A1(\mem[10][6] ),
    .A2(_0778_),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2900_ (.A1(\mem[4][6] ),
    .A2(_0837_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2901_ (.A1(_0746_),
    .A2(\mem[3][6] ),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2902_ (.I0(_1373_),
    .I1(_1374_),
    .I2(_1375_),
    .I3(_1376_),
    .S0(_0865_),
    .S1(_0815_),
    .Z(_1377_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2903_ (.I(\mem[7][6] ),
    .ZN(_1378_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2904_ (.I(\mem[11][6] ),
    .ZN(_1379_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2905_ (.A1(_1378_),
    .A2(_0737_),
    .B1(_0739_),
    .B2(_1379_),
    .ZN(_1380_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2906_ (.A1(\mem[2][6] ),
    .A2(_0755_),
    .B1(_0791_),
    .B2(\mem[14][6] ),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2907_ (.I(_1381_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2908_ (.A1(_0809_),
    .A2(_1380_),
    .B1(_1382_),
    .B2(_0817_),
    .ZN(_1383_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2909_ (.A1(_0728_),
    .A2(\mem[12][6] ),
    .A3(_0711_),
    .Z(_1384_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2910_ (.A1(_0992_),
    .A2(\mem[9][6] ),
    .A3(_0712_),
    .Z(_1385_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2911_ (.A1(_1384_),
    .A2(_1385_),
    .Z(_1386_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2912_ (.A1(\mem[5][6] ),
    .A2(_0752_),
    .B1(_1386_),
    .B2(_0807_),
    .C(_0757_),
    .ZN(_1387_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2913_ (.A1(_1372_),
    .A2(_1377_),
    .A3(_1383_),
    .A4(_1387_),
    .Z(_1388_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2914_ (.A1(\mem[0][6] ),
    .A2(_1229_),
    .ZN(_1389_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2915_ (.A1(net73),
    .A2(_0761_),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2916_ (.A1(_1232_),
    .A2(_1388_),
    .A3(_1389_),
    .B(_1390_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2917_ (.A1(\mem[3][7] ),
    .A2(_0805_),
    .B(_0719_),
    .ZN(_1391_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_4 _2918_ (.A1(_1023_),
    .A2(\mem[7][7] ),
    .B1(\mem[4][7] ),
    .B2(_0820_),
    .C1(_0731_),
    .C2(\mem[6][7] ),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2919_ (.A1(\mem[10][7] ),
    .A2(_0813_),
    .B(_0774_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2920_ (.A1(\mem[14][7] ),
    .A2(_0811_),
    .B1(_0727_),
    .B2(\mem[13][7] ),
    .C1(\mem[12][7] ),
    .C2(_0722_),
    .ZN(_1394_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2921_ (.A1(_1391_),
    .A2(_1392_),
    .B1(_1393_),
    .B2(_1394_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2922_ (.A1(_1391_),
    .A2(_1393_),
    .B(_0709_),
    .ZN(_1396_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2923_ (.A1(_0598_),
    .A2(\mem[1][7] ),
    .A3(_0818_),
    .Z(_1397_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2924_ (.A1(\mem[11][7] ),
    .A2(_0849_),
    .B(_1397_),
    .ZN(_1398_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2925_ (.A1(_1073_),
    .A2(\mem[5][7] ),
    .A3(_1031_),
    .Z(_1399_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2926_ (.A1(_0595_),
    .A2(\mem[2][7] ),
    .A3(_0714_),
    .Z(_1400_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2927_ (.A1(_1399_),
    .A2(_1400_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2928_ (.A1(_0734_),
    .A2(_1398_),
    .B1(_1401_),
    .B2(_0800_),
    .ZN(_1402_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2929_ (.A1(\mem[8][7] ),
    .A2(_0810_),
    .B1(_0819_),
    .B2(\mem[9][7] ),
    .ZN(_1403_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2930_ (.A1(\mem[15][7] ),
    .A2(_0842_),
    .ZN(_1404_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2931_ (.A1(_0740_),
    .A2(_1403_),
    .B(_1404_),
    .C(_0763_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2932_ (.A1(_1395_),
    .A2(_1396_),
    .B(_1402_),
    .C(_1405_),
    .ZN(_1406_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2933_ (.A1(\mem[0][7] ),
    .A2(_1229_),
    .ZN(_1407_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2934_ (.A1(net74),
    .A2(_0761_),
    .ZN(_1408_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2935_ (.A1(_1232_),
    .A2(_1406_),
    .A3(_1407_),
    .B(_1408_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2936_ (.A1(_0782_),
    .A2(\mem[15][8] ),
    .ZN(_1409_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2937_ (.A1(\mem[6][8] ),
    .A2(_0724_),
    .ZN(_1410_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2938_ (.A1(\mem[8][8] ),
    .A2(_0780_),
    .ZN(_1411_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2939_ (.A1(\mem[1][8] ),
    .A2(_0776_),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2940_ (.I0(_1409_),
    .I1(_1410_),
    .I2(_1411_),
    .I3(_1412_),
    .S0(_0716_),
    .S1(_0596_),
    .Z(_1413_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2941_ (.A1(\mem[13][8] ),
    .A2(_0857_),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2942_ (.A1(\mem[10][8] ),
    .A2(_0832_),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2943_ (.A1(\mem[4][8] ),
    .A2(_0837_),
    .ZN(_1416_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2944_ (.A1(_0746_),
    .A2(\mem[3][8] ),
    .ZN(_1417_));
 gf180mcu_fd_sc_mcu9t5v0__mux4_2 _2945_ (.I0(_1414_),
    .I1(_1415_),
    .I2(_1416_),
    .I3(_1417_),
    .S0(_0865_),
    .S1(_0815_),
    .Z(_1418_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2946_ (.I(\mem[7][8] ),
    .ZN(_1419_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2947_ (.I(\mem[11][8] ),
    .ZN(_1420_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2948_ (.A1(_1419_),
    .A2(_0737_),
    .B1(_0739_),
    .B2(_1420_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2949_ (.A1(\mem[2][8] ),
    .A2(_0755_),
    .B1(_0791_),
    .B2(\mem[14][8] ),
    .ZN(_1422_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _2950_ (.I(_1422_),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2951_ (.A1(_0809_),
    .A2(_1421_),
    .B1(_1423_),
    .B2(_0817_),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2952_ (.A1(_0728_),
    .A2(\mem[12][8] ),
    .A3(_0711_),
    .Z(_1425_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2953_ (.A1(_0992_),
    .A2(\mem[9][8] ),
    .A3(_0712_),
    .Z(_1426_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _2954_ (.A1(_1425_),
    .A2(_1426_),
    .Z(_1427_));
 gf180mcu_fd_sc_mcu9t5v0__aoi221_2 _2955_ (.A1(\mem[5][8] ),
    .A2(_0752_),
    .B1(_1427_),
    .B2(_0807_),
    .C(_0757_),
    .ZN(_1428_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _2956_ (.A1(_1413_),
    .A2(_1418_),
    .A3(_1424_),
    .A4(_1428_),
    .Z(_1429_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2957_ (.A1(\mem[0][8] ),
    .A2(_0764_),
    .ZN(_1430_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2958_ (.A1(net75),
    .A2(_0761_),
    .ZN(_1431_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2959_ (.A1(_1232_),
    .A2(_1429_),
    .A3(_1430_),
    .B(_1431_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2960_ (.A1(\mem[3][9] ),
    .A2(_0805_),
    .B(_0719_),
    .ZN(_1432_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2961_ (.A1(_0743_),
    .A2(\mem[7][9] ),
    .B1(\mem[4][9] ),
    .B2(_0820_),
    .C1(_0731_),
    .C2(\mem[6][9] ),
    .ZN(_1433_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2962_ (.A1(\mem[10][9] ),
    .A2(_0813_),
    .B(_0774_),
    .ZN(_1434_));
 gf180mcu_fd_sc_mcu9t5v0__aoi222_2 _2963_ (.A1(\mem[14][9] ),
    .A2(_0811_),
    .B1(_0727_),
    .B2(\mem[13][9] ),
    .C1(\mem[12][9] ),
    .C2(_0722_),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2964_ (.A1(_1432_),
    .A2(_1433_),
    .B1(_1434_),
    .B2(_1435_),
    .ZN(_1436_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _2965_ (.A1(_1432_),
    .A2(_1434_),
    .B(_0709_),
    .ZN(_1437_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2966_ (.A1(_0598_),
    .A2(\mem[1][9] ),
    .A3(_0818_),
    .Z(_1438_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _2967_ (.A1(\mem[11][9] ),
    .A2(_0849_),
    .B(_1438_),
    .ZN(_1439_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2968_ (.A1(_1073_),
    .A2(\mem[5][9] ),
    .A3(_0827_),
    .Z(_1440_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2969_ (.A1(_0595_),
    .A2(\mem[2][9] ),
    .A3(_0714_),
    .Z(_1441_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2970_ (.A1(_1440_),
    .A2(_1441_),
    .ZN(_1442_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _2971_ (.A1(_0734_),
    .A2(_1439_),
    .B1(_1442_),
    .B2(_0800_),
    .ZN(_1443_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _2972_ (.A1(\mem[8][9] ),
    .A2(_0810_),
    .B1(_0819_),
    .B2(\mem[9][9] ),
    .ZN(_1444_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2973_ (.A1(\mem[15][9] ),
    .A2(_0842_),
    .ZN(_1445_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _2974_ (.A1(_0740_),
    .A2(_1444_),
    .B(_1445_),
    .C(_0763_),
    .ZN(_1446_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _2975_ (.A1(_1436_),
    .A2(_1437_),
    .B(_1443_),
    .C(_1446_),
    .ZN(_1447_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _2976_ (.A1(\mem[0][9] ),
    .A2(_0764_),
    .ZN(_1448_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2977_ (.A1(net76),
    .A2(_0761_),
    .ZN(_1449_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _2978_ (.A1(_0762_),
    .A2(_1447_),
    .A3(_1448_),
    .B(_1449_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _2979_ (.A1(net3),
    .A2(_0593_),
    .Z(_1450_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2980_ (.A1(_0002_),
    .A2(_1450_),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2981_ (.I0(\rd_ptr_bin[1] ),
    .I1(_0003_),
    .S(_1450_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2982_ (.A1(_0809_),
    .A2(_1450_),
    .ZN(_1451_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2983_ (.A1(_0824_),
    .A2(_1451_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _2984_ (.A1(_0728_),
    .A2(\rd_ptr_bin[0] ),
    .A3(\rd_ptr_bin[1] ),
    .Z(_1452_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2985_ (.A1(_1450_),
    .A2(_1452_),
    .Z(_1453_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2986_ (.A1(_1499_),
    .A2(_1453_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2987_ (.A1(\rd_ptr_bin[0] ),
    .A2(_0003_),
    .ZN(_1454_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2988_ (.I0(\rd_ptr_gray[0] ),
    .I1(_1454_),
    .S(_1450_),
    .Z(_0552_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _2989_ (.A1(_0728_),
    .A2(_0710_),
    .A3(_0003_),
    .Z(_1455_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2990_ (.I0(\rd_ptr_gray[1] ),
    .I1(_1455_),
    .S(_1450_),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2991_ (.A1(\rd_ptr_bin[3] ),
    .A2(_1452_),
    .ZN(_1456_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _2992_ (.A1(_0728_),
    .A2(_1519_),
    .A3(_1456_),
    .ZN(_1457_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2993_ (.I0(\rd_ptr_gray[2] ),
    .I1(_1457_),
    .S(_1450_),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _2994_ (.A1(\rd_ptr_bin[4] ),
    .A2(_0842_),
    .A3(_1456_),
    .ZN(_1458_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _2995_ (.I0(\rd_ptr_gray[3] ),
    .I1(_1458_),
    .S(_1450_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _2996_ (.A1(_1450_),
    .A2(_0843_),
    .ZN(_1459_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2997_ (.A1(\rd_ptr_bin[4] ),
    .A2(_1459_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _2998_ (.A1(net37),
    .A2(_0568_),
    .Z(_1460_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _2999_ (.A1(_0000_),
    .A2(_1460_),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3000_ (.I0(\wr_ptr_bin[1] ),
    .I1(_0001_),
    .S(_1460_),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3001_ (.A1(_1512_),
    .A2(_1460_),
    .Z(_1461_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _3002_ (.A1(_0600_),
    .A2(_1461_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _3003_ (.A1(\wr_ptr_bin[2] ),
    .A2(\wr_ptr_bin[0] ),
    .A3(\wr_ptr_bin[1] ),
    .A4(_1460_),
    .Z(_1462_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _3004_ (.A1(_0601_),
    .A2(_1462_),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _3005_ (.A1(\wr_ptr_bin[0] ),
    .A2(_0001_),
    .ZN(_1463_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3006_ (.I0(\wr_ptr_gray[0] ),
    .I1(_1463_),
    .S(_1460_),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _3007_ (.A1(\wr_ptr_bin[2] ),
    .A2(_1512_),
    .A3(_0001_),
    .Z(_1464_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3008_ (.I0(\wr_ptr_gray[1] ),
    .I1(_1464_),
    .S(_1460_),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3009_ (.A1(\wr_ptr_bin[0] ),
    .A2(\wr_ptr_bin[1] ),
    .ZN(_1465_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3010_ (.A1(\wr_ptr_bin[2] ),
    .A2(_1465_),
    .Z(_1466_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _3011_ (.A1(_0601_),
    .A2(_1512_),
    .A3(_1466_),
    .ZN(_1467_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3012_ (.I0(\wr_ptr_gray[2] ),
    .I1(_1467_),
    .S(_1460_),
    .Z(_0563_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3013_ (.A1(\wr_ptr_bin[2] ),
    .A2(_1512_),
    .ZN(_1468_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _3014_ (.A1(\wr_ptr_bin[0] ),
    .A2(\wr_ptr_bin[1] ),
    .B1(_1468_),
    .B2(\wr_ptr_bin[3] ),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_2 _3015_ (.A1(_0600_),
    .A2(_0601_),
    .A3(_1512_),
    .A4(_1465_),
    .ZN(_1470_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _3016_ (.A1(_0602_),
    .A2(_1469_),
    .A3(_1470_),
    .Z(_1471_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _3017_ (.A1(\wr_ptr_bin[4] ),
    .A2(_1471_),
    .ZN(_1472_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _3018_ (.I0(\wr_ptr_gray[3] ),
    .I1(_1472_),
    .S(_1460_),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _3019_ (.A1(_1512_),
    .A2(_0651_),
    .A3(_1460_),
    .Z(_1473_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _3020_ (.A1(\wr_ptr_bin[4] ),
    .A2(_1473_),
    .Z(_0565_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _3021_ (.A1(net40),
    .A2(net41),
    .Z(_1474_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _3022_ (.A1(net42),
    .A2(net77),
    .A3(_1474_),
    .Z(_1475_));
 gf180mcu_fd_sc_mcu9t5v0__nor3_2 _3023_ (.A1(net43),
    .A2(net44),
    .A3(_1475_),
    .ZN(net39));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _3024_ (.I(_1481_),
    .ZN(net80));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _3025_ (.A1(_1480_),
    .A2(_1491_),
    .ZN(net81));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _3026_ (.A1(net80),
    .A2(net81),
    .ZN(_1476_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _3027_ (.A1(_0573_),
    .A2(_1476_),
    .B(_0578_),
    .ZN(net78));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _3028_ (.A(_1477_),
    .B(_1478_),
    .CI(_1479_),
    .CO(_1480_),
    .S(_1481_));
 gf180mcu_fd_sc_mcu9t5v0__addf_1 _3029_ (.A(\rd_ptr_bin[1] ),
    .B(_1483_),
    .CI(_1484_),
    .CO(_1485_),
    .S(_1486_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3030_ (.A(\wr_ptr_bin[1] ),
    .B(_1482_),
    .CO(_1487_),
    .S(_1488_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3031_ (.A(\wr_ptr_bin[2] ),
    .B(_1489_),
    .CO(_1490_),
    .S(_1491_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3032_ (.A(\wr_ptr_bin[3] ),
    .B(_1492_),
    .CO(_1493_),
    .S(_1494_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3033_ (.A(_1495_),
    .B(_1496_),
    .CO(_1497_),
    .S(_1498_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3034_ (.A(_1499_),
    .B(_1500_),
    .CO(_1501_),
    .S(_1502_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3035_ (.A(_1503_),
    .B(_1504_),
    .CO(_1505_),
    .S(_1506_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3036_ (.A(_0000_),
    .B(_1477_),
    .CO(_1507_),
    .S(_0001_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3037_ (.A(_0000_),
    .B(\wr_ptr_bin[1] ),
    .CO(_1508_),
    .S(_1509_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3038_ (.A(\wr_ptr_bin[0] ),
    .B(_1477_),
    .CO(_1510_),
    .S(_1511_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3039_ (.A(\wr_ptr_bin[0] ),
    .B(\wr_ptr_bin[1] ),
    .CO(_1512_),
    .S(_1513_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _3040_ (.A(_0002_),
    .B(_1495_),
    .CO(_1514_),
    .S(_0003_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _3041_ (.A(_0002_),
    .B(\rd_ptr_bin[1] ),
    .CO(_1515_),
    .S(_1516_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _3042_ (.A(\rd_ptr_bin[0] ),
    .B(_1495_),
    .CO(_1517_),
    .S(_1518_));
 gf180mcu_fd_sc_mcu9t5v0__addh_4 _3043_ (.A(\rd_ptr_bin[0] ),
    .B(\rd_ptr_bin[1] ),
    .CO(_1519_),
    .S(_1520_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3044_ (.A(\rd_ptr_bin[0] ),
    .B(_1521_),
    .CO(_1483_),
    .S(_1522_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _3045_ (.A(_0000_),
    .B(_1523_),
    .CO(_1478_),
    .S(_1524_));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][0]$_DFFE_PP_  (.D(_0004_),
    .CLK(clknet_leaf_10_wr_clk),
    .Q(\mem[0][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][10]$_DFFE_PP_  (.D(_0005_),
    .CLK(clknet_leaf_10_wr_clk),
    .Q(\mem[0][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][11]$_DFFE_PP_  (.D(_0006_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[0][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][12]$_DFFE_PP_  (.D(_0007_),
    .CLK(clknet_leaf_10_wr_clk),
    .Q(\mem[0][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][13]$_DFFE_PP_  (.D(_0008_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[0][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][14]$_DFFE_PP_  (.D(_0009_),
    .CLK(clknet_leaf_10_wr_clk),
    .Q(\mem[0][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][15]$_DFFE_PP_  (.D(_0010_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[0][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][16]$_DFFE_PP_  (.D(_0011_),
    .CLK(clknet_leaf_10_wr_clk),
    .Q(\mem[0][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][17]$_DFFE_PP_  (.D(_0012_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[0][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][18]$_DFFE_PP_  (.D(_0013_),
    .CLK(clknet_leaf_10_wr_clk),
    .Q(\mem[0][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][19]$_DFFE_PP_  (.D(_0014_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[0][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][1]$_DFFE_PP_  (.D(_0015_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[0][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][20]$_DFFE_PP_  (.D(_0016_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[0][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][21]$_DFFE_PP_  (.D(_0017_),
    .CLK(clknet_leaf_4_wr_clk),
    .Q(\mem[0][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][22]$_DFFE_PP_  (.D(_0018_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[0][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][23]$_DFFE_PP_  (.D(_0019_),
    .CLK(clknet_leaf_4_wr_clk),
    .Q(\mem[0][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][24]$_DFFE_PP_  (.D(_0020_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[0][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][25]$_DFFE_PP_  (.D(_0021_),
    .CLK(clknet_leaf_2_wr_clk),
    .Q(\mem[0][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][26]$_DFFE_PP_  (.D(_0022_),
    .CLK(clknet_leaf_2_wr_clk),
    .Q(\mem[0][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][27]$_DFFE_PP_  (.D(_0023_),
    .CLK(clknet_leaf_2_wr_clk),
    .Q(\mem[0][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][28]$_DFFE_PP_  (.D(_0024_),
    .CLK(clknet_leaf_18_wr_clk),
    .Q(\mem[0][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][29]$_DFFE_PP_  (.D(_0025_),
    .CLK(clknet_leaf_18_wr_clk),
    .Q(\mem[0][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][2]$_DFFE_PP_  (.D(_0026_),
    .CLK(clknet_leaf_18_wr_clk),
    .Q(\mem[0][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][30]$_DFFE_PP_  (.D(_0027_),
    .CLK(clknet_leaf_18_wr_clk),
    .Q(\mem[0][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][31]$_DFFE_PP_  (.D(_0028_),
    .CLK(clknet_leaf_19_wr_clk),
    .Q(\mem[0][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][3]$_DFFE_PP_  (.D(_0029_),
    .CLK(clknet_leaf_19_wr_clk),
    .Q(\mem[0][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][4]$_DFFE_PP_  (.D(_0030_),
    .CLK(clknet_leaf_18_wr_clk),
    .Q(\mem[0][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][5]$_DFFE_PP_  (.D(_0031_),
    .CLK(clknet_leaf_18_wr_clk),
    .Q(\mem[0][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][6]$_DFFE_PP_  (.D(_0032_),
    .CLK(clknet_leaf_15_wr_clk),
    .Q(\mem[0][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][7]$_DFFE_PP_  (.D(_0033_),
    .CLK(clknet_leaf_17_wr_clk),
    .Q(\mem[0][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][8]$_DFFE_PP_  (.D(_0034_),
    .CLK(clknet_leaf_14_wr_clk),
    .Q(\mem[0][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[0][9]$_DFFE_PP_  (.D(_0035_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[0][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][0]$_DFFE_PP_  (.D(_0036_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[10][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][10]$_DFFE_PP_  (.D(_0037_),
    .CLK(clknet_leaf_10_wr_clk),
    .Q(\mem[10][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][11]$_DFFE_PP_  (.D(_0038_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[10][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][12]$_DFFE_PP_  (.D(_0039_),
    .CLK(clknet_leaf_10_wr_clk),
    .Q(\mem[10][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][13]$_DFFE_PP_  (.D(_0040_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[10][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][14]$_DFFE_PP_  (.D(_0041_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[10][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][15]$_DFFE_PP_  (.D(_0042_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[10][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][16]$_DFFE_PP_  (.D(_0043_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[10][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][17]$_DFFE_PP_  (.D(_0044_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[10][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][18]$_DFFE_PP_  (.D(_0045_),
    .CLK(clknet_leaf_10_wr_clk),
    .Q(\mem[10][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][19]$_DFFE_PP_  (.D(_0046_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[10][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][1]$_DFFE_PP_  (.D(_0047_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[10][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][20]$_DFFE_PP_  (.D(_0048_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[10][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][21]$_DFFE_PP_  (.D(_0049_),
    .CLK(clknet_leaf_4_wr_clk),
    .Q(\mem[10][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][22]$_DFFE_PP_  (.D(_0050_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[10][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][23]$_DFFE_PP_  (.D(_0051_),
    .CLK(clknet_leaf_4_wr_clk),
    .Q(\mem[10][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][24]$_DFFE_PP_  (.D(_0052_),
    .CLK(clknet_leaf_6_wr_clk),
    .Q(\mem[10][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][25]$_DFFE_PP_  (.D(_0053_),
    .CLK(clknet_leaf_2_wr_clk),
    .Q(\mem[10][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][26]$_DFFE_PP_  (.D(_0054_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[10][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][27]$_DFFE_PP_  (.D(_0055_),
    .CLK(clknet_leaf_2_wr_clk),
    .Q(\mem[10][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][28]$_DFFE_PP_  (.D(_0056_),
    .CLK(clknet_leaf_18_wr_clk),
    .Q(\mem[10][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][29]$_DFFE_PP_  (.D(_0057_),
    .CLK(clknet_leaf_0_wr_clk),
    .Q(\mem[10][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][2]$_DFFE_PP_  (.D(_0058_),
    .CLK(clknet_leaf_18_wr_clk),
    .Q(\mem[10][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][30]$_DFFE_PP_  (.D(_0059_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[10][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][31]$_DFFE_PP_  (.D(_0060_),
    .CLK(clknet_leaf_19_wr_clk),
    .Q(\mem[10][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][3]$_DFFE_PP_  (.D(_0061_),
    .CLK(clknet_leaf_19_wr_clk),
    .Q(\mem[10][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][4]$_DFFE_PP_  (.D(_0062_),
    .CLK(clknet_leaf_15_wr_clk),
    .Q(\mem[10][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][5]$_DFFE_PP_  (.D(_0063_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[10][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][6]$_DFFE_PP_  (.D(_0064_),
    .CLK(clknet_leaf_15_wr_clk),
    .Q(\mem[10][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][7]$_DFFE_PP_  (.D(_0065_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[10][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][8]$_DFFE_PP_  (.D(_0066_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[10][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[10][9]$_DFFE_PP_  (.D(_0067_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[10][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][0]$_DFFE_PP_  (.D(_0068_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[11][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][10]$_DFFE_PP_  (.D(_0069_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[11][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][11]$_DFFE_PP_  (.D(_0070_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[11][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][12]$_DFFE_PP_  (.D(_0071_),
    .CLK(clknet_leaf_13_wr_clk),
    .Q(\mem[11][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][13]$_DFFE_PP_  (.D(_0072_),
    .CLK(clknet_leaf_10_wr_clk),
    .Q(\mem[11][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][14]$_DFFE_PP_  (.D(_0073_),
    .CLK(clknet_leaf_13_wr_clk),
    .Q(\mem[11][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][15]$_DFFE_PP_  (.D(_0074_),
    .CLK(clknet_leaf_10_wr_clk),
    .Q(\mem[11][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][16]$_DFFE_PP_  (.D(_0075_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[11][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][17]$_DFFE_PP_  (.D(_0076_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[11][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][18]$_DFFE_PP_  (.D(_0077_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[11][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][19]$_DFFE_PP_  (.D(_0078_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[11][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][1]$_DFFE_PP_  (.D(_0079_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[11][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][20]$_DFFE_PP_  (.D(_0080_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[11][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][21]$_DFFE_PP_  (.D(_0081_),
    .CLK(clknet_leaf_4_wr_clk),
    .Q(\mem[11][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][22]$_DFFE_PP_  (.D(_0082_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[11][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][23]$_DFFE_PP_  (.D(_0083_),
    .CLK(clknet_leaf_4_wr_clk),
    .Q(\mem[11][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][24]$_DFFE_PP_  (.D(_0084_),
    .CLK(clknet_leaf_6_wr_clk),
    .Q(\mem[11][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][25]$_DFFE_PP_  (.D(_0085_),
    .CLK(clknet_leaf_2_wr_clk),
    .Q(\mem[11][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][26]$_DFFE_PP_  (.D(_0086_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[11][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][27]$_DFFE_PP_  (.D(_0087_),
    .CLK(clknet_leaf_2_wr_clk),
    .Q(\mem[11][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][28]$_DFFE_PP_  (.D(_0088_),
    .CLK(clknet_leaf_17_wr_clk),
    .Q(\mem[11][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][29]$_DFFE_PP_  (.D(_0089_),
    .CLK(clknet_leaf_0_wr_clk),
    .Q(\mem[11][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][2]$_DFFE_PP_  (.D(_0090_),
    .CLK(clknet_leaf_17_wr_clk),
    .Q(\mem[11][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][30]$_DFFE_PP_  (.D(_0091_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[11][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][31]$_DFFE_PP_  (.D(_0092_),
    .CLK(clknet_leaf_0_wr_clk),
    .Q(\mem[11][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][3]$_DFFE_PP_  (.D(_0093_),
    .CLK(clknet_leaf_0_wr_clk),
    .Q(\mem[11][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][4]$_DFFE_PP_  (.D(_0094_),
    .CLK(clknet_leaf_17_wr_clk),
    .Q(\mem[11][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][5]$_DFFE_PP_  (.D(_0095_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[11][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][6]$_DFFE_PP_  (.D(_0096_),
    .CLK(clknet_leaf_15_wr_clk),
    .Q(\mem[11][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][7]$_DFFE_PP_  (.D(_0097_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[11][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][8]$_DFFE_PP_  (.D(_0098_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[11][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[11][9]$_DFFE_PP_  (.D(_0099_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[11][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][0]$_DFFE_PP_  (.D(_0100_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[12][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][10]$_DFFE_PP_  (.D(_0101_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[12][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][11]$_DFFE_PP_  (.D(_0102_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[12][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][12]$_DFFE_PP_  (.D(_0103_),
    .CLK(clknet_leaf_10_wr_clk),
    .Q(\mem[12][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][13]$_DFFE_PP_  (.D(_0104_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[12][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][14]$_DFFE_PP_  (.D(_0105_),
    .CLK(clknet_leaf_13_wr_clk),
    .Q(\mem[12][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][15]$_DFFE_PP_  (.D(_0106_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[12][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][16]$_DFFE_PP_  (.D(_0107_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[12][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][17]$_DFFE_PP_  (.D(_0108_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[12][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][18]$_DFFE_PP_  (.D(_0109_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[12][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][19]$_DFFE_PP_  (.D(_0110_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[12][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][1]$_DFFE_PP_  (.D(_0111_),
    .CLK(clknet_leaf_4_wr_clk),
    .Q(\mem[12][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][20]$_DFFE_PP_  (.D(_0112_),
    .CLK(clknet_leaf_6_wr_clk),
    .Q(\mem[12][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][21]$_DFFE_PP_  (.D(_0113_),
    .CLK(clknet_leaf_4_wr_clk),
    .Q(\mem[12][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][22]$_DFFE_PP_  (.D(_0114_),
    .CLK(clknet_leaf_6_wr_clk),
    .Q(\mem[12][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][23]$_DFFE_PP_  (.D(_0115_),
    .CLK(clknet_leaf_4_wr_clk),
    .Q(\mem[12][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][24]$_DFFE_PP_  (.D(_0116_),
    .CLK(clknet_leaf_6_wr_clk),
    .Q(\mem[12][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][25]$_DFFE_PP_  (.D(_0117_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[12][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][26]$_DFFE_PP_  (.D(_0118_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[12][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][27]$_DFFE_PP_  (.D(_0119_),
    .CLK(clknet_leaf_2_wr_clk),
    .Q(\mem[12][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][28]$_DFFE_PP_  (.D(_0120_),
    .CLK(clknet_leaf_17_wr_clk),
    .Q(\mem[12][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][29]$_DFFE_PP_  (.D(_0121_),
    .CLK(clknet_leaf_19_wr_clk),
    .Q(\mem[12][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][2]$_DFFE_PP_  (.D(_0122_),
    .CLK(clknet_leaf_17_wr_clk),
    .Q(\mem[12][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][30]$_DFFE_PP_  (.D(_0123_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[12][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][31]$_DFFE_PP_  (.D(_0124_),
    .CLK(clknet_leaf_19_wr_clk),
    .Q(\mem[12][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][3]$_DFFE_PP_  (.D(_0125_),
    .CLK(clknet_leaf_19_wr_clk),
    .Q(\mem[12][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][4]$_DFFE_PP_  (.D(_0126_),
    .CLK(clknet_leaf_17_wr_clk),
    .Q(\mem[12][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][5]$_DFFE_PP_  (.D(_0127_),
    .CLK(clknet_leaf_18_wr_clk),
    .Q(\mem[12][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][6]$_DFFE_PP_  (.D(_0128_),
    .CLK(clknet_leaf_15_wr_clk),
    .Q(\mem[12][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][7]$_DFFE_PP_  (.D(_0129_),
    .CLK(clknet_leaf_17_wr_clk),
    .Q(\mem[12][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][8]$_DFFE_PP_  (.D(_0130_),
    .CLK(clknet_leaf_15_wr_clk),
    .Q(\mem[12][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[12][9]$_DFFE_PP_  (.D(_0131_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[12][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][0]$_DFFE_PP_  (.D(_0132_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[13][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][10]$_DFFE_PP_  (.D(_0133_),
    .CLK(clknet_leaf_10_wr_clk),
    .Q(\mem[13][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][11]$_DFFE_PP_  (.D(_0134_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[13][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][12]$_DFFE_PP_  (.D(_0135_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[13][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][13]$_DFFE_PP_  (.D(_0136_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[13][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][14]$_DFFE_PP_  (.D(_0137_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[13][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][15]$_DFFE_PP_  (.D(_0138_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[13][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][16]$_DFFE_PP_  (.D(_0139_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[13][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][17]$_DFFE_PP_  (.D(_0140_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[13][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][18]$_DFFE_PP_  (.D(_0141_),
    .CLK(clknet_leaf_10_wr_clk),
    .Q(\mem[13][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][19]$_DFFE_PP_  (.D(_0142_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[13][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][1]$_DFFE_PP_  (.D(_0143_),
    .CLK(clknet_leaf_4_wr_clk),
    .Q(\mem[13][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][20]$_DFFE_PP_  (.D(_0144_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[13][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][21]$_DFFE_PP_  (.D(_0145_),
    .CLK(clknet_leaf_4_wr_clk),
    .Q(\mem[13][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][22]$_DFFE_PP_  (.D(_0146_),
    .CLK(clknet_leaf_6_wr_clk),
    .Q(\mem[13][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][23]$_DFFE_PP_  (.D(_0147_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[13][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][24]$_DFFE_PP_  (.D(_0148_),
    .CLK(clknet_leaf_6_wr_clk),
    .Q(\mem[13][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][25]$_DFFE_PP_  (.D(_0149_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[13][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][26]$_DFFE_PP_  (.D(_0150_),
    .CLK(clknet_leaf_6_wr_clk),
    .Q(\mem[13][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][27]$_DFFE_PP_  (.D(_0151_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[13][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][28]$_DFFE_PP_  (.D(_0152_),
    .CLK(clknet_leaf_18_wr_clk),
    .Q(\mem[13][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][29]$_DFFE_PP_  (.D(_0153_),
    .CLK(clknet_leaf_19_wr_clk),
    .Q(\mem[13][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][2]$_DFFE_PP_  (.D(_0154_),
    .CLK(clknet_leaf_18_wr_clk),
    .Q(\mem[13][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][30]$_DFFE_PP_  (.D(_0155_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[13][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][31]$_DFFE_PP_  (.D(_0156_),
    .CLK(clknet_leaf_19_wr_clk),
    .Q(\mem[13][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][3]$_DFFE_PP_  (.D(_0157_),
    .CLK(clknet_leaf_19_wr_clk),
    .Q(\mem[13][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][4]$_DFFE_PP_  (.D(_0158_),
    .CLK(clknet_leaf_15_wr_clk),
    .Q(\mem[13][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][5]$_DFFE_PP_  (.D(_0159_),
    .CLK(clknet_leaf_18_wr_clk),
    .Q(\mem[13][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][6]$_DFFE_PP_  (.D(_0160_),
    .CLK(clknet_leaf_15_wr_clk),
    .Q(\mem[13][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][7]$_DFFE_PP_  (.D(_0161_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[13][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][8]$_DFFE_PP_  (.D(_0162_),
    .CLK(clknet_leaf_14_wr_clk),
    .Q(\mem[13][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[13][9]$_DFFE_PP_  (.D(_0163_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[13][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][0]$_DFFE_PP_  (.D(_0164_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[14][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][10]$_DFFE_PP_  (.D(_0165_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[14][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][11]$_DFFE_PP_  (.D(_0166_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[14][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][12]$_DFFE_PP_  (.D(_0167_),
    .CLK(clknet_leaf_13_wr_clk),
    .Q(\mem[14][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][13]$_DFFE_PP_  (.D(_0168_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[14][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][14]$_DFFE_PP_  (.D(_0169_),
    .CLK(clknet_leaf_13_wr_clk),
    .Q(\mem[14][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][15]$_DFFE_PP_  (.D(_0170_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[14][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][16]$_DFFE_PP_  (.D(_0171_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[14][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][17]$_DFFE_PP_  (.D(_0172_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[14][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][18]$_DFFE_PP_  (.D(_0173_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[14][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][19]$_DFFE_PP_  (.D(_0174_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[14][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][1]$_DFFE_PP_  (.D(_0175_),
    .CLK(clknet_leaf_4_wr_clk),
    .Q(\mem[14][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][20]$_DFFE_PP_  (.D(_0176_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[14][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][21]$_DFFE_PP_  (.D(_0177_),
    .CLK(clknet_leaf_4_wr_clk),
    .Q(\mem[14][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][22]$_DFFE_PP_  (.D(_0178_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[14][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][23]$_DFFE_PP_  (.D(_0179_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[14][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][24]$_DFFE_PP_  (.D(_0180_),
    .CLK(clknet_leaf_2_wr_clk),
    .Q(\mem[14][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][25]$_DFFE_PP_  (.D(_0181_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[14][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][26]$_DFFE_PP_  (.D(_0182_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[14][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][27]$_DFFE_PP_  (.D(_0183_),
    .CLK(clknet_leaf_2_wr_clk),
    .Q(\mem[14][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][28]$_DFFE_PP_  (.D(_0184_),
    .CLK(clknet_leaf_18_wr_clk),
    .Q(\mem[14][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][29]$_DFFE_PP_  (.D(_0185_),
    .CLK(clknet_leaf_18_wr_clk),
    .Q(\mem[14][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][2]$_DFFE_PP_  (.D(_0186_),
    .CLK(clknet_leaf_17_wr_clk),
    .Q(\mem[14][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][30]$_DFFE_PP_  (.D(_0187_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[14][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][31]$_DFFE_PP_  (.D(_0188_),
    .CLK(clknet_leaf_19_wr_clk),
    .Q(\mem[14][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][3]$_DFFE_PP_  (.D(_0189_),
    .CLK(clknet_leaf_19_wr_clk),
    .Q(\mem[14][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][4]$_DFFE_PP_  (.D(_0190_),
    .CLK(clknet_leaf_15_wr_clk),
    .Q(\mem[14][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][5]$_DFFE_PP_  (.D(_0191_),
    .CLK(clknet_leaf_18_wr_clk),
    .Q(\mem[14][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][6]$_DFFE_PP_  (.D(_0192_),
    .CLK(clknet_leaf_15_wr_clk),
    .Q(\mem[14][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][7]$_DFFE_PP_  (.D(_0193_),
    .CLK(clknet_leaf_17_wr_clk),
    .Q(\mem[14][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][8]$_DFFE_PP_  (.D(_0194_),
    .CLK(clknet_leaf_15_wr_clk),
    .Q(\mem[14][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[14][9]$_DFFE_PP_  (.D(_0195_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[14][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][0]$_DFFE_PP_  (.D(_0196_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[15][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][10]$_DFFE_PP_  (.D(_0197_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[15][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][11]$_DFFE_PP_  (.D(_0198_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[15][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][12]$_DFFE_PP_  (.D(_0199_),
    .CLK(clknet_leaf_13_wr_clk),
    .Q(\mem[15][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][13]$_DFFE_PP_  (.D(_0200_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[15][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][14]$_DFFE_PP_  (.D(_0201_),
    .CLK(clknet_leaf_13_wr_clk),
    .Q(\mem[15][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][15]$_DFFE_PP_  (.D(_0202_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[15][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][16]$_DFFE_PP_  (.D(_0203_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[15][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][17]$_DFFE_PP_  (.D(_0204_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[15][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][18]$_DFFE_PP_  (.D(_0205_),
    .CLK(clknet_leaf_10_wr_clk),
    .Q(\mem[15][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][19]$_DFFE_PP_  (.D(_0206_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[15][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][1]$_DFFE_PP_  (.D(_0207_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[15][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][20]$_DFFE_PP_  (.D(_0208_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[15][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][21]$_DFFE_PP_  (.D(_0209_),
    .CLK(clknet_leaf_4_wr_clk),
    .Q(\mem[15][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][22]$_DFFE_PP_  (.D(_0210_),
    .CLK(clknet_leaf_6_wr_clk),
    .Q(\mem[15][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][23]$_DFFE_PP_  (.D(_0211_),
    .CLK(clknet_leaf_4_wr_clk),
    .Q(\mem[15][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][24]$_DFFE_PP_  (.D(_0212_),
    .CLK(clknet_leaf_2_wr_clk),
    .Q(\mem[15][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][25]$_DFFE_PP_  (.D(_0213_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[15][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][26]$_DFFE_PP_  (.D(_0214_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[15][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][27]$_DFFE_PP_  (.D(_0215_),
    .CLK(clknet_leaf_2_wr_clk),
    .Q(\mem[15][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][28]$_DFFE_PP_  (.D(_0216_),
    .CLK(clknet_leaf_18_wr_clk),
    .Q(\mem[15][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][29]$_DFFE_PP_  (.D(_0217_),
    .CLK(clknet_leaf_0_wr_clk),
    .Q(\mem[15][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][2]$_DFFE_PP_  (.D(_0218_),
    .CLK(clknet_leaf_17_wr_clk),
    .Q(\mem[15][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][30]$_DFFE_PP_  (.D(_0219_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[15][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][31]$_DFFE_PP_  (.D(_0220_),
    .CLK(clknet_leaf_19_wr_clk),
    .Q(\mem[15][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][3]$_DFFE_PP_  (.D(_0221_),
    .CLK(clknet_leaf_19_wr_clk),
    .Q(\mem[15][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][4]$_DFFE_PP_  (.D(_0222_),
    .CLK(clknet_leaf_15_wr_clk),
    .Q(\mem[15][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][5]$_DFFE_PP_  (.D(_0223_),
    .CLK(clknet_leaf_18_wr_clk),
    .Q(\mem[15][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][6]$_DFFE_PP_  (.D(_0224_),
    .CLK(clknet_leaf_15_wr_clk),
    .Q(\mem[15][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][7]$_DFFE_PP_  (.D(_0225_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[15][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][8]$_DFFE_PP_  (.D(_0226_),
    .CLK(clknet_leaf_14_wr_clk),
    .Q(\mem[15][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[15][9]$_DFFE_PP_  (.D(_0227_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[15][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][0]$_DFFE_PP_  (.D(_0228_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[1][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][10]$_DFFE_PP_  (.D(_0229_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[1][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][11]$_DFFE_PP_  (.D(_0230_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[1][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][12]$_DFFE_PP_  (.D(_0231_),
    .CLK(clknet_leaf_13_wr_clk),
    .Q(\mem[1][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][13]$_DFFE_PP_  (.D(_0232_),
    .CLK(clknet_leaf_10_wr_clk),
    .Q(\mem[1][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][14]$_DFFE_PP_  (.D(_0233_),
    .CLK(clknet_leaf_13_wr_clk),
    .Q(\mem[1][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][15]$_DFFE_PP_  (.D(_0234_),
    .CLK(clknet_leaf_10_wr_clk),
    .Q(\mem[1][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][16]$_DFFE_PP_  (.D(_0235_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[1][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][17]$_DFFE_PP_  (.D(_0236_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[1][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][18]$_DFFE_PP_  (.D(_0237_),
    .CLK(clknet_leaf_10_wr_clk),
    .Q(\mem[1][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][19]$_DFFE_PP_  (.D(_0238_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[1][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][1]$_DFFE_PP_  (.D(_0239_),
    .CLK(clknet_leaf_6_wr_clk),
    .Q(\mem[1][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][20]$_DFFE_PP_  (.D(_0240_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[1][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][21]$_DFFE_PP_  (.D(_0241_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[1][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][22]$_DFFE_PP_  (.D(_0242_),
    .CLK(clknet_leaf_6_wr_clk),
    .Q(\mem[1][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][23]$_DFFE_PP_  (.D(_0243_),
    .CLK(clknet_leaf_4_wr_clk),
    .Q(\mem[1][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][24]$_DFFE_PP_  (.D(_0244_),
    .CLK(clknet_leaf_2_wr_clk),
    .Q(\mem[1][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][25]$_DFFE_PP_  (.D(_0245_),
    .CLK(clknet_leaf_2_wr_clk),
    .Q(\mem[1][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][26]$_DFFE_PP_  (.D(_0246_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[1][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][27]$_DFFE_PP_  (.D(_0247_),
    .CLK(clknet_leaf_2_wr_clk),
    .Q(\mem[1][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][28]$_DFFE_PP_  (.D(_0248_),
    .CLK(clknet_leaf_18_wr_clk),
    .Q(\mem[1][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][29]$_DFFE_PP_  (.D(_0249_),
    .CLK(clknet_leaf_2_wr_clk),
    .Q(\mem[1][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][2]$_DFFE_PP_  (.D(_0250_),
    .CLK(clknet_leaf_18_wr_clk),
    .Q(\mem[1][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][30]$_DFFE_PP_  (.D(_0251_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[1][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][31]$_DFFE_PP_  (.D(_0252_),
    .CLK(clknet_leaf_0_wr_clk),
    .Q(\mem[1][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][3]$_DFFE_PP_  (.D(_0253_),
    .CLK(clknet_leaf_0_wr_clk),
    .Q(\mem[1][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][4]$_DFFE_PP_  (.D(_0254_),
    .CLK(clknet_leaf_17_wr_clk),
    .Q(\mem[1][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][5]$_DFFE_PP_  (.D(_0255_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[1][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][6]$_DFFE_PP_  (.D(_0256_),
    .CLK(clknet_leaf_15_wr_clk),
    .Q(\mem[1][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][7]$_DFFE_PP_  (.D(_0257_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[1][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][8]$_DFFE_PP_  (.D(_0258_),
    .CLK(clknet_leaf_15_wr_clk),
    .Q(\mem[1][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[1][9]$_DFFE_PP_  (.D(_0259_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[1][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][0]$_DFFE_PP_  (.D(_0260_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[2][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][10]$_DFFE_PP_  (.D(_0261_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[2][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][11]$_DFFE_PP_  (.D(_0262_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[2][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][12]$_DFFE_PP_  (.D(_0263_),
    .CLK(clknet_leaf_10_wr_clk),
    .Q(\mem[2][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][13]$_DFFE_PP_  (.D(_0264_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[2][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][14]$_DFFE_PP_  (.D(_0265_),
    .CLK(clknet_leaf_13_wr_clk),
    .Q(\mem[2][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][15]$_DFFE_PP_  (.D(_0266_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[2][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][16]$_DFFE_PP_  (.D(_0267_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[2][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][17]$_DFFE_PP_  (.D(_0268_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[2][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][18]$_DFFE_PP_  (.D(_0269_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[2][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][19]$_DFFE_PP_  (.D(_0270_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[2][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][1]$_DFFE_PP_  (.D(_0271_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[2][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][20]$_DFFE_PP_  (.D(_0272_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[2][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][21]$_DFFE_PP_  (.D(_0273_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[2][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][22]$_DFFE_PP_  (.D(_0274_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[2][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][23]$_DFFE_PP_  (.D(_0275_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[2][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][24]$_DFFE_PP_  (.D(_0276_),
    .CLK(clknet_leaf_6_wr_clk),
    .Q(\mem[2][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][25]$_DFFE_PP_  (.D(_0277_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[2][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][26]$_DFFE_PP_  (.D(_0278_),
    .CLK(clknet_leaf_2_wr_clk),
    .Q(\mem[2][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][27]$_DFFE_PP_  (.D(_0279_),
    .CLK(clknet_leaf_2_wr_clk),
    .Q(\mem[2][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][28]$_DFFE_PP_  (.D(_0280_),
    .CLK(clknet_leaf_18_wr_clk),
    .Q(\mem[2][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][29]$_DFFE_PP_  (.D(_0281_),
    .CLK(clknet_leaf_0_wr_clk),
    .Q(\mem[2][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][2]$_DFFE_PP_  (.D(_0282_),
    .CLK(clknet_leaf_17_wr_clk),
    .Q(\mem[2][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][30]$_DFFE_PP_  (.D(_0283_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[2][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][31]$_DFFE_PP_  (.D(_0284_),
    .CLK(clknet_leaf_0_wr_clk),
    .Q(\mem[2][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][3]$_DFFE_PP_  (.D(_0285_),
    .CLK(clknet_leaf_0_wr_clk),
    .Q(\mem[2][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][4]$_DFFE_PP_  (.D(_0286_),
    .CLK(clknet_leaf_15_wr_clk),
    .Q(\mem[2][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][5]$_DFFE_PP_  (.D(_0287_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[2][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][6]$_DFFE_PP_  (.D(_0288_),
    .CLK(clknet_leaf_15_wr_clk),
    .Q(\mem[2][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][7]$_DFFE_PP_  (.D(_0289_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[2][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][8]$_DFFE_PP_  (.D(_0290_),
    .CLK(clknet_leaf_14_wr_clk),
    .Q(\mem[2][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[2][9]$_DFFE_PP_  (.D(_0291_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[2][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][0]$_DFFE_PP_  (.D(_0292_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[3][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][10]$_DFFE_PP_  (.D(_0293_),
    .CLK(clknet_leaf_10_wr_clk),
    .Q(\mem[3][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][11]$_DFFE_PP_  (.D(_0294_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[3][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][12]$_DFFE_PP_  (.D(_0295_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[3][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][13]$_DFFE_PP_  (.D(_0296_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[3][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][14]$_DFFE_PP_  (.D(_0297_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[3][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][15]$_DFFE_PP_  (.D(_0298_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[3][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][16]$_DFFE_PP_  (.D(_0299_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[3][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][17]$_DFFE_PP_  (.D(_0300_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[3][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][18]$_DFFE_PP_  (.D(_0301_),
    .CLK(clknet_leaf_10_wr_clk),
    .Q(\mem[3][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][19]$_DFFE_PP_  (.D(_0302_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[3][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][1]$_DFFE_PP_  (.D(_0303_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[3][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][20]$_DFFE_PP_  (.D(_0304_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[3][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][21]$_DFFE_PP_  (.D(_0305_),
    .CLK(clknet_leaf_4_wr_clk),
    .Q(\mem[3][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][22]$_DFFE_PP_  (.D(_0306_),
    .CLK(clknet_leaf_6_wr_clk),
    .Q(\mem[3][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][23]$_DFFE_PP_  (.D(_0307_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[3][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][24]$_DFFE_PP_  (.D(_0308_),
    .CLK(clknet_leaf_6_wr_clk),
    .Q(\mem[3][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][25]$_DFFE_PP_  (.D(_0309_),
    .CLK(clknet_leaf_2_wr_clk),
    .Q(\mem[3][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][26]$_DFFE_PP_  (.D(_0310_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[3][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][27]$_DFFE_PP_  (.D(_0311_),
    .CLK(clknet_leaf_2_wr_clk),
    .Q(\mem[3][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][28]$_DFFE_PP_  (.D(_0312_),
    .CLK(clknet_leaf_18_wr_clk),
    .Q(\mem[3][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][29]$_DFFE_PP_  (.D(_0313_),
    .CLK(clknet_leaf_0_wr_clk),
    .Q(\mem[3][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][2]$_DFFE_PP_  (.D(_0314_),
    .CLK(clknet_leaf_18_wr_clk),
    .Q(\mem[3][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][30]$_DFFE_PP_  (.D(_0315_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[3][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][31]$_DFFE_PP_  (.D(_0316_),
    .CLK(clknet_leaf_0_wr_clk),
    .Q(\mem[3][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][3]$_DFFE_PP_  (.D(_0317_),
    .CLK(clknet_leaf_19_wr_clk),
    .Q(\mem[3][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][4]$_DFFE_PP_  (.D(_0318_),
    .CLK(clknet_leaf_17_wr_clk),
    .Q(\mem[3][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][5]$_DFFE_PP_  (.D(_0319_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[3][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][6]$_DFFE_PP_  (.D(_0320_),
    .CLK(clknet_leaf_15_wr_clk),
    .Q(\mem[3][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][7]$_DFFE_PP_  (.D(_0321_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[3][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][8]$_DFFE_PP_  (.D(_0322_),
    .CLK(clknet_leaf_14_wr_clk),
    .Q(\mem[3][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[3][9]$_DFFE_PP_  (.D(_0323_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[3][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][0]$_DFFE_PP_  (.D(_0324_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[4][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][10]$_DFFE_PP_  (.D(_0325_),
    .CLK(clknet_leaf_10_wr_clk),
    .Q(\mem[4][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][11]$_DFFE_PP_  (.D(_0326_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[4][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][12]$_DFFE_PP_  (.D(_0327_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[4][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][13]$_DFFE_PP_  (.D(_0328_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[4][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][14]$_DFFE_PP_  (.D(_0329_),
    .CLK(clknet_leaf_13_wr_clk),
    .Q(\mem[4][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][15]$_DFFE_PP_  (.D(_0330_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[4][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][16]$_DFFE_PP_  (.D(_0331_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[4][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][17]$_DFFE_PP_  (.D(_0332_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[4][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][18]$_DFFE_PP_  (.D(_0333_),
    .CLK(clknet_leaf_10_wr_clk),
    .Q(\mem[4][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][19]$_DFFE_PP_  (.D(_0334_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[4][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][1]$_DFFE_PP_  (.D(_0335_),
    .CLK(clknet_leaf_4_wr_clk),
    .Q(\mem[4][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][20]$_DFFE_PP_  (.D(_0336_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[4][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][21]$_DFFE_PP_  (.D(_0337_),
    .CLK(clknet_leaf_4_wr_clk),
    .Q(\mem[4][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][22]$_DFFE_PP_  (.D(_0338_),
    .CLK(clknet_leaf_6_wr_clk),
    .Q(\mem[4][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][23]$_DFFE_PP_  (.D(_0339_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[4][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][24]$_DFFE_PP_  (.D(_0340_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[4][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][25]$_DFFE_PP_  (.D(_0341_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[4][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][26]$_DFFE_PP_  (.D(_0342_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[4][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][27]$_DFFE_PP_  (.D(_0343_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[4][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][28]$_DFFE_PP_  (.D(_0344_),
    .CLK(clknet_leaf_18_wr_clk),
    .Q(\mem[4][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][29]$_DFFE_PP_  (.D(_0345_),
    .CLK(clknet_leaf_0_wr_clk),
    .Q(\mem[4][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][2]$_DFFE_PP_  (.D(_0346_),
    .CLK(clknet_leaf_18_wr_clk),
    .Q(\mem[4][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][30]$_DFFE_PP_  (.D(_0347_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[4][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][31]$_DFFE_PP_  (.D(_0348_),
    .CLK(clknet_leaf_19_wr_clk),
    .Q(\mem[4][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][3]$_DFFE_PP_  (.D(_0349_),
    .CLK(clknet_leaf_19_wr_clk),
    .Q(\mem[4][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][4]$_DFFE_PP_  (.D(_0350_),
    .CLK(clknet_leaf_17_wr_clk),
    .Q(\mem[4][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][5]$_DFFE_PP_  (.D(_0351_),
    .CLK(clknet_leaf_19_wr_clk),
    .Q(\mem[4][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][6]$_DFFE_PP_  (.D(_0352_),
    .CLK(clknet_leaf_15_wr_clk),
    .Q(\mem[4][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][7]$_DFFE_PP_  (.D(_0353_),
    .CLK(clknet_leaf_0_wr_clk),
    .Q(\mem[4][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][8]$_DFFE_PP_  (.D(_0354_),
    .CLK(clknet_leaf_15_wr_clk),
    .Q(\mem[4][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[4][9]$_DFFE_PP_  (.D(_0355_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[4][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][0]$_DFFE_PP_  (.D(_0356_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[5][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][10]$_DFFE_PP_  (.D(_0357_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[5][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][11]$_DFFE_PP_  (.D(_0358_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[5][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][12]$_DFFE_PP_  (.D(_0359_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[5][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][13]$_DFFE_PP_  (.D(_0360_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[5][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][14]$_DFFE_PP_  (.D(_0361_),
    .CLK(clknet_leaf_13_wr_clk),
    .Q(\mem[5][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][15]$_DFFE_PP_  (.D(_0362_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[5][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][16]$_DFFE_PP_  (.D(_0363_),
    .CLK(clknet_leaf_13_wr_clk),
    .Q(\mem[5][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][17]$_DFFE_PP_  (.D(_0364_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[5][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][18]$_DFFE_PP_  (.D(_0365_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[5][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][19]$_DFFE_PP_  (.D(_0366_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[5][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][1]$_DFFE_PP_  (.D(_0367_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[5][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][20]$_DFFE_PP_  (.D(_0368_),
    .CLK(clknet_leaf_6_wr_clk),
    .Q(\mem[5][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][21]$_DFFE_PP_  (.D(_0369_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[5][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][22]$_DFFE_PP_  (.D(_0370_),
    .CLK(clknet_leaf_6_wr_clk),
    .Q(\mem[5][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][23]$_DFFE_PP_  (.D(_0371_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[5][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][24]$_DFFE_PP_  (.D(_0372_),
    .CLK(clknet_leaf_2_wr_clk),
    .Q(\mem[5][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][25]$_DFFE_PP_  (.D(_0373_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[5][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][26]$_DFFE_PP_  (.D(_0374_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[5][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][27]$_DFFE_PP_  (.D(_0375_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[5][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][28]$_DFFE_PP_  (.D(_0376_),
    .CLK(clknet_leaf_17_wr_clk),
    .Q(\mem[5][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][29]$_DFFE_PP_  (.D(_0377_),
    .CLK(clknet_leaf_0_wr_clk),
    .Q(\mem[5][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][2]$_DFFE_PP_  (.D(_0378_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[5][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][30]$_DFFE_PP_  (.D(_0379_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[5][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][31]$_DFFE_PP_  (.D(_0380_),
    .CLK(clknet_leaf_0_wr_clk),
    .Q(\mem[5][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][3]$_DFFE_PP_  (.D(_0381_),
    .CLK(clknet_leaf_0_wr_clk),
    .Q(\mem[5][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][4]$_DFFE_PP_  (.D(_0382_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[5][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][5]$_DFFE_PP_  (.D(_0383_),
    .CLK(clknet_leaf_0_wr_clk),
    .Q(\mem[5][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][6]$_DFFE_PP_  (.D(_0384_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[5][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][7]$_DFFE_PP_  (.D(_0385_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[5][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][8]$_DFFE_PP_  (.D(_0386_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[5][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[5][9]$_DFFE_PP_  (.D(_0387_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[5][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][0]$_DFFE_PP_  (.D(_0388_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[6][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][10]$_DFFE_PP_  (.D(_0389_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[6][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][11]$_DFFE_PP_  (.D(_0390_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[6][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][12]$_DFFE_PP_  (.D(_0391_),
    .CLK(clknet_leaf_13_wr_clk),
    .Q(\mem[6][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][13]$_DFFE_PP_  (.D(_0392_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[6][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][14]$_DFFE_PP_  (.D(_0393_),
    .CLK(clknet_leaf_13_wr_clk),
    .Q(\mem[6][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][15]$_DFFE_PP_  (.D(_0394_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[6][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][16]$_DFFE_PP_  (.D(_0395_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[6][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][17]$_DFFE_PP_  (.D(_0396_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[6][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][18]$_DFFE_PP_  (.D(_0397_),
    .CLK(clknet_leaf_10_wr_clk),
    .Q(\mem[6][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][19]$_DFFE_PP_  (.D(_0398_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[6][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][1]$_DFFE_PP_  (.D(_0399_),
    .CLK(clknet_leaf_4_wr_clk),
    .Q(\mem[6][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][20]$_DFFE_PP_  (.D(_0400_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[6][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][21]$_DFFE_PP_  (.D(_0401_),
    .CLK(clknet_leaf_4_wr_clk),
    .Q(\mem[6][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][22]$_DFFE_PP_  (.D(_0402_),
    .CLK(clknet_leaf_6_wr_clk),
    .Q(\mem[6][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][23]$_DFFE_PP_  (.D(_0403_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[6][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][24]$_DFFE_PP_  (.D(_0404_),
    .CLK(clknet_leaf_2_wr_clk),
    .Q(\mem[6][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][25]$_DFFE_PP_  (.D(_0405_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[6][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][26]$_DFFE_PP_  (.D(_0406_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[6][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][27]$_DFFE_PP_  (.D(_0407_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[6][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][28]$_DFFE_PP_  (.D(_0408_),
    .CLK(clknet_leaf_18_wr_clk),
    .Q(\mem[6][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][29]$_DFFE_PP_  (.D(_0409_),
    .CLK(clknet_leaf_0_wr_clk),
    .Q(\mem[6][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][2]$_DFFE_PP_  (.D(_0410_),
    .CLK(clknet_leaf_17_wr_clk),
    .Q(\mem[6][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][30]$_DFFE_PP_  (.D(_0411_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[6][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][31]$_DFFE_PP_  (.D(_0412_),
    .CLK(clknet_leaf_19_wr_clk),
    .Q(\mem[6][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][3]$_DFFE_PP_  (.D(_0413_),
    .CLK(clknet_leaf_19_wr_clk),
    .Q(\mem[6][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][4]$_DFFE_PP_  (.D(_0414_),
    .CLK(clknet_leaf_17_wr_clk),
    .Q(\mem[6][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][5]$_DFFE_PP_  (.D(_0415_),
    .CLK(clknet_leaf_19_wr_clk),
    .Q(\mem[6][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][6]$_DFFE_PP_  (.D(_0416_),
    .CLK(clknet_leaf_15_wr_clk),
    .Q(\mem[6][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][7]$_DFFE_PP_  (.D(_0417_),
    .CLK(clknet_leaf_0_wr_clk),
    .Q(\mem[6][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][8]$_DFFE_PP_  (.D(_0418_),
    .CLK(clknet_leaf_15_wr_clk),
    .Q(\mem[6][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[6][9]$_DFFE_PP_  (.D(_0419_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[6][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][0]$_DFFE_PP_  (.D(_0420_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[7][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][10]$_DFFE_PP_  (.D(_0421_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[7][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][11]$_DFFE_PP_  (.D(_0422_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[7][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][12]$_DFFE_PP_  (.D(_0423_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[7][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][13]$_DFFE_PP_  (.D(_0424_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[7][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][14]$_DFFE_PP_  (.D(_0425_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[7][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][15]$_DFFE_PP_  (.D(_0426_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[7][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][16]$_DFFE_PP_  (.D(_0427_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[7][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][17]$_DFFE_PP_  (.D(_0428_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[7][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][18]$_DFFE_PP_  (.D(_0429_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[7][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][19]$_DFFE_PP_  (.D(_0430_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[7][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][1]$_DFFE_PP_  (.D(_0431_),
    .CLK(clknet_leaf_4_wr_clk),
    .Q(\mem[7][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][20]$_DFFE_PP_  (.D(_0432_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[7][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][21]$_DFFE_PP_  (.D(_0433_),
    .CLK(clknet_leaf_4_wr_clk),
    .Q(\mem[7][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][22]$_DFFE_PP_  (.D(_0434_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[7][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][23]$_DFFE_PP_  (.D(_0435_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[7][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][24]$_DFFE_PP_  (.D(_0436_),
    .CLK(clknet_leaf_6_wr_clk),
    .Q(\mem[7][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][25]$_DFFE_PP_  (.D(_0437_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[7][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][26]$_DFFE_PP_  (.D(_0438_),
    .CLK(clknet_leaf_2_wr_clk),
    .Q(\mem[7][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][27]$_DFFE_PP_  (.D(_0439_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[7][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][28]$_DFFE_PP_  (.D(_0440_),
    .CLK(clknet_leaf_17_wr_clk),
    .Q(\mem[7][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][29]$_DFFE_PP_  (.D(_0441_),
    .CLK(clknet_leaf_0_wr_clk),
    .Q(\mem[7][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][2]$_DFFE_PP_  (.D(_0442_),
    .CLK(clknet_leaf_17_wr_clk),
    .Q(\mem[7][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][30]$_DFFE_PP_  (.D(_0443_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[7][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][31]$_DFFE_PP_  (.D(_0444_),
    .CLK(clknet_leaf_0_wr_clk),
    .Q(\mem[7][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][3]$_DFFE_PP_  (.D(_0445_),
    .CLK(clknet_leaf_19_wr_clk),
    .Q(\mem[7][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][4]$_DFFE_PP_  (.D(_0446_),
    .CLK(clknet_leaf_17_wr_clk),
    .Q(\mem[7][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][5]$_DFFE_PP_  (.D(_0447_),
    .CLK(clknet_leaf_19_wr_clk),
    .Q(\mem[7][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][6]$_DFFE_PP_  (.D(_0448_),
    .CLK(clknet_leaf_15_wr_clk),
    .Q(\mem[7][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][7]$_DFFE_PP_  (.D(_0449_),
    .CLK(clknet_leaf_0_wr_clk),
    .Q(\mem[7][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][8]$_DFFE_PP_  (.D(_0450_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[7][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[7][9]$_DFFE_PP_  (.D(_0451_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[7][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][0]$_DFFE_PP_  (.D(_0452_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[8][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][10]$_DFFE_PP_  (.D(_0453_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[8][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][11]$_DFFE_PP_  (.D(_0454_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[8][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][12]$_DFFE_PP_  (.D(_0455_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[8][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][13]$_DFFE_PP_  (.D(_0456_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[8][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][14]$_DFFE_PP_  (.D(_0457_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[8][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][15]$_DFFE_PP_  (.D(_0458_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[8][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][16]$_DFFE_PP_  (.D(_0459_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[8][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][17]$_DFFE_PP_  (.D(_0460_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[8][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][18]$_DFFE_PP_  (.D(_0461_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[8][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][19]$_DFFE_PP_  (.D(_0462_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[8][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][1]$_DFFE_PP_  (.D(_0463_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[8][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][20]$_DFFE_PP_  (.D(_0464_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[8][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][21]$_DFFE_PP_  (.D(_0465_),
    .CLK(clknet_leaf_4_wr_clk),
    .Q(\mem[8][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][22]$_DFFE_PP_  (.D(_0466_),
    .CLK(clknet_leaf_6_wr_clk),
    .Q(\mem[8][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][23]$_DFFE_PP_  (.D(_0467_),
    .CLK(clknet_leaf_4_wr_clk),
    .Q(\mem[8][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][24]$_DFFE_PP_  (.D(_0468_),
    .CLK(clknet_leaf_2_wr_clk),
    .Q(\mem[8][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][25]$_DFFE_PP_  (.D(_0469_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[8][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][26]$_DFFE_PP_  (.D(_0470_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[8][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][27]$_DFFE_PP_  (.D(_0471_),
    .CLK(clknet_leaf_2_wr_clk),
    .Q(\mem[8][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][28]$_DFFE_PP_  (.D(_0472_),
    .CLK(clknet_leaf_18_wr_clk),
    .Q(\mem[8][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][29]$_DFFE_PP_  (.D(_0473_),
    .CLK(clknet_leaf_0_wr_clk),
    .Q(\mem[8][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][2]$_DFFE_PP_  (.D(_0474_),
    .CLK(clknet_leaf_17_wr_clk),
    .Q(\mem[8][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][30]$_DFFE_PP_  (.D(_0475_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[8][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][31]$_DFFE_PP_  (.D(_0476_),
    .CLK(clknet_leaf_0_wr_clk),
    .Q(\mem[8][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][3]$_DFFE_PP_  (.D(_0477_),
    .CLK(clknet_leaf_19_wr_clk),
    .Q(\mem[8][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][4]$_DFFE_PP_  (.D(_0478_),
    .CLK(clknet_leaf_17_wr_clk),
    .Q(\mem[8][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][5]$_DFFE_PP_  (.D(_0479_),
    .CLK(clknet_leaf_19_wr_clk),
    .Q(\mem[8][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][6]$_DFFE_PP_  (.D(_0480_),
    .CLK(clknet_leaf_15_wr_clk),
    .Q(\mem[8][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][7]$_DFFE_PP_  (.D(_0481_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[8][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][8]$_DFFE_PP_  (.D(_0482_),
    .CLK(clknet_leaf_15_wr_clk),
    .Q(\mem[8][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[8][9]$_DFFE_PP_  (.D(_0483_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[8][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][0]$_DFFE_PP_  (.D(_0484_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[9][0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][10]$_DFFE_PP_  (.D(_0485_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[9][10] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][11]$_DFFE_PP_  (.D(_0486_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[9][11] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][12]$_DFFE_PP_  (.D(_0487_),
    .CLK(clknet_leaf_11_wr_clk),
    .Q(\mem[9][12] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][13]$_DFFE_PP_  (.D(_0488_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[9][13] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][14]$_DFFE_PP_  (.D(_0489_),
    .CLK(clknet_leaf_13_wr_clk),
    .Q(\mem[9][14] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][15]$_DFFE_PP_  (.D(_0490_),
    .CLK(clknet_leaf_9_wr_clk),
    .Q(\mem[9][15] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][16]$_DFFE_PP_  (.D(_0491_),
    .CLK(clknet_leaf_12_wr_clk),
    .Q(\mem[9][16] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][17]$_DFFE_PP_  (.D(_0492_),
    .CLK(clknet_leaf_8_wr_clk),
    .Q(\mem[9][17] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][18]$_DFFE_PP_  (.D(_0493_),
    .CLK(clknet_leaf_7_wr_clk),
    .Q(\mem[9][18] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][19]$_DFFE_PP_  (.D(_0494_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[9][19] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][1]$_DFFE_PP_  (.D(_0495_),
    .CLK(clknet_leaf_5_wr_clk),
    .Q(\mem[9][1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][20]$_DFFE_PP_  (.D(_0496_),
    .CLK(clknet_leaf_6_wr_clk),
    .Q(\mem[9][20] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][21]$_DFFE_PP_  (.D(_0497_),
    .CLK(clknet_leaf_4_wr_clk),
    .Q(\mem[9][21] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][22]$_DFFE_PP_  (.D(_0498_),
    .CLK(clknet_leaf_6_wr_clk),
    .Q(\mem[9][22] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][23]$_DFFE_PP_  (.D(_0499_),
    .CLK(clknet_leaf_4_wr_clk),
    .Q(\mem[9][23] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][24]$_DFFE_PP_  (.D(_0500_),
    .CLK(clknet_leaf_2_wr_clk),
    .Q(\mem[9][24] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][25]$_DFFE_PP_  (.D(_0501_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[9][25] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][26]$_DFFE_PP_  (.D(_0502_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[9][26] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][27]$_DFFE_PP_  (.D(_0503_),
    .CLK(clknet_leaf_3_wr_clk),
    .Q(\mem[9][27] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][28]$_DFFE_PP_  (.D(_0504_),
    .CLK(clknet_leaf_17_wr_clk),
    .Q(\mem[9][28] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][29]$_DFFE_PP_  (.D(_0505_),
    .CLK(clknet_leaf_0_wr_clk),
    .Q(\mem[9][29] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][2]$_DFFE_PP_  (.D(_0506_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[9][2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][30]$_DFFE_PP_  (.D(_0507_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[9][30] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][31]$_DFFE_PP_  (.D(_0508_),
    .CLK(clknet_leaf_0_wr_clk),
    .Q(\mem[9][31] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][3]$_DFFE_PP_  (.D(_0509_),
    .CLK(clknet_leaf_19_wr_clk),
    .Q(\mem[9][3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][4]$_DFFE_PP_  (.D(_0510_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[9][4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][5]$_DFFE_PP_  (.D(_0511_),
    .CLK(clknet_leaf_19_wr_clk),
    .Q(\mem[9][5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][6]$_DFFE_PP_  (.D(_0512_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[9][6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][7]$_DFFE_PP_  (.D(_0513_),
    .CLK(clknet_leaf_1_wr_clk),
    .Q(\mem[9][7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][8]$_DFFE_PP_  (.D(_0514_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[9][8] ));
 gf180mcu_fd_sc_mcu9t5v0__dffq_2 \mem[9][9]$_DFFE_PP_  (.D(_0515_),
    .CLK(clknet_leaf_16_wr_clk),
    .Q(\mem[9][9] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[0]$_DFFE_PN0P_  (.D(_0516_),
    .RN(net4),
    .CLK(net2),
    .Q(net45));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[10]$_DFFE_PN0P_  (.D(_0517_),
    .RN(net4),
    .CLK(net2),
    .Q(net46));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[11]$_DFFE_PN0P_  (.D(_0518_),
    .RN(net4),
    .CLK(net2),
    .Q(net47));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[12]$_DFFE_PN0P_  (.D(_0519_),
    .RN(net4),
    .CLK(net2),
    .Q(net48));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[13]$_DFFE_PN0P_  (.D(_0520_),
    .RN(net4),
    .CLK(net2),
    .Q(net49));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[14]$_DFFE_PN0P_  (.D(_0521_),
    .RN(net4),
    .CLK(net2),
    .Q(net50));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[15]$_DFFE_PN0P_  (.D(_0522_),
    .RN(net4),
    .CLK(net2),
    .Q(net51));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[16]$_DFFE_PN0P_  (.D(_0523_),
    .RN(net4),
    .CLK(net2),
    .Q(net52));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[17]$_DFFE_PN0P_  (.D(_0524_),
    .RN(net4),
    .CLK(net2),
    .Q(net53));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[18]$_DFFE_PN0P_  (.D(_0525_),
    .RN(net4),
    .CLK(net2),
    .Q(net54));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[19]$_DFFE_PN0P_  (.D(_0526_),
    .RN(net4),
    .CLK(net2),
    .Q(net55));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[1]$_DFFE_PN0P_  (.D(_0527_),
    .RN(net4),
    .CLK(net2),
    .Q(net56));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[20]$_DFFE_PN0P_  (.D(_0528_),
    .RN(net4),
    .CLK(net2),
    .Q(net57));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[21]$_DFFE_PN0P_  (.D(_0529_),
    .RN(net4),
    .CLK(net2),
    .Q(net58));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[22]$_DFFE_PN0P_  (.D(_0530_),
    .RN(net4),
    .CLK(net2),
    .Q(net59));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[23]$_DFFE_PN0P_  (.D(_0531_),
    .RN(net4),
    .CLK(net2),
    .Q(net60));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[24]$_DFFE_PN0P_  (.D(_0532_),
    .RN(net4),
    .CLK(net2),
    .Q(net61));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[25]$_DFFE_PN0P_  (.D(_0533_),
    .RN(net4),
    .CLK(net2),
    .Q(net62));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[26]$_DFFE_PN0P_  (.D(_0534_),
    .RN(net4),
    .CLK(net2),
    .Q(net63));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[27]$_DFFE_PN0P_  (.D(_0535_),
    .RN(net4),
    .CLK(net2),
    .Q(net64));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[28]$_DFFE_PN0P_  (.D(_0536_),
    .RN(net4),
    .CLK(net2),
    .Q(net65));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[29]$_DFFE_PN0P_  (.D(_0537_),
    .RN(net4),
    .CLK(net2),
    .Q(net66));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[2]$_DFFE_PN0P_  (.D(_0538_),
    .RN(net4),
    .CLK(net2),
    .Q(net67));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[30]$_DFFE_PN0P_  (.D(_0539_),
    .RN(net4),
    .CLK(net2),
    .Q(net68));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[31]$_DFFE_PN0P_  (.D(_0540_),
    .RN(net4),
    .CLK(net2),
    .Q(net69));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[3]$_DFFE_PN0P_  (.D(_0541_),
    .RN(net4),
    .CLK(net2),
    .Q(net70));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[4]$_DFFE_PN0P_  (.D(_0542_),
    .RN(net4),
    .CLK(net2),
    .Q(net71));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[5]$_DFFE_PN0P_  (.D(_0543_),
    .RN(net4),
    .CLK(net2),
    .Q(net72));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[6]$_DFFE_PN0P_  (.D(_0544_),
    .RN(net4),
    .CLK(net2),
    .Q(net73));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[7]$_DFFE_PN0P_  (.D(_0545_),
    .RN(net4),
    .CLK(net2),
    .Q(net74));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[8]$_DFFE_PN0P_  (.D(_0546_),
    .RN(net4),
    .CLK(net2),
    .Q(net75));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_data[9]$_DFFE_PN0P_  (.D(_0547_),
    .RN(net4),
    .CLK(net2),
    .Q(net76));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_ptr_bin[0]$_DFFE_PN0P_  (.D(_0548_),
    .RN(net4),
    .CLK(net2),
    .Q(\rd_ptr_bin[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_ptr_bin[1]$_DFFE_PN0P_  (.D(_0549_),
    .RN(net4),
    .CLK(net2),
    .Q(\rd_ptr_bin[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_ptr_bin[2]$_DFFE_PN0P_  (.D(_0550_),
    .RN(net4),
    .CLK(net2),
    .Q(\rd_ptr_bin[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \rd_ptr_bin[3]$_DFFE_PN0P_  (.D(_0551_),
    .RN(net4),
    .CLK(net2),
    .Q(\rd_ptr_bin[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_ptr_gray[0]$_DFFE_PN0P_  (.D(_0552_),
    .RN(net4),
    .CLK(net2),
    .Q(\rd_ptr_gray[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_ptr_gray[1]$_DFFE_PN0P_  (.D(_0553_),
    .RN(net4),
    .CLK(net2),
    .Q(\rd_ptr_gray[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_ptr_gray[2]$_DFFE_PN0P_  (.D(_0554_),
    .RN(net4),
    .CLK(net2),
    .Q(\rd_ptr_gray[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_ptr_gray[3]$_DFFE_PN0P_  (.D(_0555_),
    .RN(net4),
    .CLK(net2),
    .Q(\rd_ptr_gray[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_ptr_gray[4]$_DFFE_PN0P_  (.D(_0556_),
    .RN(net4),
    .CLK(net2),
    .Q(\rd_ptr_bin[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_ptr_gray_sync1[0]$_DFF_PN0_  (.D(\rd_ptr_gray[0] ),
    .RN(net1),
    .CLK(clknet_leaf_14_wr_clk),
    .Q(\rd_ptr_gray_sync1[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_ptr_gray_sync1[1]$_DFF_PN0_  (.D(\rd_ptr_gray[1] ),
    .RN(net1),
    .CLK(clknet_leaf_14_wr_clk),
    .Q(\rd_ptr_gray_sync1[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_ptr_gray_sync1[2]$_DFF_PN0_  (.D(\rd_ptr_gray[2] ),
    .RN(net1),
    .CLK(clknet_leaf_14_wr_clk),
    .Q(\rd_ptr_gray_sync1[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_ptr_gray_sync1[3]$_DFF_PN0_  (.D(\rd_ptr_gray[3] ),
    .RN(net1),
    .CLK(clknet_leaf_14_wr_clk),
    .Q(\rd_ptr_gray_sync1[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_ptr_gray_sync1[4]$_DFF_PN0_  (.D(\rd_ptr_bin[4] ),
    .RN(net1),
    .CLK(clknet_leaf_14_wr_clk),
    .Q(\rd_ptr_gray_sync1[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_ptr_gray_sync2[0]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[0] ),
    .RN(net1),
    .CLK(clknet_leaf_14_wr_clk),
    .Q(\rd_ptr_gray_sync2[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_ptr_gray_sync2[1]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[1] ),
    .RN(net1),
    .CLK(clknet_leaf_14_wr_clk),
    .Q(\rd_ptr_gray_sync2[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_ptr_gray_sync2[2]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[2] ),
    .RN(net1),
    .CLK(clknet_leaf_14_wr_clk),
    .Q(\rd_ptr_gray_sync2[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_ptr_gray_sync2[3]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[3] ),
    .RN(net1),
    .CLK(clknet_leaf_14_wr_clk),
    .Q(\rd_ptr_gray_sync2[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rd_ptr_gray_sync2[4]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[4] ),
    .RN(net1),
    .CLK(clknet_leaf_14_wr_clk),
    .Q(\rd_ptr_gray_sync2[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr_bin[0]$_DFFE_PN0P_  (.D(_0557_),
    .RN(net1),
    .CLK(clknet_leaf_14_wr_clk),
    .Q(\wr_ptr_bin[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr_bin[1]$_DFFE_PN0P_  (.D(_0558_),
    .RN(net1),
    .CLK(clknet_leaf_14_wr_clk),
    .Q(\wr_ptr_bin[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr_bin[2]$_DFFE_PN0P_  (.D(_0559_),
    .RN(net1),
    .CLK(clknet_leaf_14_wr_clk),
    .Q(\wr_ptr_bin[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr_bin[3]$_DFFE_PN0P_  (.D(_0560_),
    .RN(net1),
    .CLK(clknet_leaf_14_wr_clk),
    .Q(\wr_ptr_bin[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr_gray[0]$_DFFE_PN0P_  (.D(_0561_),
    .RN(net1),
    .CLK(clknet_leaf_14_wr_clk),
    .Q(\wr_ptr_gray[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr_gray[1]$_DFFE_PN0P_  (.D(_0562_),
    .RN(net1),
    .CLK(clknet_leaf_14_wr_clk),
    .Q(\wr_ptr_gray[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr_gray[2]$_DFFE_PN0P_  (.D(_0563_),
    .RN(net1),
    .CLK(clknet_leaf_14_wr_clk),
    .Q(\wr_ptr_gray[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr_gray[3]$_DFFE_PN0P_  (.D(_0564_),
    .RN(net1),
    .CLK(clknet_leaf_14_wr_clk),
    .Q(\wr_ptr_gray[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr_gray[4]$_DFFE_PN0P_  (.D(_0565_),
    .RN(net1),
    .CLK(clknet_leaf_14_wr_clk),
    .Q(\wr_ptr_bin[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr_gray_sync1[0]$_DFF_PN0_  (.D(\wr_ptr_gray[0] ),
    .RN(net4),
    .CLK(net2),
    .Q(\wr_ptr_gray_sync1[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr_gray_sync1[1]$_DFF_PN0_  (.D(\wr_ptr_gray[1] ),
    .RN(net4),
    .CLK(net2),
    .Q(\wr_ptr_gray_sync1[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr_gray_sync1[2]$_DFF_PN0_  (.D(\wr_ptr_gray[2] ),
    .RN(net4),
    .CLK(net2),
    .Q(\wr_ptr_gray_sync1[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr_gray_sync1[3]$_DFF_PN0_  (.D(\wr_ptr_gray[3] ),
    .RN(net4),
    .CLK(net2),
    .Q(\wr_ptr_gray_sync1[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr_gray_sync1[4]$_DFF_PN0_  (.D(\wr_ptr_bin[4] ),
    .RN(net4),
    .CLK(net2),
    .Q(\wr_ptr_gray_sync1[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr_gray_sync2[0]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[0] ),
    .RN(net4),
    .CLK(net2),
    .Q(\wr_ptr_gray_sync2[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr_gray_sync2[1]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[1] ),
    .RN(net4),
    .CLK(net2),
    .Q(\wr_ptr_gray_sync2[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr_gray_sync2[2]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[2] ),
    .RN(net4),
    .CLK(net2),
    .Q(\wr_ptr_gray_sync2[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr_gray_sync2[3]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[3] ),
    .RN(net4),
    .CLK(net2),
    .Q(\wr_ptr_gray_sync2[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \wr_ptr_gray_sync2[4]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[4] ),
    .RN(net4),
    .CLK(net2),
    .Q(\wr_ptr_gray_sync2[4] ));
 gf180mcu_fd_sc_mcu9t5v0__buf_8 hold1 (.I(net38),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_103 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_104 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_105 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_106 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_107 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_108 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_109 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_110 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_111 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_112 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_113 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_114 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_115 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_116 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_117 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_118 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_119 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_120 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_121 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_122 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_123 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_124 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_125 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_126 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_127 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_128 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_129 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_130 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_131 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_132 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_133 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_134 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_135 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_136 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_137 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_138 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_139 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_140 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_141 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_142 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_143 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_144 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Left_145 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Left_146 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Left_147 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Left_148 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Left_149 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Left_150 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Left_151 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Left_152 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Left_153 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Left_154 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Left_155 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Left_156 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Left_157 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Left_158 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Left_159 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Left_160 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Left_161 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Left_162 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Left_163 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Left_164 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Left_165 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Left_166 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Left_167 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_65_Left_168 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_66_Left_169 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_67_Left_170 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_68_Left_171 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_69_Left_172 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_70_Left_173 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_71_Left_174 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_72_Left_175 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_73_Left_176 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_74_Left_177 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_75_Left_178 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_76_Left_179 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_77_Left_180 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_78_Left_181 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_79_Left_182 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_80_Left_183 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_81_Left_184 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_82_Left_185 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_83_Left_186 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_84_Left_187 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_85_Left_188 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_86_Left_189 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_87_Left_190 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_88_Left_191 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_89_Left_192 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_90_Left_193 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_91_Left_194 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_92_Left_195 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_93_Left_196 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_94_Left_197 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_95_Left_198 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_96_Left_199 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_97_Left_200 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_98_Left_201 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_99_Left_202 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_100_Left_203 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_101_Left_204 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_102_Left_205 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_206 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_207 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_208 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_209 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_210 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_211 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_212 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_213 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_214 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_215 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_216 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_217 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_218 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_219 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_220 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_221 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_222 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_223 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_224 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_225 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_226 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_227 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_228 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_229 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_230 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_231 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_232 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_233 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_234 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_235 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_236 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_237 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_238 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_239 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_240 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_241 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_242 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_243 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_244 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_245 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_246 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_247 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_248 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_249 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_250 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_251 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_252 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_253 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_254 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_255 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_256 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_257 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_258 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_259 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_260 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_261 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_262 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_263 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_264 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_265 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_266 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_267 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_268 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_269 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_270 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_271 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_272 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_273 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_274 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_275 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_276 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_277 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_278 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_279 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_280 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_281 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_282 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_283 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_284 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_285 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_286 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_287 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_288 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_289 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_290 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_291 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_292 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_293 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_294 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_295 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_296 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_297 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_298 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_299 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_300 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_301 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_302 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_303 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_304 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_305 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_306 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_307 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_308 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_309 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_310 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_311 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_312 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_313 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_314 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_315 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_316 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_317 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_318 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_319 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_320 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_321 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_322 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_323 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_324 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_325 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_326 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_327 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_328 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_329 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_330 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_331 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_332 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_333 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_334 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_335 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_336 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_337 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_338 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_339 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_340 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_341 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_342 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_343 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_344 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_345 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_346 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_347 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_348 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_349 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_350 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_351 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_352 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_353 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_354 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_355 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_356 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_357 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_358 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_359 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_360 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_361 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_362 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_363 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_364 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_365 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_366 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_367 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_368 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_369 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_370 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_371 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_65_372 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_373 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_374 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_66_375 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_376 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_67_377 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_378 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_379 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_68_380 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_381 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_69_382 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_383 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_384 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_70_385 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_386 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_71_387 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_388 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_389 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_72_390 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_391 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_73_392 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_393 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_394 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_74_395 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_396 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_75_397 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_398 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_399 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_76_400 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_401 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_77_402 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_403 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_404 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_78_405 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_406 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_79_407 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_408 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_409 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_80_410 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_411 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_81_412 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_413 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_414 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_82_415 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_416 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_83_417 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_418 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_419 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_84_420 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_421 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_85_422 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_423 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_424 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_86_425 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_426 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_87_427 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_428 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_429 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_88_430 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_431 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_89_432 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_433 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_434 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_90_435 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_436 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_91_437 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_438 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_439 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_92_440 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_441 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_93_442 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_443 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_444 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_94_445 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_446 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_95_447 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_448 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_449 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_96_450 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_451 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_97_452 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_453 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_454 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_98_455 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_456 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_99_457 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_458 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_459 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_100_460 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_461 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_101_462 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_463 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_464 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_465 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_466 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_102_467 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_16 input1 (.I(rd_clk),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input2 (.I(rd_en),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__buf_20 input3 (.I(rd_rst_n),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input4 (.I(net113),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input5 (.I(net103),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input6 (.I(net89),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input7 (.I(net105),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input8 (.I(net87),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input9 (.I(net96),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input10 (.I(net97),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input11 (.I(net104),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input12 (.I(net100),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input13 (.I(net116),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input14 (.I(net90),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input15 (.I(net92),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input16 (.I(net107),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input17 (.I(net94),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input18 (.I(net110),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input19 (.I(net99),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input20 (.I(net115),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input21 (.I(net88),
    .Z(net22));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input22 (.I(net114),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input23 (.I(net86),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input24 (.I(net98),
    .Z(net25));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input25 (.I(net101),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input26 (.I(net93),
    .Z(net27));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input27 (.I(net117),
    .Z(net28));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input28 (.I(net91),
    .Z(net29));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input29 (.I(net109),
    .Z(net30));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input30 (.I(net95),
    .Z(net31));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input31 (.I(net111),
    .Z(net32));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input32 (.I(net108),
    .Z(net33));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input33 (.I(net102),
    .Z(net34));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input34 (.I(net112),
    .Z(net35));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 input35 (.I(net106),
    .Z(net36));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input36 (.I(wr_en),
    .Z(net37));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input37 (.I(net85),
    .Z(net38));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output38 (.I(net39),
    .Z(rd_almost_empty));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output39 (.I(net40),
    .Z(rd_count[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output40 (.I(net41),
    .Z(rd_count[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output41 (.I(net42),
    .Z(rd_count[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output42 (.I(net43),
    .Z(rd_count[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output43 (.I(net44),
    .Z(rd_count[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output44 (.I(net45),
    .Z(rd_data[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output45 (.I(net46),
    .Z(rd_data[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output46 (.I(net47),
    .Z(rd_data[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output47 (.I(net48),
    .Z(rd_data[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output48 (.I(net49),
    .Z(rd_data[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output49 (.I(net50),
    .Z(rd_data[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output50 (.I(net51),
    .Z(rd_data[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output51 (.I(net52),
    .Z(rd_data[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output52 (.I(net53),
    .Z(rd_data[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output53 (.I(net54),
    .Z(rd_data[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output54 (.I(net55),
    .Z(rd_data[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output55 (.I(net56),
    .Z(rd_data[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output56 (.I(net57),
    .Z(rd_data[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output57 (.I(net58),
    .Z(rd_data[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output58 (.I(net59),
    .Z(rd_data[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output59 (.I(net60),
    .Z(rd_data[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output60 (.I(net61),
    .Z(rd_data[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output61 (.I(net62),
    .Z(rd_data[25]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output62 (.I(net63),
    .Z(rd_data[26]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output63 (.I(net64),
    .Z(rd_data[27]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output64 (.I(net65),
    .Z(rd_data[28]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output65 (.I(net66),
    .Z(rd_data[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output66 (.I(net67),
    .Z(rd_data[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output67 (.I(net68),
    .Z(rd_data[30]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output68 (.I(net69),
    .Z(rd_data[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output69 (.I(net70),
    .Z(rd_data[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output70 (.I(net71),
    .Z(rd_data[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output71 (.I(net72),
    .Z(rd_data[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output72 (.I(net73),
    .Z(rd_data[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output73 (.I(net74),
    .Z(rd_data[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output74 (.I(net75),
    .Z(rd_data[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output75 (.I(net76),
    .Z(rd_data[9]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output76 (.I(net77),
    .Z(rd_empty));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output77 (.I(net78),
    .Z(wr_almost_full));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output78 (.I(net79),
    .Z(wr_count[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output79 (.I(net80),
    .Z(wr_count[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output80 (.I(net81),
    .Z(wr_count[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output81 (.I(net82),
    .Z(wr_count[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output82 (.I(net83),
    .Z(wr_count[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output83 (.I(net84),
    .Z(wr_full));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_0_wr_clk (.I(clknet_1_0__leaf_wr_clk),
    .Z(clknet_leaf_0_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_1_wr_clk (.I(clknet_1_0__leaf_wr_clk),
    .Z(clknet_leaf_1_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_2_wr_clk (.I(clknet_1_1__leaf_wr_clk),
    .Z(clknet_leaf_2_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_3_wr_clk (.I(clknet_1_1__leaf_wr_clk),
    .Z(clknet_leaf_3_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_4_wr_clk (.I(clknet_1_1__leaf_wr_clk),
    .Z(clknet_leaf_4_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_5_wr_clk (.I(clknet_1_1__leaf_wr_clk),
    .Z(clknet_leaf_5_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_6_wr_clk (.I(clknet_1_1__leaf_wr_clk),
    .Z(clknet_leaf_6_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_7_wr_clk (.I(clknet_1_1__leaf_wr_clk),
    .Z(clknet_leaf_7_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_8_wr_clk (.I(clknet_1_1__leaf_wr_clk),
    .Z(clknet_leaf_8_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_9_wr_clk (.I(clknet_1_1__leaf_wr_clk),
    .Z(clknet_leaf_9_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_10_wr_clk (.I(clknet_1_1__leaf_wr_clk),
    .Z(clknet_leaf_10_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_11_wr_clk (.I(clknet_1_1__leaf_wr_clk),
    .Z(clknet_leaf_11_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_12_wr_clk (.I(clknet_1_0__leaf_wr_clk),
    .Z(clknet_leaf_12_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_13_wr_clk (.I(clknet_1_0__leaf_wr_clk),
    .Z(clknet_leaf_13_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_14_wr_clk (.I(clknet_1_0__leaf_wr_clk),
    .Z(clknet_leaf_14_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_15_wr_clk (.I(clknet_1_0__leaf_wr_clk),
    .Z(clknet_leaf_15_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_16_wr_clk (.I(clknet_1_0__leaf_wr_clk),
    .Z(clknet_leaf_16_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_17_wr_clk (.I(clknet_1_0__leaf_wr_clk),
    .Z(clknet_leaf_17_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_18_wr_clk (.I(clknet_1_0__leaf_wr_clk),
    .Z(clknet_leaf_18_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 clkbuf_leaf_19_wr_clk (.I(clknet_1_0__leaf_wr_clk),
    .Z(clknet_leaf_19_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_0_wr_clk (.I(wr_clk),
    .Z(clknet_0_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_1_0__f_wr_clk (.I(clknet_0_wr_clk),
    .Z(clknet_1_0__leaf_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkbuf_1_1__f_wr_clk (.I(clknet_0_wr_clk),
    .Z(clknet_1_1__leaf_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload0 (.I(clknet_leaf_0_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 clkload1 (.I(clknet_leaf_1_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_1 clkload2 (.I(clknet_leaf_12_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_12 clkload3 (.I(clknet_leaf_13_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload4 (.I(clknet_leaf_14_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload5 (.I(clknet_leaf_15_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload6 (.I(clknet_leaf_17_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload7 (.I(clknet_leaf_18_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload8 (.I(clknet_leaf_19_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload9 (.I(clknet_leaf_2_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload10 (.I(clknet_leaf_3_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 clkload11 (.I(clknet_leaf_4_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload12 (.I(clknet_leaf_5_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 clkload13 (.I(clknet_leaf_6_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload14 (.I(clknet_leaf_8_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload15 (.I(clknet_leaf_9_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 clkload16 (.I(clknet_leaf_10_wr_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(wr_rst_n),
    .Z(net85));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold3 (.I(wr_data[27]),
    .Z(net86));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold4 (.I(wr_data[13]),
    .Z(net87));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold5 (.I(wr_data[25]),
    .Z(net88));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold6 (.I(wr_data[11]),
    .Z(net89));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold7 (.I(wr_data[19]),
    .Z(net90));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold8 (.I(wr_data[31]),
    .Z(net91));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold9 (.I(wr_data[1]),
    .Z(net92));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold10 (.I(wr_data[2]),
    .Z(net93));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold11 (.I(wr_data[21]),
    .Z(net94));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold12 (.I(wr_data[4]),
    .Z(net95));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold13 (.I(wr_data[14]),
    .Z(net96));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold14 (.I(wr_data[15]),
    .Z(net97));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold15 (.I(wr_data[28]),
    .Z(net98));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold16 (.I(wr_data[23]),
    .Z(net99));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold17 (.I(wr_data[17]),
    .Z(net100));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold18 (.I(wr_data[29]),
    .Z(net101));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold19 (.I(wr_data[7]),
    .Z(net102));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold20 (.I(wr_data[10]),
    .Z(net103));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold21 (.I(wr_data[16]),
    .Z(net104));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold22 (.I(wr_data[12]),
    .Z(net105));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold23 (.I(wr_data[9]),
    .Z(net106));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold24 (.I(wr_data[20]),
    .Z(net107));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold25 (.I(wr_data[6]),
    .Z(net108));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold26 (.I(wr_data[3]),
    .Z(net109));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold27 (.I(wr_data[22]),
    .Z(net110));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold28 (.I(wr_data[5]),
    .Z(net111));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold29 (.I(wr_data[8]),
    .Z(net112));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold30 (.I(wr_data[0]),
    .Z(net113));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold31 (.I(wr_data[26]),
    .Z(net114));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold32 (.I(wr_data[24]),
    .Z(net115));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold33 (.I(wr_data[18]),
    .Z(net116));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold34 (.I(wr_data[30]),
    .Z(net117));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_537 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_555 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_699 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_809 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_876 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_841 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_897 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_905 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_789 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_831 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_301 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_813 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_901 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_587 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_649 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_31_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_32_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_277 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_70 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_791 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_37_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_393 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_522 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_530 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_38_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_39_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_39_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_482 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_41_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_869 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_41_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_42_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_828 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_843 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_43_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_43_847 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_283 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_883 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_896 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_45_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_909 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_45_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_46_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_801 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_875 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_47_907 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_47_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_270 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_329 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_49_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_832 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_49_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_898 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_50_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_381 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_554 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_654 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_664 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_716 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_51_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_867 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_51_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_499 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_629 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_645 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_793 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_799 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_817 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_52_848 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_377 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_429 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_495 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_679 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_53_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_733 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_753 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_834 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_858 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_913 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_54_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_291 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_459 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_506 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_514 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_55_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_55_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_378 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_56_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_469 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_856 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_57_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_57_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_371 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_660 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_732 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_839 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_923 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_58_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_512 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_599 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_603 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_59_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_812 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_849 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_59_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_375 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_458 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_489 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_620 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_850 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_553 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_724 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_798 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_833 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_845 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_425 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_678 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_682 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_772 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_20 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_309 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_63_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_766 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_787 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_859 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_879 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_385 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_65_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_763 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_65_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_795 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_65_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_65_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_65_830 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_65_894 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_65_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_465 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_66_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_652 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_737 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_66_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_837 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_66_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_66_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_66_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_66_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_305 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_483 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_546 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_67_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_728 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_67_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_835 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_67_852 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_860 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_862 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_67_899 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_67_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_67_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_472 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_68_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_613 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_657 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_739 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_741 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_68_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_68_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_68_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_68_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_69_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_457 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_480 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_69_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_621 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_625 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_69_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_69_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_882 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_890 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_69_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_294 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_407 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_70_749 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_70_853 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_70_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_70_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_70_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_70_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_70_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_419 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_71_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_796 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_827 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_71_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_71_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_71_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_71_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_71_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_71_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_637 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_653 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_661 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_72_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_758 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_777 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_783 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_881 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_72_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_72_900 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_72_902 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_72_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_36 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_547 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_73_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_628 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_630 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_73_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_73_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_73_844 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_846 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_73_865 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_73_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_73_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_411 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_498 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_74_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_74_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_806 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_822 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_74_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_74_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_74_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_74_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_74_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_75_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_370 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_543 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_75_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_75_863 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_75_895 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_75_911 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_75_915 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_917 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_75_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_382 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_632 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_640 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_713 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_721 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_754 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_770 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_76_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_782 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_76_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_76_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_76_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_76_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_76_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_76_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_307 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_388 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_607 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_623 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_77_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_77_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_77_903 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_77_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_77_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_77_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_77_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_303 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_359 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_363 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_542 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_591 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_78_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_78_667 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_78_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_854 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_78_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_78_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_78_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_297 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_379 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_387 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_452 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_79_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_79_690 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_744 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_79_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_765 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_79_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_79_771 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_79_866 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_79_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_273 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_576 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_752 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_784 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_80_788 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_80_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_80_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_80_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_80_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_80_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_80_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_254 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_413 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_439 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_722 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_726 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_81_773 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_781 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_81_785 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_81_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_81_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_81_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_81_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_81_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_193 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_279 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_281 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_320 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_404 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_528 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_82_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_615 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_697 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_82_729 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_748 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_82_825 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_82_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_82_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_82_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_492 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_524 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_83_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_662 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_686 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_83_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_745 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_761 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_769 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_819 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_83_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_83_904 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_83_920 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_83_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_83_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_64 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_84_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_383 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_478 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_510 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_635 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_702 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_735 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_767 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_775 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_779 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_805 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_84_861 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_84_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_84_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_84_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_84_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_83 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_390 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_394 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_441 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_505 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_521 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_608 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_85_691 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_707 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_85_797 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_85_855 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_85_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_85_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_85_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_85_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_267 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_275 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_330 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_365 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_369 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_386 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_86_627 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_641 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_677 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_725 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_86_757 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_821 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_829 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_86_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_86_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_86_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_86_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_346 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_464 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_87_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_586 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_87_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_87_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_87_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_87_921 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_87_929 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_87_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_290 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_298 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_432 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_88_471 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_573 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_585 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_655 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_694 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_698 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_700 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_715 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_723 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_727 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_751 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_755 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_786 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_877 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_88_885 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_88_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_88_908 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_88_916 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_88_918 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_164 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_300 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_304 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_366 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_89_562 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_631 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_639 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_89_658 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_674 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_688 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_731 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_89_794 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_802 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_818 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_820 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_89_836 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_89_838 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_89_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_89_870 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_136 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_90_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_367 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_442 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_90_461 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_571 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_575 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_618 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_626 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_644 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_663 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_671 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_675 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_685 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_693 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_695 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_803 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_90_811 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_857 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_90_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_90_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_90_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_285 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_317 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_319 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_364 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_418 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_437 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_445 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_91_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_511 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_656 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_672 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_705 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_91_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_740 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_91_816 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_91_880 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_91_912 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_91_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_91_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_29 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_280 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_288 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_332 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_356 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_362 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_408 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_424 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_497 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_501 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_503 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_545 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_549 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_92_551 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_614 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_692 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_756 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_764 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_768 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_92_804 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_92_868 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_92_884 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_92_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_92_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_92_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_30 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_257 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_296 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_328 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_405 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_466 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_477 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_624 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_650 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_666 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_93_710 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_93_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_93_734 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_750 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_93_814 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_93_878 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_93_910 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_93_926 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_454 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_515 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_94_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_670 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_94_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_717 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_94_719 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_760 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_94_824 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_94_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_94_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_94_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_271 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_306 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_323 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_343 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_376 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_403 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_435 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_484 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_488 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_490 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_516 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_520 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_609 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_95_642 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_759 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_95_823 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_95_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_95_919 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_95_927 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_95_931 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_95_933 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_314 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_395 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_399 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_401 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_451 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_467 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_475 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_597 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_96_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_647 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_681 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_96_704 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_738 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_96_776 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_840 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_96_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_96_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_96_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_96_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_97_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_402 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_410 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_414 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_446 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_97_474 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_494 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_601 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_97_617 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_648 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_778 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_97_842 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_97_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_97_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_268 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_315 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_368 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_400 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_416 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_450 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_509 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_525 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_98_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_566 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_583 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_600 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_604 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_651 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_98_683 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_98_689 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_706 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_762 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_98_826 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_98_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_98_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_98_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_278 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_295 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_327 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_335 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_339 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_341 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_444 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_508 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_556 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_596 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_616 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_633 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_665 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_669 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_701 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_99_730 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_746 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_99_810 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_99_874 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_99_906 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_99_930 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_340 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_360 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_396 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_476 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_507 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_523 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_598 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_606 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_610 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_612 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_643 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_659 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_100_708 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_712 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_743 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_100_807 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_100_871 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_887 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_100_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_100_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_100_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_292 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_326 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_406 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_430 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_434 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_443 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_447 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_463 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_535 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_539 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_541 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_557 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_579 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_611 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_619 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_101_636 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_668 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_101_687 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_101_703 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_711 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_101_720 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_736 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_800 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_101_864 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_101_928 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_101_932 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_380 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_384 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_427 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_473 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_540 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_572 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_588 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_622 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_638 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_646 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_680 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_696 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_102_714 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_718 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_742 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_774 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_790 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_102_792 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_102_808 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_102_872 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_888 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_102_892 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_102_924 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_102_932 ();
endmodule
