module network_interface_cdc (dst_clk,
    dst_rst_n,
    mem_read,
    mem_ready,
    mem_write,
    router_in_ready,
    router_in_valid,
    router_out_ready,
    router_out_valid,
    src_clk,
    src_rst_n,
    dest_id,
    mem_addr,
    mem_rdata,
    mem_wdata,
    msg_type,
    router_in_data,
    router_out_data);
 input dst_clk;
 input dst_rst_n;
 input mem_read;
 output mem_ready;
 input mem_write;
 input router_in_ready;
 output router_in_valid;
 output router_out_ready;
 input router_out_valid;
 input src_clk;
 input src_rst_n;
 input [7:0] dest_id;
 input [31:0] mem_addr;
 output [31:0] mem_rdata;
 input [31:0] mem_wdata;
 input [2:0] msg_type;
 output [31:0] router_in_data;
 input [31:0] router_out_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire dst_ack;
 wire dst_ack_prev;
 wire dst_ack_sync;
 wire \dst_ack_sync_reg[0] ;
 wire dst_data_valid;
 wire dst_data_valid_sync;
 wire \dst_data_valid_sync_reg[0] ;
 wire dst_is_write_op;
 wire \dst_state[0] ;
 wire \dst_state[1] ;
 wire \dst_state[2] ;
 wire \dst_state[3] ;
 wire \dst_to_src_data[0] ;
 wire \dst_to_src_data[10] ;
 wire \dst_to_src_data[11] ;
 wire \dst_to_src_data[12] ;
 wire \dst_to_src_data[13] ;
 wire \dst_to_src_data[14] ;
 wire \dst_to_src_data[15] ;
 wire \dst_to_src_data[16] ;
 wire \dst_to_src_data[17] ;
 wire \dst_to_src_data[18] ;
 wire \dst_to_src_data[19] ;
 wire \dst_to_src_data[1] ;
 wire \dst_to_src_data[20] ;
 wire \dst_to_src_data[21] ;
 wire \dst_to_src_data[22] ;
 wire \dst_to_src_data[23] ;
 wire \dst_to_src_data[24] ;
 wire \dst_to_src_data[25] ;
 wire \dst_to_src_data[26] ;
 wire \dst_to_src_data[27] ;
 wire \dst_to_src_data[28] ;
 wire \dst_to_src_data[29] ;
 wire \dst_to_src_data[2] ;
 wire \dst_to_src_data[30] ;
 wire \dst_to_src_data[31] ;
 wire \dst_to_src_data[3] ;
 wire \dst_to_src_data[4] ;
 wire \dst_to_src_data[5] ;
 wire \dst_to_src_data[6] ;
 wire \dst_to_src_data[7] ;
 wire \dst_to_src_data[8] ;
 wire \dst_to_src_data[9] ;
 wire src_data_valid;
 wire src_data_valid_sync;
 wire \src_data_valid_sync_reg[0] ;
 wire src_is_write_op_flag;
 wire src_is_write_op_sync;
 wire \src_is_write_op_sync_reg[0] ;
 wire src_req;
 wire src_req_prev;
 wire src_req_sync;
 wire \src_req_sync_reg[0] ;
 wire \src_state[0] ;
 wire \src_state[1] ;
 wire \src_state[2] ;
 wire \src_state[3] ;
 wire \src_to_dst_data[0] ;
 wire \src_to_dst_data[10] ;
 wire \src_to_dst_data[11] ;
 wire \src_to_dst_data[12] ;
 wire \src_to_dst_data[13] ;
 wire \src_to_dst_data[14] ;
 wire \src_to_dst_data[15] ;
 wire \src_to_dst_data[16] ;
 wire \src_to_dst_data[17] ;
 wire \src_to_dst_data[18] ;
 wire \src_to_dst_data[19] ;
 wire \src_to_dst_data[1] ;
 wire \src_to_dst_data[20] ;
 wire \src_to_dst_data[21] ;
 wire \src_to_dst_data[22] ;
 wire \src_to_dst_data[23] ;
 wire \src_to_dst_data[24] ;
 wire \src_to_dst_data[25] ;
 wire \src_to_dst_data[26] ;
 wire \src_to_dst_data[27] ;
 wire \src_to_dst_data[28] ;
 wire \src_to_dst_data[29] ;
 wire \src_to_dst_data[2] ;
 wire \src_to_dst_data[30] ;
 wire \src_to_dst_data[31] ;
 wire \src_to_dst_data[3] ;
 wire \src_to_dst_data[4] ;
 wire \src_to_dst_data[5] ;
 wire \src_to_dst_data[6] ;
 wire \src_to_dst_data[7] ;
 wire \src_to_dst_data[8] ;
 wire \src_to_dst_data[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;

 sky130_fd_sc_hd__clkbuf_2 _233_ (.A(src_data_valid_sync),
    .X(_141_));
 sky130_fd_sc_hd__xor2_4 _234_ (.A(src_req_prev),
    .B(src_req_sync),
    .X(_142_));
 sky130_fd_sc_hd__nand2_1 _235_ (.A(net170),
    .B(net69),
    .Y(_143_));
 sky130_fd_sc_hd__a32o_1 _236_ (.A1(_141_),
    .A2(\dst_state[0] ),
    .A3(_142_),
    .B1(_143_),
    .B2(\dst_state[2] ),
    .X(_003_));
 sky130_fd_sc_hd__buf_2 _237_ (.A(src_is_write_op_flag),
    .X(_144_));
 sky130_fd_sc_hd__xor2_2 _238_ (.A(dst_ack_prev),
    .B(dst_ack_sync),
    .X(_145_));
 sky130_fd_sc_hd__nor3b_2 _239_ (.A(net65),
    .B(net32),
    .C_N(\src_state[0] ),
    .Y(_146_));
 sky130_fd_sc_hd__a311o_1 _240_ (.A1(_144_),
    .A2(\src_state[1] ),
    .A3(_145_),
    .B1(_146_),
    .C1(\src_state[3] ),
    .X(_005_));
 sky130_fd_sc_hd__clkbuf_4 _241_ (.A(\src_state[2] ),
    .X(_147_));
 sky130_fd_sc_hd__buf_2 _242_ (.A(_147_),
    .X(_148_));
 sky130_fd_sc_hd__xnor2_4 _243_ (.A(dst_ack_prev),
    .B(dst_ack_sync),
    .Y(_149_));
 sky130_fd_sc_hd__nor2_1 _244_ (.A(_144_),
    .B(dst_data_valid_sync),
    .Y(_150_));
 sky130_fd_sc_hd__a21o_1 _245_ (.A1(_144_),
    .A2(_149_),
    .B1(_150_),
    .X(_151_));
 sky130_fd_sc_hd__a22o_1 _246_ (.A1(_148_),
    .A2(_145_),
    .B1(_151_),
    .B2(\src_state[1] ),
    .X(_006_));
 sky130_fd_sc_hd__nand2_1 _247_ (.A(_141_),
    .B(_142_),
    .Y(_152_));
 sky130_fd_sc_hd__nand3_1 _248_ (.A(net170),
    .B(net69),
    .C(dst_is_write_op),
    .Y(_153_));
 sky130_fd_sc_hd__o21ai_0 _249_ (.A1(_141_),
    .A2(dst_is_write_op),
    .B1(_153_),
    .Y(_154_));
 sky130_fd_sc_hd__a22o_1 _250_ (.A1(\dst_state[0] ),
    .A2(_152_),
    .B1(_154_),
    .B2(\dst_state[3] ),
    .X(_001_));
 sky130_fd_sc_hd__nor2b_1 _251_ (.A(dst_is_write_op),
    .B_N(net102),
    .Y(_155_));
 sky130_fd_sc_hd__a31oi_1 _252_ (.A1(_141_),
    .A2(dst_is_write_op),
    .A3(_142_),
    .B1(_155_),
    .Y(_156_));
 sky130_fd_sc_hd__a32o_1 _253_ (.A1(net170),
    .A2(net69),
    .A3(\dst_state[2] ),
    .B1(\dst_state[1] ),
    .B2(_156_),
    .X(_002_));
 sky130_fd_sc_hd__inv_1 _254_ (.A(\dst_state[3] ),
    .Y(_157_));
 sky130_fd_sc_hd__inv_1 _255_ (.A(\dst_state[1] ),
    .Y(_158_));
 sky130_fd_sc_hd__o22ai_1 _256_ (.A1(_157_),
    .A2(_154_),
    .B1(_156_),
    .B2(_158_),
    .Y(_004_));
 sky130_fd_sc_hd__o21ai_2 _257_ (.A1(net65),
    .A2(net32),
    .B1(\src_state[0] ),
    .Y(_159_));
 sky130_fd_sc_hd__buf_2 _258_ (.A(_159_),
    .X(_160_));
 sky130_fd_sc_hd__nand2_1 _259_ (.A(_148_),
    .B(_149_),
    .Y(_161_));
 sky130_fd_sc_hd__nand2_1 _260_ (.A(_160_),
    .B(_161_),
    .Y(_007_));
 sky130_fd_sc_hd__nand2_1 _261_ (.A(_157_),
    .B(_158_),
    .Y(net171));
 sky130_fd_sc_hd__nand2_2 _262_ (.A(\dst_state[1] ),
    .B(_155_),
    .Y(_162_));
 sky130_fd_sc_hd__clkbuf_4 _263_ (.A(_162_),
    .X(_163_));
 sky130_fd_sc_hd__o21ai_1 _264_ (.A1(_157_),
    .A2(dst_is_write_op),
    .B1(_163_),
    .Y(_231_));
 sky130_fd_sc_hd__a31o_1 _265_ (.A1(_141_),
    .A2(\dst_state[1] ),
    .A3(_142_),
    .B1(\dst_state[3] ),
    .X(_164_));
 sky130_fd_sc_hd__a21o_1 _266_ (.A1(dst_is_write_op),
    .A2(_164_),
    .B1(_003_),
    .X(_232_));
 sky130_fd_sc_hd__inv_1 _267_ (.A(_144_),
    .Y(_165_));
 sky130_fd_sc_hd__a21oi_1 _268_ (.A1(\src_state[1] ),
    .A2(_149_),
    .B1(_148_),
    .Y(_166_));
 sky130_fd_sc_hd__o211ai_1 _269_ (.A1(_165_),
    .A2(_166_),
    .B1(_161_),
    .C1(_160_),
    .Y(_230_));
 sky130_fd_sc_hd__nand3_4 _270_ (.A(_165_),
    .B(\src_state[1] ),
    .C(dst_data_valid_sync),
    .Y(_167_));
 sky130_fd_sc_hd__clkbuf_4 _271_ (.A(_167_),
    .X(_168_));
 sky130_fd_sc_hd__inv_1 _272_ (.A(_168_),
    .Y(_000_));
 sky130_fd_sc_hd__mux2_1 _273_ (.A0(\dst_state[0] ),
    .A1(dst_is_write_op),
    .S(\dst_state[1] ),
    .X(_169_));
 sky130_fd_sc_hd__nand3_4 _274_ (.A(_141_),
    .B(_142_),
    .C(_169_),
    .Y(_170_));
 sky130_fd_sc_hd__buf_6 _275_ (.A(_170_),
    .X(_171_));
 sky130_fd_sc_hd__xnor2_1 _276_ (.A(dst_ack),
    .B(_171_),
    .Y(_008_));
 sky130_fd_sc_hd__mux2_1 _277_ (.A0(\src_to_dst_data[0] ),
    .A1(net138),
    .S(_171_),
    .X(_009_));
 sky130_fd_sc_hd__mux2_1 _278_ (.A0(\src_to_dst_data[10] ),
    .A1(net139),
    .S(_171_),
    .X(_010_));
 sky130_fd_sc_hd__mux2_1 _279_ (.A0(\src_to_dst_data[11] ),
    .A1(net140),
    .S(_171_),
    .X(_011_));
 sky130_fd_sc_hd__mux2_1 _280_ (.A0(\src_to_dst_data[12] ),
    .A1(net141),
    .S(_171_),
    .X(_012_));
 sky130_fd_sc_hd__mux2_1 _281_ (.A0(\src_to_dst_data[13] ),
    .A1(net142),
    .S(_171_),
    .X(_013_));
 sky130_fd_sc_hd__mux2_1 _282_ (.A0(\src_to_dst_data[14] ),
    .A1(net143),
    .S(_171_),
    .X(_014_));
 sky130_fd_sc_hd__mux2_1 _283_ (.A0(\src_to_dst_data[15] ),
    .A1(net144),
    .S(_171_),
    .X(_015_));
 sky130_fd_sc_hd__mux2_1 _284_ (.A0(\src_to_dst_data[16] ),
    .A1(net145),
    .S(_171_),
    .X(_016_));
 sky130_fd_sc_hd__mux2_1 _285_ (.A0(\src_to_dst_data[17] ),
    .A1(net146),
    .S(_171_),
    .X(_017_));
 sky130_fd_sc_hd__buf_6 _286_ (.A(_170_),
    .X(_172_));
 sky130_fd_sc_hd__mux2_1 _287_ (.A0(\src_to_dst_data[18] ),
    .A1(net147),
    .S(_172_),
    .X(_018_));
 sky130_fd_sc_hd__mux2_1 _288_ (.A0(\src_to_dst_data[19] ),
    .A1(net148),
    .S(_172_),
    .X(_019_));
 sky130_fd_sc_hd__mux2_1 _289_ (.A0(\src_to_dst_data[1] ),
    .A1(net149),
    .S(_172_),
    .X(_020_));
 sky130_fd_sc_hd__mux2_1 _290_ (.A0(\src_to_dst_data[20] ),
    .A1(net150),
    .S(_172_),
    .X(_021_));
 sky130_fd_sc_hd__mux2_1 _291_ (.A0(\src_to_dst_data[21] ),
    .A1(net151),
    .S(_172_),
    .X(_022_));
 sky130_fd_sc_hd__mux2_1 _292_ (.A0(\src_to_dst_data[22] ),
    .A1(net152),
    .S(_172_),
    .X(_023_));
 sky130_fd_sc_hd__mux2_1 _293_ (.A0(\src_to_dst_data[23] ),
    .A1(net153),
    .S(_172_),
    .X(_024_));
 sky130_fd_sc_hd__mux2_1 _294_ (.A0(\src_to_dst_data[24] ),
    .A1(net154),
    .S(_172_),
    .X(_025_));
 sky130_fd_sc_hd__mux2_1 _295_ (.A0(\src_to_dst_data[25] ),
    .A1(net155),
    .S(_172_),
    .X(_026_));
 sky130_fd_sc_hd__mux2_1 _296_ (.A0(\src_to_dst_data[26] ),
    .A1(net156),
    .S(_172_),
    .X(_027_));
 sky130_fd_sc_hd__buf_6 _297_ (.A(_170_),
    .X(_173_));
 sky130_fd_sc_hd__mux2_1 _298_ (.A0(\src_to_dst_data[27] ),
    .A1(net157),
    .S(_173_),
    .X(_028_));
 sky130_fd_sc_hd__mux2_1 _299_ (.A0(\src_to_dst_data[28] ),
    .A1(net158),
    .S(_173_),
    .X(_029_));
 sky130_fd_sc_hd__mux2_1 _300_ (.A0(\src_to_dst_data[29] ),
    .A1(net159),
    .S(_173_),
    .X(_030_));
 sky130_fd_sc_hd__mux2_1 _301_ (.A0(\src_to_dst_data[2] ),
    .A1(net160),
    .S(_173_),
    .X(_031_));
 sky130_fd_sc_hd__mux2_1 _302_ (.A0(\src_to_dst_data[30] ),
    .A1(net161),
    .S(_173_),
    .X(_032_));
 sky130_fd_sc_hd__mux2_1 _303_ (.A0(\src_to_dst_data[31] ),
    .A1(net162),
    .S(_173_),
    .X(_033_));
 sky130_fd_sc_hd__mux2_1 _304_ (.A0(\src_to_dst_data[3] ),
    .A1(net163),
    .S(_173_),
    .X(_034_));
 sky130_fd_sc_hd__mux2_1 _305_ (.A0(\src_to_dst_data[4] ),
    .A1(net164),
    .S(_173_),
    .X(_035_));
 sky130_fd_sc_hd__mux2_1 _306_ (.A0(\src_to_dst_data[5] ),
    .A1(net165),
    .S(_173_),
    .X(_036_));
 sky130_fd_sc_hd__mux2_1 _307_ (.A0(\src_to_dst_data[6] ),
    .A1(net166),
    .S(_173_),
    .X(_037_));
 sky130_fd_sc_hd__mux2_1 _308_ (.A0(\src_to_dst_data[7] ),
    .A1(net167),
    .S(_170_),
    .X(_038_));
 sky130_fd_sc_hd__mux2_1 _309_ (.A0(\src_to_dst_data[8] ),
    .A1(net168),
    .S(_170_),
    .X(_039_));
 sky130_fd_sc_hd__mux2_1 _310_ (.A0(\src_to_dst_data[9] ),
    .A1(net169),
    .S(_170_),
    .X(_040_));
 sky130_fd_sc_hd__nand3_1 _311_ (.A(_141_),
    .B(\dst_state[0] ),
    .C(_142_),
    .Y(_174_));
 sky130_fd_sc_hd__mux2_1 _312_ (.A0(src_is_write_op_sync),
    .A1(dst_is_write_op),
    .S(_174_),
    .X(_041_));
 sky130_fd_sc_hd__mux2_1 _313_ (.A0(net70),
    .A1(\dst_to_src_data[0] ),
    .S(_163_),
    .X(_042_));
 sky130_fd_sc_hd__mux2_1 _314_ (.A0(net71),
    .A1(\dst_to_src_data[10] ),
    .S(_163_),
    .X(_043_));
 sky130_fd_sc_hd__mux2_1 _315_ (.A0(net72),
    .A1(\dst_to_src_data[11] ),
    .S(_163_),
    .X(_044_));
 sky130_fd_sc_hd__mux2_1 _316_ (.A0(net73),
    .A1(\dst_to_src_data[12] ),
    .S(_163_),
    .X(_045_));
 sky130_fd_sc_hd__mux2_1 _317_ (.A0(net74),
    .A1(\dst_to_src_data[13] ),
    .S(_163_),
    .X(_046_));
 sky130_fd_sc_hd__mux2_1 _318_ (.A0(net75),
    .A1(\dst_to_src_data[14] ),
    .S(_163_),
    .X(_047_));
 sky130_fd_sc_hd__mux2_1 _319_ (.A0(net76),
    .A1(\dst_to_src_data[15] ),
    .S(_163_),
    .X(_048_));
 sky130_fd_sc_hd__mux2_1 _320_ (.A0(net77),
    .A1(\dst_to_src_data[16] ),
    .S(_163_),
    .X(_049_));
 sky130_fd_sc_hd__mux2_1 _321_ (.A0(net78),
    .A1(\dst_to_src_data[17] ),
    .S(_163_),
    .X(_050_));
 sky130_fd_sc_hd__buf_4 _322_ (.A(_162_),
    .X(_175_));
 sky130_fd_sc_hd__mux2_1 _323_ (.A0(net79),
    .A1(\dst_to_src_data[18] ),
    .S(_175_),
    .X(_051_));
 sky130_fd_sc_hd__mux2_1 _324_ (.A0(net80),
    .A1(\dst_to_src_data[19] ),
    .S(_175_),
    .X(_052_));
 sky130_fd_sc_hd__mux2_1 _325_ (.A0(net81),
    .A1(\dst_to_src_data[1] ),
    .S(_175_),
    .X(_053_));
 sky130_fd_sc_hd__mux2_1 _326_ (.A0(net82),
    .A1(\dst_to_src_data[20] ),
    .S(_175_),
    .X(_054_));
 sky130_fd_sc_hd__mux2_1 _327_ (.A0(net83),
    .A1(\dst_to_src_data[21] ),
    .S(_175_),
    .X(_055_));
 sky130_fd_sc_hd__mux2_1 _328_ (.A0(net84),
    .A1(\dst_to_src_data[22] ),
    .S(_175_),
    .X(_056_));
 sky130_fd_sc_hd__mux2_1 _329_ (.A0(net85),
    .A1(\dst_to_src_data[23] ),
    .S(_175_),
    .X(_057_));
 sky130_fd_sc_hd__mux2_1 _330_ (.A0(net86),
    .A1(\dst_to_src_data[24] ),
    .S(_175_),
    .X(_058_));
 sky130_fd_sc_hd__mux2_1 _331_ (.A0(net87),
    .A1(\dst_to_src_data[25] ),
    .S(_175_),
    .X(_059_));
 sky130_fd_sc_hd__mux2_1 _332_ (.A0(net88),
    .A1(\dst_to_src_data[26] ),
    .S(_175_),
    .X(_060_));
 sky130_fd_sc_hd__buf_4 _333_ (.A(_162_),
    .X(_176_));
 sky130_fd_sc_hd__mux2_1 _334_ (.A0(net89),
    .A1(\dst_to_src_data[27] ),
    .S(_176_),
    .X(_061_));
 sky130_fd_sc_hd__mux2_1 _335_ (.A0(net90),
    .A1(\dst_to_src_data[28] ),
    .S(_176_),
    .X(_062_));
 sky130_fd_sc_hd__mux2_1 _336_ (.A0(net91),
    .A1(\dst_to_src_data[29] ),
    .S(_176_),
    .X(_063_));
 sky130_fd_sc_hd__mux2_1 _337_ (.A0(net92),
    .A1(\dst_to_src_data[2] ),
    .S(_176_),
    .X(_064_));
 sky130_fd_sc_hd__mux2_1 _338_ (.A0(net93),
    .A1(\dst_to_src_data[30] ),
    .S(_176_),
    .X(_065_));
 sky130_fd_sc_hd__mux2_1 _339_ (.A0(net94),
    .A1(\dst_to_src_data[31] ),
    .S(_176_),
    .X(_066_));
 sky130_fd_sc_hd__mux2_1 _340_ (.A0(net95),
    .A1(\dst_to_src_data[3] ),
    .S(_176_),
    .X(_067_));
 sky130_fd_sc_hd__mux2_1 _341_ (.A0(net96),
    .A1(\dst_to_src_data[4] ),
    .S(_176_),
    .X(_068_));
 sky130_fd_sc_hd__mux2_1 _342_ (.A0(net97),
    .A1(\dst_to_src_data[5] ),
    .S(_176_),
    .X(_069_));
 sky130_fd_sc_hd__mux2_1 _343_ (.A0(net98),
    .A1(\dst_to_src_data[6] ),
    .S(_176_),
    .X(_070_));
 sky130_fd_sc_hd__mux2_1 _344_ (.A0(net99),
    .A1(\dst_to_src_data[7] ),
    .S(_162_),
    .X(_071_));
 sky130_fd_sc_hd__mux2_1 _345_ (.A0(net100),
    .A1(\dst_to_src_data[8] ),
    .S(_162_),
    .X(_072_));
 sky130_fd_sc_hd__mux2_1 _346_ (.A0(net101),
    .A1(\dst_to_src_data[9] ),
    .S(_162_),
    .X(_073_));
 sky130_fd_sc_hd__mux2_1 _347_ (.A0(\dst_to_src_data[0] ),
    .A1(net105),
    .S(_168_),
    .X(_074_));
 sky130_fd_sc_hd__mux2_1 _348_ (.A0(\dst_to_src_data[10] ),
    .A1(net106),
    .S(_168_),
    .X(_075_));
 sky130_fd_sc_hd__mux2_1 _349_ (.A0(\dst_to_src_data[11] ),
    .A1(net107),
    .S(_168_),
    .X(_076_));
 sky130_fd_sc_hd__mux2_1 _350_ (.A0(\dst_to_src_data[12] ),
    .A1(net108),
    .S(_168_),
    .X(_077_));
 sky130_fd_sc_hd__mux2_1 _351_ (.A0(\dst_to_src_data[13] ),
    .A1(net109),
    .S(_168_),
    .X(_078_));
 sky130_fd_sc_hd__mux2_1 _352_ (.A0(\dst_to_src_data[14] ),
    .A1(net110),
    .S(_168_),
    .X(_079_));
 sky130_fd_sc_hd__mux2_1 _353_ (.A0(\dst_to_src_data[15] ),
    .A1(net111),
    .S(_168_),
    .X(_080_));
 sky130_fd_sc_hd__mux2_1 _354_ (.A0(\dst_to_src_data[16] ),
    .A1(net112),
    .S(_168_),
    .X(_081_));
 sky130_fd_sc_hd__mux2_1 _355_ (.A0(\dst_to_src_data[17] ),
    .A1(net113),
    .S(_168_),
    .X(_082_));
 sky130_fd_sc_hd__clkbuf_4 _356_ (.A(_167_),
    .X(_177_));
 sky130_fd_sc_hd__mux2_1 _357_ (.A0(\dst_to_src_data[18] ),
    .A1(net114),
    .S(_177_),
    .X(_083_));
 sky130_fd_sc_hd__mux2_1 _358_ (.A0(\dst_to_src_data[19] ),
    .A1(net115),
    .S(_177_),
    .X(_084_));
 sky130_fd_sc_hd__mux2_1 _359_ (.A0(\dst_to_src_data[1] ),
    .A1(net116),
    .S(_177_),
    .X(_085_));
 sky130_fd_sc_hd__mux2_1 _360_ (.A0(\dst_to_src_data[20] ),
    .A1(net117),
    .S(_177_),
    .X(_086_));
 sky130_fd_sc_hd__mux2_1 _361_ (.A0(\dst_to_src_data[21] ),
    .A1(net118),
    .S(_177_),
    .X(_087_));
 sky130_fd_sc_hd__mux2_1 _362_ (.A0(\dst_to_src_data[22] ),
    .A1(net119),
    .S(_177_),
    .X(_088_));
 sky130_fd_sc_hd__mux2_1 _363_ (.A0(\dst_to_src_data[23] ),
    .A1(net120),
    .S(_177_),
    .X(_089_));
 sky130_fd_sc_hd__mux2_1 _364_ (.A0(\dst_to_src_data[24] ),
    .A1(net121),
    .S(_177_),
    .X(_090_));
 sky130_fd_sc_hd__mux2_1 _365_ (.A0(\dst_to_src_data[25] ),
    .A1(net122),
    .S(_177_),
    .X(_091_));
 sky130_fd_sc_hd__mux2_1 _366_ (.A0(\dst_to_src_data[26] ),
    .A1(net123),
    .S(_177_),
    .X(_092_));
 sky130_fd_sc_hd__buf_4 _367_ (.A(_167_),
    .X(_178_));
 sky130_fd_sc_hd__mux2_1 _368_ (.A0(\dst_to_src_data[27] ),
    .A1(net124),
    .S(_178_),
    .X(_093_));
 sky130_fd_sc_hd__mux2_1 _369_ (.A0(\dst_to_src_data[28] ),
    .A1(net125),
    .S(_178_),
    .X(_094_));
 sky130_fd_sc_hd__mux2_1 _370_ (.A0(\dst_to_src_data[29] ),
    .A1(net126),
    .S(_178_),
    .X(_095_));
 sky130_fd_sc_hd__mux2_1 _371_ (.A0(\dst_to_src_data[2] ),
    .A1(net127),
    .S(_178_),
    .X(_096_));
 sky130_fd_sc_hd__mux2_1 _372_ (.A0(\dst_to_src_data[30] ),
    .A1(net128),
    .S(_178_),
    .X(_097_));
 sky130_fd_sc_hd__mux2_1 _373_ (.A0(\dst_to_src_data[31] ),
    .A1(net129),
    .S(_178_),
    .X(_098_));
 sky130_fd_sc_hd__mux2_1 _374_ (.A0(\dst_to_src_data[3] ),
    .A1(net130),
    .S(_178_),
    .X(_099_));
 sky130_fd_sc_hd__mux2_1 _375_ (.A0(\dst_to_src_data[4] ),
    .A1(net131),
    .S(_178_),
    .X(_100_));
 sky130_fd_sc_hd__mux2_1 _376_ (.A0(\dst_to_src_data[5] ),
    .A1(net132),
    .S(_178_),
    .X(_101_));
 sky130_fd_sc_hd__mux2_1 _377_ (.A0(\dst_to_src_data[6] ),
    .A1(net133),
    .S(_178_),
    .X(_102_));
 sky130_fd_sc_hd__mux2_1 _378_ (.A0(\dst_to_src_data[7] ),
    .A1(net134),
    .S(_167_),
    .X(_103_));
 sky130_fd_sc_hd__mux2_1 _379_ (.A0(\dst_to_src_data[8] ),
    .A1(net135),
    .S(_167_),
    .X(_104_));
 sky130_fd_sc_hd__mux2_1 _380_ (.A0(\dst_to_src_data[9] ),
    .A1(net136),
    .S(_167_),
    .X(_105_));
 sky130_fd_sc_hd__nor3b_1 _381_ (.A(\src_state[3] ),
    .B(\src_state[0] ),
    .C_N(net137),
    .Y(_179_));
 sky130_fd_sc_hd__or3b_1 _382_ (.A(\src_state[3] ),
    .B(\src_state[0] ),
    .C_N(\src_state[1] ),
    .X(_180_));
 sky130_fd_sc_hd__a211oi_1 _383_ (.A1(_144_),
    .A2(_149_),
    .B1(_150_),
    .C1(_180_),
    .Y(_181_));
 sky130_fd_sc_hd__a311o_1 _384_ (.A1(\src_state[1] ),
    .A2(net137),
    .A3(_151_),
    .B1(_179_),
    .C1(_181_),
    .X(_106_));
 sky130_fd_sc_hd__nand2_1 _385_ (.A(\src_state[0] ),
    .B(net32),
    .Y(_182_));
 sky130_fd_sc_hd__a22o_1 _386_ (.A1(\src_state[0] ),
    .A2(net65),
    .B1(_182_),
    .B2(_144_),
    .X(_107_));
 sky130_fd_sc_hd__mux2i_2 _387_ (.A0(\src_state[0] ),
    .A1(_144_),
    .S(\src_state[2] ),
    .Y(_183_));
 sky130_fd_sc_hd__a211oi_4 _388_ (.A1(\src_state[2] ),
    .A2(_149_),
    .B1(_146_),
    .C1(_183_),
    .Y(_184_));
 sky130_fd_sc_hd__buf_6 _389_ (.A(_184_),
    .X(_185_));
 sky130_fd_sc_hd__xor2_1 _390_ (.A(src_req),
    .B(_185_),
    .X(_108_));
 sky130_fd_sc_hd__nand4b_4 _391_ (.A_N(_146_),
    .B(_147_),
    .C(_144_),
    .D(_145_),
    .Y(_186_));
 sky130_fd_sc_hd__clkbuf_4 _392_ (.A(_186_),
    .X(_187_));
 sky130_fd_sc_hd__or3_1 _393_ (.A(_148_),
    .B(net11),
    .C(_160_),
    .X(_188_));
 sky130_fd_sc_hd__o221a_1 _394_ (.A1(\src_to_dst_data[0] ),
    .A2(_185_),
    .B1(_187_),
    .B2(net33),
    .C1(_188_),
    .X(_109_));
 sky130_fd_sc_hd__or3_1 _395_ (.A(_148_),
    .B(net12),
    .C(_160_),
    .X(_189_));
 sky130_fd_sc_hd__o221a_1 _396_ (.A1(\src_to_dst_data[10] ),
    .A2(_185_),
    .B1(_187_),
    .B2(net34),
    .C1(_189_),
    .X(_110_));
 sky130_fd_sc_hd__or3_1 _397_ (.A(_148_),
    .B(net13),
    .C(_160_),
    .X(_190_));
 sky130_fd_sc_hd__o221a_1 _398_ (.A1(\src_to_dst_data[11] ),
    .A2(_185_),
    .B1(_187_),
    .B2(net35),
    .C1(_190_),
    .X(_111_));
 sky130_fd_sc_hd__or3_1 _399_ (.A(_148_),
    .B(net14),
    .C(_160_),
    .X(_191_));
 sky130_fd_sc_hd__o221a_1 _400_ (.A1(\src_to_dst_data[12] ),
    .A2(_185_),
    .B1(_187_),
    .B2(net36),
    .C1(_191_),
    .X(_112_));
 sky130_fd_sc_hd__or3_1 _401_ (.A(_148_),
    .B(net15),
    .C(_160_),
    .X(_192_));
 sky130_fd_sc_hd__o221a_1 _402_ (.A1(\src_to_dst_data[13] ),
    .A2(_185_),
    .B1(_187_),
    .B2(net37),
    .C1(_192_),
    .X(_113_));
 sky130_fd_sc_hd__buf_2 _403_ (.A(_147_),
    .X(_193_));
 sky130_fd_sc_hd__or3_1 _404_ (.A(_193_),
    .B(net16),
    .C(_160_),
    .X(_194_));
 sky130_fd_sc_hd__o221a_1 _405_ (.A1(\src_to_dst_data[14] ),
    .A2(_185_),
    .B1(_187_),
    .B2(net38),
    .C1(_194_),
    .X(_114_));
 sky130_fd_sc_hd__or3_1 _406_ (.A(_193_),
    .B(net17),
    .C(_160_),
    .X(_195_));
 sky130_fd_sc_hd__o221a_1 _407_ (.A1(\src_to_dst_data[15] ),
    .A2(_185_),
    .B1(_187_),
    .B2(net39),
    .C1(_195_),
    .X(_115_));
 sky130_fd_sc_hd__or3_1 _408_ (.A(_193_),
    .B(net18),
    .C(_160_),
    .X(_196_));
 sky130_fd_sc_hd__o221a_1 _409_ (.A1(\src_to_dst_data[16] ),
    .A2(_185_),
    .B1(_187_),
    .B2(net40),
    .C1(_196_),
    .X(_116_));
 sky130_fd_sc_hd__clkbuf_2 _410_ (.A(_159_),
    .X(_197_));
 sky130_fd_sc_hd__or3_1 _411_ (.A(_193_),
    .B(net19),
    .C(_197_),
    .X(_198_));
 sky130_fd_sc_hd__o221a_1 _412_ (.A1(\src_to_dst_data[17] ),
    .A2(_185_),
    .B1(_187_),
    .B2(net41),
    .C1(_198_),
    .X(_117_));
 sky130_fd_sc_hd__buf_6 _413_ (.A(_184_),
    .X(_199_));
 sky130_fd_sc_hd__or3_1 _414_ (.A(_193_),
    .B(net20),
    .C(_197_),
    .X(_200_));
 sky130_fd_sc_hd__o221a_1 _415_ (.A1(\src_to_dst_data[18] ),
    .A2(_199_),
    .B1(_187_),
    .B2(net42),
    .C1(_200_),
    .X(_118_));
 sky130_fd_sc_hd__clkbuf_4 _416_ (.A(_186_),
    .X(_201_));
 sky130_fd_sc_hd__or3_1 _417_ (.A(_193_),
    .B(net21),
    .C(_197_),
    .X(_202_));
 sky130_fd_sc_hd__o221a_1 _418_ (.A1(\src_to_dst_data[19] ),
    .A2(_199_),
    .B1(_201_),
    .B2(net43),
    .C1(_202_),
    .X(_119_));
 sky130_fd_sc_hd__or3_1 _419_ (.A(_193_),
    .B(net22),
    .C(_197_),
    .X(_203_));
 sky130_fd_sc_hd__o221a_1 _420_ (.A1(\src_to_dst_data[1] ),
    .A2(_199_),
    .B1(_201_),
    .B2(net44),
    .C1(_203_),
    .X(_120_));
 sky130_fd_sc_hd__nor2_1 _421_ (.A(net65),
    .B(net23),
    .Y(_204_));
 sky130_fd_sc_hd__nand2_1 _422_ (.A(_148_),
    .B(net45),
    .Y(_205_));
 sky130_fd_sc_hd__o21ai_1 _423_ (.A1(_148_),
    .A2(_204_),
    .B1(_205_),
    .Y(_206_));
 sky130_fd_sc_hd__mux2_1 _424_ (.A0(\src_to_dst_data[20] ),
    .A1(_206_),
    .S(_184_),
    .X(_121_));
 sky130_fd_sc_hd__or3_1 _425_ (.A(_193_),
    .B(net66),
    .C(_197_),
    .X(_207_));
 sky130_fd_sc_hd__o221a_1 _426_ (.A1(\src_to_dst_data[21] ),
    .A2(_199_),
    .B1(_201_),
    .B2(net46),
    .C1(_207_),
    .X(_122_));
 sky130_fd_sc_hd__or3_1 _427_ (.A(_193_),
    .B(net67),
    .C(_197_),
    .X(_208_));
 sky130_fd_sc_hd__o221a_1 _428_ (.A1(\src_to_dst_data[22] ),
    .A2(_199_),
    .B1(_201_),
    .B2(net47),
    .C1(_208_),
    .X(_123_));
 sky130_fd_sc_hd__or3_1 _429_ (.A(_193_),
    .B(net68),
    .C(_197_),
    .X(_209_));
 sky130_fd_sc_hd__o221a_1 _430_ (.A1(\src_to_dst_data[23] ),
    .A2(_199_),
    .B1(_201_),
    .B2(net48),
    .C1(_209_),
    .X(_124_));
 sky130_fd_sc_hd__buf_2 _431_ (.A(_147_),
    .X(_210_));
 sky130_fd_sc_hd__or3_1 _432_ (.A(_210_),
    .B(net1),
    .C(_197_),
    .X(_211_));
 sky130_fd_sc_hd__o221a_1 _433_ (.A1(\src_to_dst_data[24] ),
    .A2(_199_),
    .B1(_201_),
    .B2(net49),
    .C1(_211_),
    .X(_125_));
 sky130_fd_sc_hd__or3_1 _434_ (.A(_210_),
    .B(net2),
    .C(_197_),
    .X(_212_));
 sky130_fd_sc_hd__o221a_1 _435_ (.A1(\src_to_dst_data[25] ),
    .A2(_199_),
    .B1(_201_),
    .B2(net50),
    .C1(_212_),
    .X(_126_));
 sky130_fd_sc_hd__or3_1 _436_ (.A(_210_),
    .B(net3),
    .C(_197_),
    .X(_213_));
 sky130_fd_sc_hd__o221a_1 _437_ (.A1(\src_to_dst_data[26] ),
    .A2(_199_),
    .B1(_201_),
    .B2(net51),
    .C1(_213_),
    .X(_127_));
 sky130_fd_sc_hd__clkbuf_2 _438_ (.A(_159_),
    .X(_214_));
 sky130_fd_sc_hd__or3_1 _439_ (.A(_210_),
    .B(net4),
    .C(_214_),
    .X(_215_));
 sky130_fd_sc_hd__o221a_1 _440_ (.A1(\src_to_dst_data[27] ),
    .A2(_199_),
    .B1(_201_),
    .B2(net52),
    .C1(_215_),
    .X(_128_));
 sky130_fd_sc_hd__buf_6 _441_ (.A(_184_),
    .X(_216_));
 sky130_fd_sc_hd__or3_1 _442_ (.A(_210_),
    .B(net5),
    .C(_214_),
    .X(_217_));
 sky130_fd_sc_hd__o221a_1 _443_ (.A1(\src_to_dst_data[28] ),
    .A2(_216_),
    .B1(_201_),
    .B2(net53),
    .C1(_217_),
    .X(_129_));
 sky130_fd_sc_hd__buf_2 _444_ (.A(_186_),
    .X(_218_));
 sky130_fd_sc_hd__or3_1 _445_ (.A(_210_),
    .B(net6),
    .C(_214_),
    .X(_219_));
 sky130_fd_sc_hd__o221a_1 _446_ (.A1(\src_to_dst_data[29] ),
    .A2(_216_),
    .B1(_218_),
    .B2(net54),
    .C1(_219_),
    .X(_130_));
 sky130_fd_sc_hd__or3_1 _447_ (.A(_210_),
    .B(net24),
    .C(_214_),
    .X(_220_));
 sky130_fd_sc_hd__o221a_1 _448_ (.A1(\src_to_dst_data[2] ),
    .A2(_216_),
    .B1(_218_),
    .B2(net55),
    .C1(_220_),
    .X(_131_));
 sky130_fd_sc_hd__or3_1 _449_ (.A(_210_),
    .B(net7),
    .C(_214_),
    .X(_221_));
 sky130_fd_sc_hd__o221a_1 _450_ (.A1(\src_to_dst_data[30] ),
    .A2(_216_),
    .B1(_218_),
    .B2(net56),
    .C1(_221_),
    .X(_132_));
 sky130_fd_sc_hd__or3_1 _451_ (.A(_210_),
    .B(net8),
    .C(_214_),
    .X(_222_));
 sky130_fd_sc_hd__o221a_1 _452_ (.A1(\src_to_dst_data[31] ),
    .A2(_216_),
    .B1(_218_),
    .B2(net57),
    .C1(_222_),
    .X(_133_));
 sky130_fd_sc_hd__or3_1 _453_ (.A(_210_),
    .B(net25),
    .C(_214_),
    .X(_223_));
 sky130_fd_sc_hd__o221a_1 _454_ (.A1(\src_to_dst_data[3] ),
    .A2(_216_),
    .B1(_218_),
    .B2(net58),
    .C1(_223_),
    .X(_134_));
 sky130_fd_sc_hd__or3_1 _455_ (.A(_147_),
    .B(net26),
    .C(_214_),
    .X(_224_));
 sky130_fd_sc_hd__o221a_1 _456_ (.A1(\src_to_dst_data[4] ),
    .A2(_216_),
    .B1(_218_),
    .B2(net59),
    .C1(_224_),
    .X(_135_));
 sky130_fd_sc_hd__or3_1 _457_ (.A(_147_),
    .B(net27),
    .C(_214_),
    .X(_225_));
 sky130_fd_sc_hd__o221a_1 _458_ (.A1(\src_to_dst_data[5] ),
    .A2(_216_),
    .B1(_218_),
    .B2(net60),
    .C1(_225_),
    .X(_136_));
 sky130_fd_sc_hd__or3_1 _459_ (.A(_147_),
    .B(net28),
    .C(_214_),
    .X(_226_));
 sky130_fd_sc_hd__o221a_1 _460_ (.A1(\src_to_dst_data[6] ),
    .A2(_216_),
    .B1(_218_),
    .B2(net61),
    .C1(_226_),
    .X(_137_));
 sky130_fd_sc_hd__or3_1 _461_ (.A(_147_),
    .B(net29),
    .C(_159_),
    .X(_227_));
 sky130_fd_sc_hd__o221a_1 _462_ (.A1(\src_to_dst_data[7] ),
    .A2(_216_),
    .B1(_218_),
    .B2(net62),
    .C1(_227_),
    .X(_138_));
 sky130_fd_sc_hd__or3_1 _463_ (.A(_147_),
    .B(net30),
    .C(_159_),
    .X(_228_));
 sky130_fd_sc_hd__o221a_1 _464_ (.A1(\src_to_dst_data[8] ),
    .A2(_184_),
    .B1(_218_),
    .B2(net63),
    .C1(_228_),
    .X(_139_));
 sky130_fd_sc_hd__or3_1 _465_ (.A(_147_),
    .B(net31),
    .C(_159_),
    .X(_229_));
 sky130_fd_sc_hd__o221a_1 _466_ (.A1(\src_to_dst_data[9] ),
    .A2(_184_),
    .B1(_186_),
    .B2(net64),
    .C1(_229_),
    .X(_140_));
 sky130_fd_sc_hd__dfrtp_1 \dst_ack$_DFFE_PN0P_  (.D(_008_),
    .Q(dst_ack),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_2 \dst_ack_prev$_DFF_PN0_  (.D(dst_ack_sync),
    .Q(dst_ack_prev),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \dst_ack_sync_reg[0]$_DFF_PN0_  (.D(dst_ack),
    .Q(\dst_ack_sync_reg[0] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_2 \dst_ack_sync_reg[1]$_DFF_PN0_  (.D(\dst_ack_sync_reg[0] ),
    .Q(dst_ack_sync),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[0]$_DFFE_PN0P_  (.D(_009_),
    .Q(net138),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[10]$_DFFE_PN0P_  (.D(_010_),
    .Q(net139),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[11]$_DFFE_PN0P_  (.D(_011_),
    .Q(net140),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[12]$_DFFE_PN0P_  (.D(_012_),
    .Q(net141),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[13]$_DFFE_PN0P_  (.D(_013_),
    .Q(net142),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[14]$_DFFE_PN0P_  (.D(_014_),
    .Q(net143),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[15]$_DFFE_PN0P_  (.D(_015_),
    .Q(net144),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[16]$_DFFE_PN0P_  (.D(_016_),
    .Q(net145),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[17]$_DFFE_PN0P_  (.D(_017_),
    .Q(net146),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[18]$_DFFE_PN0P_  (.D(_018_),
    .Q(net147),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[19]$_DFFE_PN0P_  (.D(_019_),
    .Q(net148),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[1]$_DFFE_PN0P_  (.D(_020_),
    .Q(net149),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[20]$_DFFE_PN0P_  (.D(_021_),
    .Q(net150),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[21]$_DFFE_PN0P_  (.D(_022_),
    .Q(net151),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[22]$_DFFE_PN0P_  (.D(_023_),
    .Q(net152),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[23]$_DFFE_PN0P_  (.D(_024_),
    .Q(net153),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[24]$_DFFE_PN0P_  (.D(_025_),
    .Q(net154),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[25]$_DFFE_PN0P_  (.D(_026_),
    .Q(net155),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[26]$_DFFE_PN0P_  (.D(_027_),
    .Q(net156),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[27]$_DFFE_PN0P_  (.D(_028_),
    .Q(net157),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[28]$_DFFE_PN0P_  (.D(_029_),
    .Q(net158),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[29]$_DFFE_PN0P_  (.D(_030_),
    .Q(net159),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[2]$_DFFE_PN0P_  (.D(_031_),
    .Q(net160),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[30]$_DFFE_PN0P_  (.D(_032_),
    .Q(net161),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[31]$_DFFE_PN0P_  (.D(_033_),
    .Q(net162),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[3]$_DFFE_PN0P_  (.D(_034_),
    .Q(net163),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[4]$_DFFE_PN0P_  (.D(_035_),
    .Q(net164),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[5]$_DFFE_PN0P_  (.D(_036_),
    .Q(net165),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[6]$_DFFE_PN0P_  (.D(_037_),
    .Q(net166),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[7]$_DFFE_PN0P_  (.D(_038_),
    .Q(net167),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[8]$_DFFE_PN0P_  (.D(_039_),
    .Q(net168),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_reg[9]$_DFFE_PN0P_  (.D(_040_),
    .Q(net169),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_valid$_DFF_PN0_  (.D(_231_),
    .Q(dst_data_valid),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_valid_sync_reg[0]$_DFF_PN0_  (.D(dst_data_valid),
    .Q(\dst_data_valid_sync_reg[0] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \dst_data_valid_sync_reg[1]$_DFF_PN0_  (.D(\dst_data_valid_sync_reg[0] ),
    .Q(dst_data_valid_sync),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_2 \dst_is_write_op$_DFFE_PN0P_  (.D(_041_),
    .Q(dst_is_write_op),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfstp_1 \dst_state[0]$_DFF_PN1_  (.D(_001_),
    .Q(\dst_state[0] ),
    .SET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_state[1]$_DFF_PN0_  (.D(_002_),
    .Q(\dst_state[1] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_state[2]$_DFF_PN0_  (.D(_003_),
    .Q(\dst_state[2] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_state[3]$_DFF_PN0_  (.D(_004_),
    .Q(\dst_state[3] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[0]$_DFFE_PN0P_  (.D(_042_),
    .Q(\dst_to_src_data[0] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[10]$_DFFE_PN0P_  (.D(_043_),
    .Q(\dst_to_src_data[10] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[11]$_DFFE_PN0P_  (.D(_044_),
    .Q(\dst_to_src_data[11] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[12]$_DFFE_PN0P_  (.D(_045_),
    .Q(\dst_to_src_data[12] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[13]$_DFFE_PN0P_  (.D(_046_),
    .Q(\dst_to_src_data[13] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[14]$_DFFE_PN0P_  (.D(_047_),
    .Q(\dst_to_src_data[14] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[15]$_DFFE_PN0P_  (.D(_048_),
    .Q(\dst_to_src_data[15] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[16]$_DFFE_PN0P_  (.D(_049_),
    .Q(\dst_to_src_data[16] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[17]$_DFFE_PN0P_  (.D(_050_),
    .Q(\dst_to_src_data[17] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[18]$_DFFE_PN0P_  (.D(_051_),
    .Q(\dst_to_src_data[18] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[19]$_DFFE_PN0P_  (.D(_052_),
    .Q(\dst_to_src_data[19] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[1]$_DFFE_PN0P_  (.D(_053_),
    .Q(\dst_to_src_data[1] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[20]$_DFFE_PN0P_  (.D(_054_),
    .Q(\dst_to_src_data[20] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[21]$_DFFE_PN0P_  (.D(_055_),
    .Q(\dst_to_src_data[21] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[22]$_DFFE_PN0P_  (.D(_056_),
    .Q(\dst_to_src_data[22] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[23]$_DFFE_PN0P_  (.D(_057_),
    .Q(\dst_to_src_data[23] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[24]$_DFFE_PN0P_  (.D(_058_),
    .Q(\dst_to_src_data[24] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[25]$_DFFE_PN0P_  (.D(_059_),
    .Q(\dst_to_src_data[25] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[26]$_DFFE_PN0P_  (.D(_060_),
    .Q(\dst_to_src_data[26] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[27]$_DFFE_PN0P_  (.D(_061_),
    .Q(\dst_to_src_data[27] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[28]$_DFFE_PN0P_  (.D(_062_),
    .Q(\dst_to_src_data[28] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[29]$_DFFE_PN0P_  (.D(_063_),
    .Q(\dst_to_src_data[29] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[2]$_DFFE_PN0P_  (.D(_064_),
    .Q(\dst_to_src_data[2] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[30]$_DFFE_PN0P_  (.D(_065_),
    .Q(\dst_to_src_data[30] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[31]$_DFFE_PN0P_  (.D(_066_),
    .Q(\dst_to_src_data[31] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[3]$_DFFE_PN0P_  (.D(_067_),
    .Q(\dst_to_src_data[3] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[4]$_DFFE_PN0P_  (.D(_068_),
    .Q(\dst_to_src_data[4] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[5]$_DFFE_PN0P_  (.D(_069_),
    .Q(\dst_to_src_data[5] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[6]$_DFFE_PN0P_  (.D(_070_),
    .Q(\dst_to_src_data[6] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[7]$_DFFE_PN0P_  (.D(_071_),
    .Q(\dst_to_src_data[7] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[8]$_DFFE_PN0P_  (.D(_072_),
    .Q(\dst_to_src_data[8] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_to_src_data[9]$_DFFE_PN0P_  (.D(_073_),
    .Q(\dst_to_src_data[9] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \dst_valid$_DFF_PN0_  (.D(_232_),
    .Q(net170),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[0]$_DFFE_PN0P_  (.D(_074_),
    .Q(net105),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[10]$_DFFE_PN0P_  (.D(_075_),
    .Q(net106),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[11]$_DFFE_PN0P_  (.D(_076_),
    .Q(net107),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[12]$_DFFE_PN0P_  (.D(_077_),
    .Q(net108),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[13]$_DFFE_PN0P_  (.D(_078_),
    .Q(net109),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[14]$_DFFE_PN0P_  (.D(_079_),
    .Q(net110),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[15]$_DFFE_PN0P_  (.D(_080_),
    .Q(net111),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[16]$_DFFE_PN0P_  (.D(_081_),
    .Q(net112),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[17]$_DFFE_PN0P_  (.D(_082_),
    .Q(net113),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[18]$_DFFE_PN0P_  (.D(_083_),
    .Q(net114),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[19]$_DFFE_PN0P_  (.D(_084_),
    .Q(net115),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[1]$_DFFE_PN0P_  (.D(_085_),
    .Q(net116),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[20]$_DFFE_PN0P_  (.D(_086_),
    .Q(net117),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[21]$_DFFE_PN0P_  (.D(_087_),
    .Q(net118),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[22]$_DFFE_PN0P_  (.D(_088_),
    .Q(net119),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[23]$_DFFE_PN0P_  (.D(_089_),
    .Q(net120),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[24]$_DFFE_PN0P_  (.D(_090_),
    .Q(net121),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[25]$_DFFE_PN0P_  (.D(_091_),
    .Q(net122),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[26]$_DFFE_PN0P_  (.D(_092_),
    .Q(net123),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[27]$_DFFE_PN0P_  (.D(_093_),
    .Q(net124),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[28]$_DFFE_PN0P_  (.D(_094_),
    .Q(net125),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[29]$_DFFE_PN0P_  (.D(_095_),
    .Q(net126),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[2]$_DFFE_PN0P_  (.D(_096_),
    .Q(net127),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[30]$_DFFE_PN0P_  (.D(_097_),
    .Q(net128),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[31]$_DFFE_PN0P_  (.D(_098_),
    .Q(net129),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[3]$_DFFE_PN0P_  (.D(_099_),
    .Q(net130),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[4]$_DFFE_PN0P_  (.D(_100_),
    .Q(net131),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[5]$_DFFE_PN0P_  (.D(_101_),
    .Q(net132),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[6]$_DFFE_PN0P_  (.D(_102_),
    .Q(net133),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[7]$_DFFE_PN0P_  (.D(_103_),
    .Q(net134),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[8]$_DFFE_PN0P_  (.D(_104_),
    .Q(net135),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[9]$_DFFE_PN0P_  (.D(_105_),
    .Q(net136),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \mem_ready$_DFFE_PN0P_  (.D(_106_),
    .Q(net137),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_data_valid$_DFF_PN0_  (.D(_230_),
    .Q(src_data_valid),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_data_valid_sync_reg[0]$_DFF_PN0_  (.D(src_data_valid),
    .Q(\src_data_valid_sync_reg[0] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \src_data_valid_sync_reg[1]$_DFF_PN0_  (.D(\src_data_valid_sync_reg[0] ),
    .Q(src_data_valid_sync),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \src_is_write_op$_DFFE_PN0P_  (.D(_107_),
    .Q(src_is_write_op_flag),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_is_write_op_sync_reg[0]$_DFF_PN0_  (.D(src_is_write_op_flag),
    .Q(\src_is_write_op_sync_reg[0] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \src_is_write_op_sync_reg[1]$_DFF_PN0_  (.D(\src_is_write_op_sync_reg[0] ),
    .Q(src_is_write_op_sync),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \src_req$_DFFE_PN0P_  (.D(_108_),
    .Q(src_req),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_req_prev$_DFF_PN0_  (.D(src_req_sync),
    .Q(src_req_prev),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \src_req_sync_reg[0]$_DFF_PN0_  (.D(src_req),
    .Q(\src_req_sync_reg[0] ),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfrtp_1 \src_req_sync_reg[1]$_DFF_PN0_  (.D(\src_req_sync_reg[0] ),
    .Q(src_req_sync),
    .RESET_B(net10),
    .CLK(net9));
 sky130_fd_sc_hd__dfstp_1 \src_state[0]$_DFF_PN1_  (.D(_005_),
    .Q(\src_state[0] ),
    .SET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_2 \src_state[1]$_DFF_PN0_  (.D(_006_),
    .Q(\src_state[1] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_2 \src_state[2]$_DFF_PN0_  (.D(_007_),
    .Q(\src_state[2] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_state[3]$_DFF_PN0_  (.D(_000_),
    .Q(\src_state[3] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[0]$_DFFE_PN0P_  (.D(_109_),
    .Q(\src_to_dst_data[0] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[10]$_DFFE_PN0P_  (.D(_110_),
    .Q(\src_to_dst_data[10] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[11]$_DFFE_PN0P_  (.D(_111_),
    .Q(\src_to_dst_data[11] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[12]$_DFFE_PN0P_  (.D(_112_),
    .Q(\src_to_dst_data[12] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[13]$_DFFE_PN0P_  (.D(_113_),
    .Q(\src_to_dst_data[13] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[14]$_DFFE_PN0P_  (.D(_114_),
    .Q(\src_to_dst_data[14] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[15]$_DFFE_PN0P_  (.D(_115_),
    .Q(\src_to_dst_data[15] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[16]$_DFFE_PN0P_  (.D(_116_),
    .Q(\src_to_dst_data[16] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[17]$_DFFE_PN0P_  (.D(_117_),
    .Q(\src_to_dst_data[17] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[18]$_DFFE_PN0P_  (.D(_118_),
    .Q(\src_to_dst_data[18] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[19]$_DFFE_PN0P_  (.D(_119_),
    .Q(\src_to_dst_data[19] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[1]$_DFFE_PN0P_  (.D(_120_),
    .Q(\src_to_dst_data[1] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[20]$_DFFE_PN0P_  (.D(_121_),
    .Q(\src_to_dst_data[20] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[21]$_DFFE_PN0P_  (.D(_122_),
    .Q(\src_to_dst_data[21] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[22]$_DFFE_PN0P_  (.D(_123_),
    .Q(\src_to_dst_data[22] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[23]$_DFFE_PN0P_  (.D(_124_),
    .Q(\src_to_dst_data[23] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[24]$_DFFE_PN0P_  (.D(_125_),
    .Q(\src_to_dst_data[24] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[25]$_DFFE_PN0P_  (.D(_126_),
    .Q(\src_to_dst_data[25] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[26]$_DFFE_PN0P_  (.D(_127_),
    .Q(\src_to_dst_data[26] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[27]$_DFFE_PN0P_  (.D(_128_),
    .Q(\src_to_dst_data[27] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[28]$_DFFE_PN0P_  (.D(_129_),
    .Q(\src_to_dst_data[28] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[29]$_DFFE_PN0P_  (.D(_130_),
    .Q(\src_to_dst_data[29] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[2]$_DFFE_PN0P_  (.D(_131_),
    .Q(\src_to_dst_data[2] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[30]$_DFFE_PN0P_  (.D(_132_),
    .Q(\src_to_dst_data[30] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[31]$_DFFE_PN0P_  (.D(_133_),
    .Q(\src_to_dst_data[31] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[3]$_DFFE_PN0P_  (.D(_134_),
    .Q(\src_to_dst_data[3] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[4]$_DFFE_PN0P_  (.D(_135_),
    .Q(\src_to_dst_data[4] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[5]$_DFFE_PN0P_  (.D(_136_),
    .Q(\src_to_dst_data[5] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[6]$_DFFE_PN0P_  (.D(_137_),
    .Q(\src_to_dst_data[6] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[7]$_DFFE_PN0P_  (.D(_138_),
    .Q(\src_to_dst_data[7] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[8]$_DFFE_PN0P_  (.D(_139_),
    .Q(\src_to_dst_data[8] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__dfrtp_1 \src_to_dst_data[9]$_DFFE_PN0P_  (.D(_140_),
    .Q(\src_to_dst_data[9] ),
    .RESET_B(net104),
    .CLK(net103));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_135 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(dest_id[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(dest_id[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(dest_id[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(dest_id[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(dest_id[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(dest_id[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(dest_id[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(dest_id[7]),
    .X(net8));
 sky130_fd_sc_hd__buf_16 input9 (.A(dst_clk),
    .X(net9));
 sky130_fd_sc_hd__buf_16 input10 (.A(dst_rst_n),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(mem_addr[0]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(mem_addr[10]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(mem_addr[11]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(mem_addr[12]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(mem_addr[13]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(mem_addr[14]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(mem_addr[15]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(mem_addr[16]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(mem_addr[17]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(mem_addr[18]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(mem_addr[19]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(mem_addr[1]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(mem_addr[20]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(mem_addr[2]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(mem_addr[3]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(mem_addr[4]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(mem_addr[5]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(mem_addr[6]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(mem_addr[7]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(mem_addr[8]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(mem_addr[9]),
    .X(net31));
 sky130_fd_sc_hd__dlymetal6s2s_1 input32 (.A(mem_read),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(mem_wdata[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(mem_wdata[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(mem_wdata[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(mem_wdata[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(mem_wdata[13]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(mem_wdata[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(mem_wdata[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(mem_wdata[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(mem_wdata[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(mem_wdata[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(mem_wdata[19]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(mem_wdata[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(mem_wdata[20]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(mem_wdata[21]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(mem_wdata[22]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(mem_wdata[23]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(mem_wdata[24]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(mem_wdata[25]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(mem_wdata[26]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(mem_wdata[27]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(mem_wdata[28]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(mem_wdata[29]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(mem_wdata[2]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(mem_wdata[30]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(mem_wdata[31]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(mem_wdata[3]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(mem_wdata[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(mem_wdata[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(mem_wdata[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(mem_wdata[7]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(mem_wdata[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(mem_wdata[9]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 input65 (.A(mem_write),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(msg_type[0]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(msg_type[1]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(msg_type[2]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(router_in_ready),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(router_out_data[0]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(router_out_data[10]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(router_out_data[11]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(router_out_data[12]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 input74 (.A(router_out_data[13]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 input75 (.A(router_out_data[14]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(router_out_data[15]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(router_out_data[16]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(router_out_data[17]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input79 (.A(router_out_data[18]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 input80 (.A(router_out_data[19]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 input81 (.A(router_out_data[1]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input82 (.A(router_out_data[20]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 input83 (.A(router_out_data[21]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(router_out_data[22]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(router_out_data[23]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(router_out_data[24]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(router_out_data[25]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(router_out_data[26]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 input89 (.A(router_out_data[27]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 input90 (.A(router_out_data[28]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(router_out_data[29]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 input92 (.A(router_out_data[2]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 input93 (.A(router_out_data[30]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 input94 (.A(router_out_data[31]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 input95 (.A(router_out_data[3]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 input96 (.A(router_out_data[4]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 input97 (.A(router_out_data[5]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 input98 (.A(router_out_data[6]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 input99 (.A(router_out_data[7]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 input100 (.A(router_out_data[8]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 input101 (.A(router_out_data[9]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 input102 (.A(router_out_valid),
    .X(net102));
 sky130_fd_sc_hd__buf_16 input103 (.A(src_clk),
    .X(net103));
 sky130_fd_sc_hd__buf_16 input104 (.A(src_rst_n),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 output105 (.A(net105),
    .X(mem_rdata[0]));
 sky130_fd_sc_hd__clkbuf_1 output106 (.A(net106),
    .X(mem_rdata[10]));
 sky130_fd_sc_hd__clkbuf_1 output107 (.A(net107),
    .X(mem_rdata[11]));
 sky130_fd_sc_hd__clkbuf_1 output108 (.A(net108),
    .X(mem_rdata[12]));
 sky130_fd_sc_hd__clkbuf_1 output109 (.A(net109),
    .X(mem_rdata[13]));
 sky130_fd_sc_hd__clkbuf_1 output110 (.A(net110),
    .X(mem_rdata[14]));
 sky130_fd_sc_hd__clkbuf_1 output111 (.A(net111),
    .X(mem_rdata[15]));
 sky130_fd_sc_hd__clkbuf_1 output112 (.A(net112),
    .X(mem_rdata[16]));
 sky130_fd_sc_hd__clkbuf_1 output113 (.A(net113),
    .X(mem_rdata[17]));
 sky130_fd_sc_hd__clkbuf_1 output114 (.A(net114),
    .X(mem_rdata[18]));
 sky130_fd_sc_hd__clkbuf_1 output115 (.A(net115),
    .X(mem_rdata[19]));
 sky130_fd_sc_hd__clkbuf_1 output116 (.A(net116),
    .X(mem_rdata[1]));
 sky130_fd_sc_hd__clkbuf_1 output117 (.A(net117),
    .X(mem_rdata[20]));
 sky130_fd_sc_hd__clkbuf_1 output118 (.A(net118),
    .X(mem_rdata[21]));
 sky130_fd_sc_hd__clkbuf_1 output119 (.A(net119),
    .X(mem_rdata[22]));
 sky130_fd_sc_hd__clkbuf_1 output120 (.A(net120),
    .X(mem_rdata[23]));
 sky130_fd_sc_hd__clkbuf_1 output121 (.A(net121),
    .X(mem_rdata[24]));
 sky130_fd_sc_hd__clkbuf_1 output122 (.A(net122),
    .X(mem_rdata[25]));
 sky130_fd_sc_hd__clkbuf_1 output123 (.A(net123),
    .X(mem_rdata[26]));
 sky130_fd_sc_hd__clkbuf_1 output124 (.A(net124),
    .X(mem_rdata[27]));
 sky130_fd_sc_hd__clkbuf_1 output125 (.A(net125),
    .X(mem_rdata[28]));
 sky130_fd_sc_hd__clkbuf_1 output126 (.A(net126),
    .X(mem_rdata[29]));
 sky130_fd_sc_hd__clkbuf_1 output127 (.A(net127),
    .X(mem_rdata[2]));
 sky130_fd_sc_hd__clkbuf_1 output128 (.A(net128),
    .X(mem_rdata[30]));
 sky130_fd_sc_hd__clkbuf_1 output129 (.A(net129),
    .X(mem_rdata[31]));
 sky130_fd_sc_hd__clkbuf_1 output130 (.A(net130),
    .X(mem_rdata[3]));
 sky130_fd_sc_hd__clkbuf_1 output131 (.A(net131),
    .X(mem_rdata[4]));
 sky130_fd_sc_hd__clkbuf_1 output132 (.A(net132),
    .X(mem_rdata[5]));
 sky130_fd_sc_hd__clkbuf_1 output133 (.A(net133),
    .X(mem_rdata[6]));
 sky130_fd_sc_hd__clkbuf_1 output134 (.A(net134),
    .X(mem_rdata[7]));
 sky130_fd_sc_hd__clkbuf_1 output135 (.A(net135),
    .X(mem_rdata[8]));
 sky130_fd_sc_hd__clkbuf_1 output136 (.A(net136),
    .X(mem_rdata[9]));
 sky130_fd_sc_hd__clkbuf_1 output137 (.A(net137),
    .X(mem_ready));
 sky130_fd_sc_hd__clkbuf_1 output138 (.A(net138),
    .X(router_in_data[0]));
 sky130_fd_sc_hd__clkbuf_1 output139 (.A(net139),
    .X(router_in_data[10]));
 sky130_fd_sc_hd__clkbuf_1 output140 (.A(net140),
    .X(router_in_data[11]));
 sky130_fd_sc_hd__clkbuf_1 output141 (.A(net141),
    .X(router_in_data[12]));
 sky130_fd_sc_hd__clkbuf_1 output142 (.A(net142),
    .X(router_in_data[13]));
 sky130_fd_sc_hd__clkbuf_1 output143 (.A(net143),
    .X(router_in_data[14]));
 sky130_fd_sc_hd__clkbuf_1 output144 (.A(net144),
    .X(router_in_data[15]));
 sky130_fd_sc_hd__clkbuf_1 output145 (.A(net145),
    .X(router_in_data[16]));
 sky130_fd_sc_hd__clkbuf_1 output146 (.A(net146),
    .X(router_in_data[17]));
 sky130_fd_sc_hd__clkbuf_1 output147 (.A(net147),
    .X(router_in_data[18]));
 sky130_fd_sc_hd__clkbuf_1 output148 (.A(net148),
    .X(router_in_data[19]));
 sky130_fd_sc_hd__clkbuf_1 output149 (.A(net149),
    .X(router_in_data[1]));
 sky130_fd_sc_hd__clkbuf_1 output150 (.A(net150),
    .X(router_in_data[20]));
 sky130_fd_sc_hd__clkbuf_1 output151 (.A(net151),
    .X(router_in_data[21]));
 sky130_fd_sc_hd__clkbuf_1 output152 (.A(net152),
    .X(router_in_data[22]));
 sky130_fd_sc_hd__clkbuf_1 output153 (.A(net153),
    .X(router_in_data[23]));
 sky130_fd_sc_hd__clkbuf_1 output154 (.A(net154),
    .X(router_in_data[24]));
 sky130_fd_sc_hd__clkbuf_1 output155 (.A(net155),
    .X(router_in_data[25]));
 sky130_fd_sc_hd__clkbuf_1 output156 (.A(net156),
    .X(router_in_data[26]));
 sky130_fd_sc_hd__clkbuf_1 output157 (.A(net157),
    .X(router_in_data[27]));
 sky130_fd_sc_hd__clkbuf_1 output158 (.A(net158),
    .X(router_in_data[28]));
 sky130_fd_sc_hd__clkbuf_1 output159 (.A(net159),
    .X(router_in_data[29]));
 sky130_fd_sc_hd__clkbuf_1 output160 (.A(net160),
    .X(router_in_data[2]));
 sky130_fd_sc_hd__clkbuf_1 output161 (.A(net161),
    .X(router_in_data[30]));
 sky130_fd_sc_hd__clkbuf_1 output162 (.A(net162),
    .X(router_in_data[31]));
 sky130_fd_sc_hd__clkbuf_1 output163 (.A(net163),
    .X(router_in_data[3]));
 sky130_fd_sc_hd__clkbuf_1 output164 (.A(net164),
    .X(router_in_data[4]));
 sky130_fd_sc_hd__clkbuf_1 output165 (.A(net165),
    .X(router_in_data[5]));
 sky130_fd_sc_hd__clkbuf_1 output166 (.A(net166),
    .X(router_in_data[6]));
 sky130_fd_sc_hd__clkbuf_1 output167 (.A(net167),
    .X(router_in_data[7]));
 sky130_fd_sc_hd__clkbuf_1 output168 (.A(net168),
    .X(router_in_data[8]));
 sky130_fd_sc_hd__clkbuf_1 output169 (.A(net169),
    .X(router_in_data[9]));
 sky130_fd_sc_hd__clkbuf_1 output170 (.A(net170),
    .X(router_in_valid));
 sky130_fd_sc_hd__clkbuf_1 output171 (.A(net171),
    .X(router_out_ready));
 sky130_fd_sc_hd__fill_4 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_84 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_186 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_113 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_21 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_194 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_54 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_25 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_186 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_19 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_90 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_126 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_57 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_92 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_186 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_220 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_225 ();
endmodule
