module parameterized_fft (busy,
    clk,
    data_ready,
    data_valid_in,
    data_valid_out,
    rst_n,
    start,
    data_in_imag,
    data_in_real,
    data_out_imag,
    data_out_real);
 output busy;
 input clk;
 output data_ready;
 input data_valid_in;
 output data_valid_out;
 input rst_n;
 input start;
 input [15:0] data_in_imag;
 input [15:0] data_in_real;
 output [127:0] data_out_imag;
 output [127:0] data_out_real;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire net56;
 wire net60;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire net22;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire net6;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire net8;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire net10;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire net7;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire net9;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire net3;
 wire _01602_;
 wire _01603_;
 wire net4;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire net33;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire net414;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire net13;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire net12;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire net16;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire net30;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire net11;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire net5;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire net52;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire net129;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire net132;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire net125;
 wire _05421_;
 wire net137;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire net156;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire net149;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire net154;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire net153;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire net152;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire net158;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire net151;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire net133;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire net58;
 wire _05836_;
 wire net57;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire net98;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire net94;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire net59;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire net97;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire clknet_leaf_0_clk;
 wire net398;
 wire \bit_rev_idx[0] ;
 wire \bit_rev_idx[1] ;
 wire \bit_rev_idx[2] ;
 wire \butterfly_count[0] ;
 wire \butterfly_count[1] ;
 wire \butterfly_count[2] ;
 wire \butterfly_in_group[0] ;
 wire \butterfly_in_group[1] ;
 wire \butterfly_in_group[2] ;
 wire \group[0] ;
 wire \group[1] ;
 wire \group[2] ;
 wire \idx1[0] ;
 wire \idx1[1] ;
 wire \idx1[2] ;
 wire \idx2[0] ;
 wire \idx2[1] ;
 wire \idx2[2] ;
 wire \sample_count[0] ;
 wire \sample_count[1] ;
 wire \sample_count[2] ;
 wire \samples_imag[0][0] ;
 wire \samples_imag[0][10] ;
 wire \samples_imag[0][11] ;
 wire \samples_imag[0][12] ;
 wire \samples_imag[0][13] ;
 wire \samples_imag[0][14] ;
 wire \samples_imag[0][15] ;
 wire \samples_imag[0][1] ;
 wire \samples_imag[0][2] ;
 wire \samples_imag[0][3] ;
 wire \samples_imag[0][4] ;
 wire \samples_imag[0][5] ;
 wire \samples_imag[0][6] ;
 wire \samples_imag[0][7] ;
 wire \samples_imag[0][8] ;
 wire \samples_imag[0][9] ;
 wire \samples_imag[1][0] ;
 wire \samples_imag[1][10] ;
 wire \samples_imag[1][11] ;
 wire \samples_imag[1][12] ;
 wire \samples_imag[1][13] ;
 wire \samples_imag[1][14] ;
 wire \samples_imag[1][15] ;
 wire \samples_imag[1][1] ;
 wire \samples_imag[1][2] ;
 wire \samples_imag[1][3] ;
 wire \samples_imag[1][4] ;
 wire \samples_imag[1][5] ;
 wire \samples_imag[1][6] ;
 wire \samples_imag[1][7] ;
 wire \samples_imag[1][8] ;
 wire \samples_imag[1][9] ;
 wire \samples_imag[2][0] ;
 wire \samples_imag[2][10] ;
 wire \samples_imag[2][11] ;
 wire \samples_imag[2][12] ;
 wire \samples_imag[2][13] ;
 wire \samples_imag[2][14] ;
 wire \samples_imag[2][15] ;
 wire \samples_imag[2][1] ;
 wire \samples_imag[2][2] ;
 wire \samples_imag[2][3] ;
 wire \samples_imag[2][4] ;
 wire \samples_imag[2][5] ;
 wire \samples_imag[2][6] ;
 wire \samples_imag[2][7] ;
 wire \samples_imag[2][8] ;
 wire \samples_imag[2][9] ;
 wire \samples_imag[3][0] ;
 wire \samples_imag[3][10] ;
 wire \samples_imag[3][11] ;
 wire \samples_imag[3][12] ;
 wire \samples_imag[3][13] ;
 wire \samples_imag[3][14] ;
 wire \samples_imag[3][15] ;
 wire \samples_imag[3][1] ;
 wire \samples_imag[3][2] ;
 wire \samples_imag[3][3] ;
 wire \samples_imag[3][4] ;
 wire \samples_imag[3][5] ;
 wire \samples_imag[3][6] ;
 wire \samples_imag[3][7] ;
 wire \samples_imag[3][8] ;
 wire \samples_imag[3][9] ;
 wire \samples_imag[4][0] ;
 wire \samples_imag[4][10] ;
 wire \samples_imag[4][11] ;
 wire \samples_imag[4][12] ;
 wire \samples_imag[4][13] ;
 wire \samples_imag[4][14] ;
 wire \samples_imag[4][15] ;
 wire \samples_imag[4][1] ;
 wire \samples_imag[4][2] ;
 wire \samples_imag[4][3] ;
 wire \samples_imag[4][4] ;
 wire \samples_imag[4][5] ;
 wire \samples_imag[4][6] ;
 wire \samples_imag[4][7] ;
 wire \samples_imag[4][8] ;
 wire \samples_imag[4][9] ;
 wire \samples_imag[5][0] ;
 wire \samples_imag[5][10] ;
 wire \samples_imag[5][11] ;
 wire \samples_imag[5][12] ;
 wire \samples_imag[5][13] ;
 wire \samples_imag[5][14] ;
 wire \samples_imag[5][15] ;
 wire \samples_imag[5][1] ;
 wire \samples_imag[5][2] ;
 wire \samples_imag[5][3] ;
 wire \samples_imag[5][4] ;
 wire \samples_imag[5][5] ;
 wire \samples_imag[5][6] ;
 wire \samples_imag[5][7] ;
 wire \samples_imag[5][8] ;
 wire \samples_imag[5][9] ;
 wire \samples_imag[6][0] ;
 wire \samples_imag[6][10] ;
 wire \samples_imag[6][11] ;
 wire \samples_imag[6][12] ;
 wire \samples_imag[6][13] ;
 wire \samples_imag[6][14] ;
 wire \samples_imag[6][15] ;
 wire \samples_imag[6][1] ;
 wire \samples_imag[6][2] ;
 wire \samples_imag[6][3] ;
 wire \samples_imag[6][4] ;
 wire \samples_imag[6][5] ;
 wire \samples_imag[6][6] ;
 wire \samples_imag[6][7] ;
 wire \samples_imag[6][8] ;
 wire \samples_imag[6][9] ;
 wire \samples_imag[7][0] ;
 wire \samples_imag[7][10] ;
 wire \samples_imag[7][11] ;
 wire \samples_imag[7][12] ;
 wire \samples_imag[7][13] ;
 wire \samples_imag[7][14] ;
 wire \samples_imag[7][15] ;
 wire \samples_imag[7][1] ;
 wire \samples_imag[7][2] ;
 wire \samples_imag[7][3] ;
 wire \samples_imag[7][4] ;
 wire \samples_imag[7][5] ;
 wire \samples_imag[7][6] ;
 wire \samples_imag[7][7] ;
 wire \samples_imag[7][8] ;
 wire \samples_imag[7][9] ;
 wire \samples_real[0][0] ;
 wire \samples_real[0][10] ;
 wire \samples_real[0][11] ;
 wire \samples_real[0][12] ;
 wire \samples_real[0][13] ;
 wire \samples_real[0][14] ;
 wire \samples_real[0][15] ;
 wire \samples_real[0][1] ;
 wire \samples_real[0][2] ;
 wire \samples_real[0][3] ;
 wire \samples_real[0][4] ;
 wire \samples_real[0][5] ;
 wire \samples_real[0][6] ;
 wire \samples_real[0][7] ;
 wire \samples_real[0][8] ;
 wire \samples_real[0][9] ;
 wire \samples_real[1][0] ;
 wire \samples_real[1][10] ;
 wire \samples_real[1][11] ;
 wire \samples_real[1][12] ;
 wire \samples_real[1][13] ;
 wire \samples_real[1][14] ;
 wire \samples_real[1][15] ;
 wire \samples_real[1][1] ;
 wire \samples_real[1][2] ;
 wire \samples_real[1][3] ;
 wire \samples_real[1][4] ;
 wire \samples_real[1][5] ;
 wire \samples_real[1][6] ;
 wire \samples_real[1][7] ;
 wire \samples_real[1][8] ;
 wire \samples_real[1][9] ;
 wire \samples_real[2][0] ;
 wire \samples_real[2][10] ;
 wire \samples_real[2][11] ;
 wire \samples_real[2][12] ;
 wire \samples_real[2][13] ;
 wire \samples_real[2][14] ;
 wire \samples_real[2][15] ;
 wire \samples_real[2][1] ;
 wire \samples_real[2][2] ;
 wire \samples_real[2][3] ;
 wire \samples_real[2][4] ;
 wire \samples_real[2][5] ;
 wire \samples_real[2][6] ;
 wire \samples_real[2][7] ;
 wire \samples_real[2][8] ;
 wire \samples_real[2][9] ;
 wire \samples_real[3][0] ;
 wire \samples_real[3][10] ;
 wire \samples_real[3][11] ;
 wire \samples_real[3][12] ;
 wire \samples_real[3][13] ;
 wire \samples_real[3][14] ;
 wire \samples_real[3][15] ;
 wire \samples_real[3][1] ;
 wire \samples_real[3][2] ;
 wire \samples_real[3][3] ;
 wire \samples_real[3][4] ;
 wire \samples_real[3][5] ;
 wire \samples_real[3][6] ;
 wire \samples_real[3][7] ;
 wire \samples_real[3][8] ;
 wire \samples_real[3][9] ;
 wire \samples_real[4][0] ;
 wire \samples_real[4][10] ;
 wire \samples_real[4][11] ;
 wire \samples_real[4][12] ;
 wire \samples_real[4][13] ;
 wire \samples_real[4][14] ;
 wire \samples_real[4][15] ;
 wire \samples_real[4][1] ;
 wire \samples_real[4][2] ;
 wire \samples_real[4][3] ;
 wire \samples_real[4][4] ;
 wire \samples_real[4][5] ;
 wire \samples_real[4][6] ;
 wire \samples_real[4][7] ;
 wire \samples_real[4][8] ;
 wire \samples_real[4][9] ;
 wire \samples_real[5][0] ;
 wire \samples_real[5][10] ;
 wire \samples_real[5][11] ;
 wire \samples_real[5][12] ;
 wire \samples_real[5][13] ;
 wire \samples_real[5][14] ;
 wire \samples_real[5][15] ;
 wire \samples_real[5][1] ;
 wire \samples_real[5][2] ;
 wire \samples_real[5][3] ;
 wire \samples_real[5][4] ;
 wire \samples_real[5][5] ;
 wire \samples_real[5][6] ;
 wire \samples_real[5][7] ;
 wire \samples_real[5][8] ;
 wire \samples_real[5][9] ;
 wire \samples_real[6][0] ;
 wire \samples_real[6][10] ;
 wire \samples_real[6][11] ;
 wire \samples_real[6][12] ;
 wire \samples_real[6][13] ;
 wire \samples_real[6][14] ;
 wire \samples_real[6][15] ;
 wire \samples_real[6][1] ;
 wire \samples_real[6][2] ;
 wire \samples_real[6][3] ;
 wire \samples_real[6][4] ;
 wire \samples_real[6][5] ;
 wire \samples_real[6][6] ;
 wire \samples_real[6][7] ;
 wire \samples_real[6][8] ;
 wire \samples_real[6][9] ;
 wire \samples_real[7][0] ;
 wire \samples_real[7][10] ;
 wire \samples_real[7][11] ;
 wire \samples_real[7][12] ;
 wire \samples_real[7][13] ;
 wire \samples_real[7][14] ;
 wire \samples_real[7][15] ;
 wire \samples_real[7][1] ;
 wire \samples_real[7][2] ;
 wire \samples_real[7][3] ;
 wire \samples_real[7][4] ;
 wire \samples_real[7][5] ;
 wire \samples_real[7][6] ;
 wire \samples_real[7][7] ;
 wire \samples_real[7][8] ;
 wire \samples_real[7][9] ;
 wire \stage[0] ;
 wire \stage[1] ;
 wire \stage[2] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire \temp_imag[0] ;
 wire \temp_real[0] ;
 wire \twiddle_idx[0] ;
 wire \twiddle_idx[1] ;
 wire net1;
 wire net2;
 wire net14;
 wire net15;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net31;
 wire net32;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net51;
 wire net53;
 wire net61;
 wire net93;
 wire net101;
 wire net104;
 wire net107;
 wire net130;
 wire net131;
 wire net138;
 wire net139;
 wire net140;
 wire net143;
 wire net144;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net54;
 wire net55;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net95;
 wire net96;
 wire net99;
 wire net100;
 wire net102;
 wire net103;
 wire net105;
 wire net106;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net126;
 wire net127;
 wire net128;
 wire net134;
 wire net135;
 wire net136;
 wire net141;
 wire net142;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net150;
 wire net155;
 wire net157;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net429;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net481;
 wire net482;
 wire net483;
 wire net491;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net512;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net520;
 wire net426;
 wire net428;
 wire net437;
 wire net438;
 wire net443;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net470;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net511;
 wire net513;
 wire net521;
 wire net522;
 wire net524;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net534;

 BUF_X2 _09753_ (.A(rst_n),
    .Z(_00841_));
 BUF_X4 _09754_ (.A(_00841_),
    .Z(_00842_));
 INV_X4 _09755_ (.A(_00842_),
    .ZN(_00843_));
 BUF_X4 _09756_ (.A(_00843_),
    .Z(_00844_));
 BUF_X4 _09757_ (.A(_00844_),
    .Z(_00845_));
 BUF_X2 _09758_ (.A(\state[1] ),
    .Z(_00846_));
 CLKBUF_X3 _09759_ (.A(\stage[2] ),
    .Z(_00847_));
 BUF_X4 _09760_ (.A(_00847_),
    .Z(_00848_));
 BUF_X2 _09761_ (.A(\stage[0] ),
    .Z(_00849_));
 BUF_X2 _09762_ (.A(\stage[1] ),
    .Z(_00850_));
 AOI21_X4 _09763_ (.A(_00848_),
    .B1(_00849_),
    .B2(_00850_),
    .ZN(_00851_));
 NAND2_X1 _09764_ (.A1(_00846_),
    .A2(_00851_),
    .ZN(_00852_));
 CLKBUF_X3 _09765_ (.A(\state[2] ),
    .Z(_00853_));
 NAND3_X1 _09766_ (.A1(net86),
    .A2(_09382_),
    .A3(_00853_),
    .ZN(_00854_));
 AOI21_X1 _09767_ (.A(_00845_),
    .B1(_00852_),
    .B2(_00854_),
    .ZN(_00011_));
 CLKBUF_X3 _09768_ (.A(_00842_),
    .Z(_00855_));
 BUF_X4 _09769_ (.A(_00855_),
    .Z(_00856_));
 BUF_X4 _09770_ (.A(\state[3] ),
    .Z(_00857_));
 INV_X4 _09771_ (.A(_00857_),
    .ZN(_00858_));
 CLKBUF_X3 _09772_ (.A(_00858_),
    .Z(_00859_));
 BUF_X2 _09773_ (.A(\state[0] ),
    .Z(_00860_));
 INV_X1 _09774_ (.A(net87),
    .ZN(_00861_));
 NAND2_X1 _09775_ (.A1(_00860_),
    .A2(_00861_),
    .ZN(_00862_));
 NAND3_X1 _09776_ (.A1(_00856_),
    .A2(_00859_),
    .A3(_00862_),
    .ZN(_00010_));
 CLKBUF_X2 split56 (.A(net61),
    .Z(net56));
 BUF_X4 clone60 (.A(net452),
    .Z(net60));
 MUX2_X1 _09779_ (.A(\samples_imag[0][15] ),
    .B(\samples_imag[2][15] ),
    .S(net56),
    .Z(_00865_));
 MUX2_X1 _09780_ (.A(\samples_imag[1][15] ),
    .B(\samples_imag[3][15] ),
    .S(net56),
    .Z(_00866_));
 BUF_X4 _09781_ (.A(_00000_),
    .Z(_00867_));
 MUX2_X1 _09782_ (.A(_00865_),
    .B(_00866_),
    .S(_00867_),
    .Z(_00868_));
 MUX2_X1 _09783_ (.A(\samples_imag[4][15] ),
    .B(\samples_imag[6][15] ),
    .S(net56),
    .Z(_00869_));
 MUX2_X1 _09784_ (.A(\samples_imag[5][15] ),
    .B(\samples_imag[7][15] ),
    .S(net56),
    .Z(_00870_));
 MUX2_X1 _09785_ (.A(_00869_),
    .B(_00870_),
    .S(_00867_),
    .Z(_00871_));
 BUF_X2 _09786_ (.A(_00002_),
    .Z(_00872_));
 MUX2_X2 _09787_ (.A(_00868_),
    .B(_00871_),
    .S(_00872_),
    .Z(_08561_));
 BUF_X16 _09788_ (.A(_00001_),
    .Z(_00873_));
 BUF_X4 _09789_ (.A(net57),
    .Z(_00874_));
 MUX2_X1 _09790_ (.A(\samples_imag[0][14] ),
    .B(\samples_imag[2][14] ),
    .S(_00874_),
    .Z(_00875_));
 MUX2_X1 _09791_ (.A(\samples_imag[1][14] ),
    .B(\samples_imag[3][14] ),
    .S(_00874_),
    .Z(_00876_));
 BUF_X4 _09792_ (.A(_00867_),
    .Z(_00877_));
 MUX2_X1 _09793_ (.A(_00875_),
    .B(_00876_),
    .S(_00877_),
    .Z(_00878_));
 MUX2_X1 _09794_ (.A(\samples_imag[4][14] ),
    .B(\samples_imag[6][14] ),
    .S(_00874_),
    .Z(_00879_));
 MUX2_X1 _09795_ (.A(\samples_imag[5][14] ),
    .B(\samples_imag[7][14] ),
    .S(_00874_),
    .Z(_00880_));
 MUX2_X1 _09796_ (.A(_00879_),
    .B(_00880_),
    .S(_00877_),
    .Z(_00881_));
 BUF_X4 _09797_ (.A(_00872_),
    .Z(_00882_));
 MUX2_X2 _09798_ (.A(_00878_),
    .B(_00881_),
    .S(_00882_),
    .Z(_08553_));
 BUF_X16 _09799_ (.A(_00873_),
    .Z(_00883_));
 MUX2_X1 _09800_ (.A(\samples_imag[0][13] ),
    .B(\samples_imag[2][13] ),
    .S(_00883_),
    .Z(_00884_));
 MUX2_X1 _09801_ (.A(\samples_imag[1][13] ),
    .B(\samples_imag[3][13] ),
    .S(_00883_),
    .Z(_00885_));
 BUF_X4 _09802_ (.A(_00867_),
    .Z(_00886_));
 MUX2_X1 _09803_ (.A(_00884_),
    .B(_00885_),
    .S(_00886_),
    .Z(_00887_));
 MUX2_X1 _09804_ (.A(\samples_imag[4][13] ),
    .B(\samples_imag[6][13] ),
    .S(_00883_),
    .Z(_00888_));
 MUX2_X1 _09805_ (.A(\samples_imag[5][13] ),
    .B(\samples_imag[7][13] ),
    .S(_00883_),
    .Z(_00889_));
 MUX2_X1 _09806_ (.A(_00888_),
    .B(_00889_),
    .S(_00886_),
    .Z(_00890_));
 MUX2_X2 _09807_ (.A(_00887_),
    .B(_00890_),
    .S(_00882_),
    .Z(_08569_));
 BUF_X4 _09808_ (.A(net57),
    .Z(_00891_));
 MUX2_X1 _09809_ (.A(\samples_imag[0][12] ),
    .B(\samples_imag[2][12] ),
    .S(_00891_),
    .Z(_00892_));
 MUX2_X1 _09810_ (.A(\samples_imag[1][12] ),
    .B(\samples_imag[3][12] ),
    .S(_00891_),
    .Z(_00893_));
 BUF_X4 _09811_ (.A(_00867_),
    .Z(_00894_));
 MUX2_X1 _09812_ (.A(_00892_),
    .B(_00893_),
    .S(_00894_),
    .Z(_00895_));
 BUF_X4 _09813_ (.A(net57),
    .Z(_00896_));
 MUX2_X1 _09814_ (.A(\samples_imag[4][12] ),
    .B(\samples_imag[6][12] ),
    .S(_00896_),
    .Z(_00897_));
 MUX2_X1 _09815_ (.A(\samples_imag[5][12] ),
    .B(\samples_imag[7][12] ),
    .S(_00896_),
    .Z(_00898_));
 BUF_X4 _09816_ (.A(_00867_),
    .Z(_00899_));
 MUX2_X1 _09817_ (.A(_00897_),
    .B(_00898_),
    .S(_00899_),
    .Z(_00900_));
 BUF_X4 _09818_ (.A(_00872_),
    .Z(_00901_));
 MUX2_X2 _09819_ (.A(_00895_),
    .B(_00900_),
    .S(_00901_),
    .Z(_08574_));
 BUF_X4 _09820_ (.A(_00873_),
    .Z(_00902_));
 MUX2_X1 _09821_ (.A(\samples_imag[0][11] ),
    .B(\samples_imag[2][11] ),
    .S(net59),
    .Z(_00903_));
 MUX2_X1 _09822_ (.A(\samples_imag[1][11] ),
    .B(\samples_imag[3][11] ),
    .S(net59),
    .Z(_00904_));
 MUX2_X1 _09823_ (.A(_00903_),
    .B(_00904_),
    .S(_00886_),
    .Z(_00905_));
 BUF_X4 _09824_ (.A(net57),
    .Z(_00906_));
 MUX2_X1 _09825_ (.A(\samples_imag[4][11] ),
    .B(\samples_imag[6][11] ),
    .S(_00906_),
    .Z(_00907_));
 MUX2_X1 _09826_ (.A(\samples_imag[5][11] ),
    .B(\samples_imag[7][11] ),
    .S(_00906_),
    .Z(_00908_));
 MUX2_X1 _09827_ (.A(_00907_),
    .B(_00908_),
    .S(_00877_),
    .Z(_00909_));
 MUX2_X2 _09828_ (.A(_00905_),
    .B(_00909_),
    .S(_00882_),
    .Z(_08579_));
 BUF_X8 _09829_ (.A(_00873_),
    .Z(_00910_));
 MUX2_X1 _09830_ (.A(\samples_imag[0][10] ),
    .B(\samples_imag[2][10] ),
    .S(net129),
    .Z(_00911_));
 MUX2_X1 _09831_ (.A(\samples_imag[1][10] ),
    .B(\samples_imag[3][10] ),
    .S(_00910_),
    .Z(_00912_));
 BUF_X4 _09832_ (.A(_00867_),
    .Z(_00913_));
 MUX2_X1 _09833_ (.A(_00911_),
    .B(_00912_),
    .S(_00913_),
    .Z(_00914_));
 MUX2_X1 _09834_ (.A(\samples_imag[4][10] ),
    .B(\samples_imag[6][10] ),
    .S(_00910_),
    .Z(_00915_));
 MUX2_X1 _09835_ (.A(\samples_imag[5][10] ),
    .B(\samples_imag[7][10] ),
    .S(_00910_),
    .Z(_00916_));
 MUX2_X1 _09836_ (.A(_00915_),
    .B(_00916_),
    .S(_00913_),
    .Z(_00917_));
 BUF_X4 _09837_ (.A(_00872_),
    .Z(_00918_));
 MUX2_X2 _09838_ (.A(_00914_),
    .B(_00917_),
    .S(_00918_),
    .Z(_08584_));
 BUF_X8 _09839_ (.A(_00001_),
    .Z(_00919_));
 MUX2_X1 _09840_ (.A(\samples_imag[0][9] ),
    .B(\samples_imag[2][9] ),
    .S(net60),
    .Z(_00920_));
 BUF_X4 _09841_ (.A(_00001_),
    .Z(_00921_));
 MUX2_X1 _09842_ (.A(\samples_imag[1][9] ),
    .B(\samples_imag[3][9] ),
    .S(_00921_),
    .Z(_00922_));
 BUF_X4 _09843_ (.A(_00867_),
    .Z(_00923_));
 MUX2_X1 _09844_ (.A(_00920_),
    .B(_00922_),
    .S(_00923_),
    .Z(_00924_));
 MUX2_X1 _09845_ (.A(\samples_imag[4][9] ),
    .B(\samples_imag[6][9] ),
    .S(_00921_),
    .Z(_00925_));
 MUX2_X1 _09846_ (.A(\samples_imag[5][9] ),
    .B(\samples_imag[7][9] ),
    .S(_00921_),
    .Z(_00926_));
 MUX2_X1 _09847_ (.A(_00925_),
    .B(_00926_),
    .S(_00923_),
    .Z(_00927_));
 MUX2_X2 _09848_ (.A(_00924_),
    .B(_00927_),
    .S(_00918_),
    .Z(_08589_));
 MUX2_X1 _09849_ (.A(\samples_imag[0][8] ),
    .B(\samples_imag[2][8] ),
    .S(_00921_),
    .Z(_00928_));
 MUX2_X1 _09850_ (.A(\samples_imag[1][8] ),
    .B(\samples_imag[3][8] ),
    .S(_00921_),
    .Z(_00929_));
 MUX2_X1 _09851_ (.A(_00928_),
    .B(_00929_),
    .S(_00923_),
    .Z(_00930_));
 BUF_X16 _09852_ (.A(_00873_),
    .Z(_00931_));
 MUX2_X1 _09853_ (.A(\samples_imag[4][8] ),
    .B(\samples_imag[6][8] ),
    .S(net476),
    .Z(_00932_));
 MUX2_X1 _09854_ (.A(\samples_imag[5][8] ),
    .B(\samples_imag[7][8] ),
    .S(net476),
    .Z(_00933_));
 MUX2_X1 _09855_ (.A(_00932_),
    .B(_00933_),
    .S(_00913_),
    .Z(_00934_));
 MUX2_X2 _09856_ (.A(_00930_),
    .B(_00934_),
    .S(_00918_),
    .Z(_08594_));
 BUF_X4 _09857_ (.A(net57),
    .Z(_00935_));
 MUX2_X1 _09858_ (.A(\samples_imag[0][7] ),
    .B(\samples_imag[2][7] ),
    .S(_00935_),
    .Z(_00936_));
 MUX2_X1 _09859_ (.A(\samples_imag[1][7] ),
    .B(\samples_imag[3][7] ),
    .S(_00935_),
    .Z(_00937_));
 MUX2_X1 _09860_ (.A(_00936_),
    .B(_00937_),
    .S(_00899_),
    .Z(_00938_));
 MUX2_X1 _09861_ (.A(\samples_imag[4][7] ),
    .B(\samples_imag[6][7] ),
    .S(_00935_),
    .Z(_00939_));
 MUX2_X1 _09862_ (.A(\samples_imag[5][7] ),
    .B(\samples_imag[7][7] ),
    .S(_00935_),
    .Z(_00940_));
 MUX2_X1 _09863_ (.A(_00939_),
    .B(_00940_),
    .S(_00899_),
    .Z(_00941_));
 MUX2_X2 _09864_ (.A(_00938_),
    .B(_00941_),
    .S(_00901_),
    .Z(_08599_));
 BUF_X8 _09865_ (.A(_00873_),
    .Z(_00942_));
 MUX2_X1 _09866_ (.A(\samples_imag[0][6] ),
    .B(\samples_imag[2][6] ),
    .S(_00942_),
    .Z(_00943_));
 MUX2_X1 _09867_ (.A(\samples_imag[1][6] ),
    .B(\samples_imag[3][6] ),
    .S(_00891_),
    .Z(_00944_));
 MUX2_X1 _09868_ (.A(_00943_),
    .B(_00944_),
    .S(_00894_),
    .Z(_00945_));
 MUX2_X1 _09869_ (.A(\samples_imag[4][6] ),
    .B(\samples_imag[6][6] ),
    .S(_00891_),
    .Z(_00946_));
 MUX2_X1 _09870_ (.A(\samples_imag[5][6] ),
    .B(\samples_imag[7][6] ),
    .S(_00891_),
    .Z(_00947_));
 MUX2_X1 _09871_ (.A(_00946_),
    .B(_00947_),
    .S(_00894_),
    .Z(_00948_));
 MUX2_X2 _09872_ (.A(_00945_),
    .B(_00948_),
    .S(_00901_),
    .Z(_08604_));
 MUX2_X1 _09873_ (.A(\samples_imag[0][5] ),
    .B(\samples_imag[2][5] ),
    .S(_00906_),
    .Z(_00949_));
 MUX2_X1 _09874_ (.A(\samples_imag[1][5] ),
    .B(\samples_imag[3][5] ),
    .S(_00906_),
    .Z(_00950_));
 MUX2_X1 _09875_ (.A(_00949_),
    .B(_00950_),
    .S(_00877_),
    .Z(_00951_));
 MUX2_X1 _09876_ (.A(\samples_imag[4][5] ),
    .B(\samples_imag[6][5] ),
    .S(_00906_),
    .Z(_00952_));
 MUX2_X1 _09877_ (.A(\samples_imag[5][5] ),
    .B(\samples_imag[7][5] ),
    .S(_00874_),
    .Z(_00953_));
 MUX2_X1 _09878_ (.A(_00952_),
    .B(_00953_),
    .S(_00877_),
    .Z(_00954_));
 MUX2_X2 _09879_ (.A(_00951_),
    .B(_00954_),
    .S(_00882_),
    .Z(_08609_));
 MUX2_X1 _09880_ (.A(\samples_imag[0][4] ),
    .B(\samples_imag[2][4] ),
    .S(_00896_),
    .Z(_00955_));
 MUX2_X1 _09881_ (.A(\samples_imag[1][4] ),
    .B(\samples_imag[3][4] ),
    .S(_00896_),
    .Z(_00956_));
 MUX2_X1 _09882_ (.A(_00955_),
    .B(_00956_),
    .S(_00899_),
    .Z(_00957_));
 MUX2_X1 _09883_ (.A(\samples_imag[4][4] ),
    .B(\samples_imag[6][4] ),
    .S(_00896_),
    .Z(_00958_));
 MUX2_X1 _09884_ (.A(\samples_imag[5][4] ),
    .B(\samples_imag[7][4] ),
    .S(_00935_),
    .Z(_00959_));
 MUX2_X1 _09885_ (.A(_00958_),
    .B(_00959_),
    .S(_00899_),
    .Z(_00960_));
 MUX2_X2 _09886_ (.A(_00957_),
    .B(_00960_),
    .S(_00901_),
    .Z(_08614_));
 MUX2_X1 _09887_ (.A(\samples_imag[0][3] ),
    .B(\samples_imag[2][3] ),
    .S(_00942_),
    .Z(_00961_));
 MUX2_X1 _09888_ (.A(\samples_imag[1][3] ),
    .B(\samples_imag[3][3] ),
    .S(_00942_),
    .Z(_00962_));
 MUX2_X1 _09889_ (.A(_00961_),
    .B(_00962_),
    .S(_00894_),
    .Z(_00963_));
 MUX2_X1 _09890_ (.A(\samples_imag[4][3] ),
    .B(\samples_imag[6][3] ),
    .S(_00942_),
    .Z(_00964_));
 MUX2_X1 _09891_ (.A(\samples_imag[5][3] ),
    .B(\samples_imag[7][3] ),
    .S(_00942_),
    .Z(_00965_));
 MUX2_X1 _09892_ (.A(_00964_),
    .B(_00965_),
    .S(_00894_),
    .Z(_00966_));
 MUX2_X2 _09893_ (.A(_00963_),
    .B(_00966_),
    .S(_00901_),
    .Z(_08619_));
 MUX2_X1 _09894_ (.A(\samples_imag[0][2] ),
    .B(\samples_imag[2][2] ),
    .S(_00883_),
    .Z(_00967_));
 MUX2_X1 _09895_ (.A(\samples_imag[1][2] ),
    .B(\samples_imag[3][2] ),
    .S(_00902_),
    .Z(_00968_));
 MUX2_X1 _09896_ (.A(_00967_),
    .B(_00968_),
    .S(_00886_),
    .Z(_00969_));
 MUX2_X1 _09897_ (.A(\samples_imag[4][2] ),
    .B(\samples_imag[6][2] ),
    .S(_00902_),
    .Z(_00970_));
 MUX2_X1 _09898_ (.A(\samples_imag[5][2] ),
    .B(\samples_imag[7][2] ),
    .S(_00902_),
    .Z(_00971_));
 MUX2_X1 _09899_ (.A(_00970_),
    .B(_00971_),
    .S(_00886_),
    .Z(_00972_));
 MUX2_X2 _09900_ (.A(_00969_),
    .B(_00972_),
    .S(_00882_),
    .Z(_08624_));
 MUX2_X1 _09901_ (.A(\samples_imag[0][1] ),
    .B(\samples_imag[2][1] ),
    .S(_00919_),
    .Z(_00973_));
 MUX2_X1 _09902_ (.A(\samples_imag[1][1] ),
    .B(\samples_imag[3][1] ),
    .S(_00919_),
    .Z(_00974_));
 MUX2_X1 _09903_ (.A(_00973_),
    .B(_00974_),
    .S(_00923_),
    .Z(_00975_));
 MUX2_X1 _09904_ (.A(\samples_imag[4][1] ),
    .B(\samples_imag[6][1] ),
    .S(_00919_),
    .Z(_00976_));
 MUX2_X1 _09905_ (.A(\samples_imag[5][1] ),
    .B(\samples_imag[7][1] ),
    .S(_00919_),
    .Z(_00977_));
 MUX2_X1 _09906_ (.A(_00976_),
    .B(_00977_),
    .S(_00923_),
    .Z(_00978_));
 MUX2_X2 _09907_ (.A(_00975_),
    .B(_00978_),
    .S(_00918_),
    .Z(_08629_));
 MUX2_X1 _09908_ (.A(\samples_imag[0][0] ),
    .B(\samples_imag[2][0] ),
    .S(net511),
    .Z(_00979_));
 MUX2_X1 _09909_ (.A(\samples_imag[1][0] ),
    .B(\samples_imag[3][0] ),
    .S(net511),
    .Z(_00980_));
 MUX2_X1 _09910_ (.A(_00979_),
    .B(_00980_),
    .S(_00913_),
    .Z(_00981_));
 MUX2_X1 _09911_ (.A(\samples_imag[4][0] ),
    .B(\samples_imag[6][0] ),
    .S(net511),
    .Z(_00982_));
 MUX2_X1 _09912_ (.A(\samples_imag[5][0] ),
    .B(\samples_imag[7][0] ),
    .S(_00910_),
    .Z(_00983_));
 MUX2_X1 _09913_ (.A(_00982_),
    .B(_00983_),
    .S(_00913_),
    .Z(_00984_));
 MUX2_X2 _09914_ (.A(_00981_),
    .B(_00984_),
    .S(_00918_),
    .Z(_08559_));
 MUX2_X1 _09915_ (.A(\samples_real[0][15] ),
    .B(\samples_real[2][15] ),
    .S(net56),
    .Z(_00985_));
 MUX2_X1 _09916_ (.A(\samples_real[1][15] ),
    .B(\samples_real[3][15] ),
    .S(net61),
    .Z(_00986_));
 MUX2_X1 _09917_ (.A(_00985_),
    .B(_00986_),
    .S(_00867_),
    .Z(_00987_));
 MUX2_X1 _09918_ (.A(\samples_real[4][15] ),
    .B(\samples_real[6][15] ),
    .S(net61),
    .Z(_00988_));
 MUX2_X1 _09919_ (.A(\samples_real[5][15] ),
    .B(\samples_real[7][15] ),
    .S(net61),
    .Z(_00989_));
 MUX2_X1 _09920_ (.A(_00988_),
    .B(_00989_),
    .S(_00867_),
    .Z(_00990_));
 MUX2_X2 _09921_ (.A(_00987_),
    .B(_00990_),
    .S(_00872_),
    .Z(_08642_));
 MUX2_X1 _09922_ (.A(\samples_real[0][14] ),
    .B(\samples_real[2][14] ),
    .S(_00874_),
    .Z(_00991_));
 MUX2_X1 _09923_ (.A(\samples_real[1][14] ),
    .B(\samples_real[3][14] ),
    .S(_00874_),
    .Z(_00992_));
 MUX2_X1 _09924_ (.A(_00991_),
    .B(_00992_),
    .S(_00877_),
    .Z(_00993_));
 MUX2_X1 _09925_ (.A(\samples_real[4][14] ),
    .B(\samples_real[6][14] ),
    .S(_00874_),
    .Z(_00994_));
 MUX2_X1 _09926_ (.A(\samples_real[5][14] ),
    .B(\samples_real[7][14] ),
    .S(_00874_),
    .Z(_00995_));
 MUX2_X1 _09927_ (.A(_00994_),
    .B(_00995_),
    .S(_00877_),
    .Z(_00996_));
 MUX2_X2 _09928_ (.A(_00993_),
    .B(_00996_),
    .S(_00882_),
    .Z(_08634_));
 MUX2_X1 _09929_ (.A(\samples_real[0][13] ),
    .B(\samples_real[2][13] ),
    .S(_00883_),
    .Z(_00997_));
 MUX2_X1 _09930_ (.A(\samples_real[1][13] ),
    .B(\samples_real[3][13] ),
    .S(_00883_),
    .Z(_00998_));
 MUX2_X1 _09931_ (.A(_00997_),
    .B(_00998_),
    .S(_00886_),
    .Z(_00999_));
 MUX2_X1 _09932_ (.A(\samples_real[4][13] ),
    .B(\samples_real[6][13] ),
    .S(_00883_),
    .Z(_01000_));
 MUX2_X1 _09933_ (.A(\samples_real[5][13] ),
    .B(\samples_real[7][13] ),
    .S(_00883_),
    .Z(_01001_));
 MUX2_X1 _09934_ (.A(_01000_),
    .B(_01001_),
    .S(_00886_),
    .Z(_01002_));
 MUX2_X2 _09935_ (.A(_00999_),
    .B(_01002_),
    .S(_00882_),
    .Z(_08650_));
 MUX2_X1 _09936_ (.A(\samples_real[0][12] ),
    .B(\samples_real[2][12] ),
    .S(_00891_),
    .Z(_01003_));
 MUX2_X1 _09937_ (.A(\samples_real[1][12] ),
    .B(\samples_real[3][12] ),
    .S(_00891_),
    .Z(_01004_));
 MUX2_X1 _09938_ (.A(_01003_),
    .B(_01004_),
    .S(_00894_),
    .Z(_01005_));
 MUX2_X1 _09939_ (.A(\samples_real[4][12] ),
    .B(\samples_real[6][12] ),
    .S(_00896_),
    .Z(_01006_));
 MUX2_X1 _09940_ (.A(\samples_real[5][12] ),
    .B(\samples_real[7][12] ),
    .S(_00896_),
    .Z(_01007_));
 MUX2_X1 _09941_ (.A(_01006_),
    .B(_01007_),
    .S(_00899_),
    .Z(_01008_));
 MUX2_X2 _09942_ (.A(_01005_),
    .B(_01008_),
    .S(_00901_),
    .Z(_08655_));
 MUX2_X1 _09943_ (.A(\samples_real[0][11] ),
    .B(\samples_real[2][11] ),
    .S(net59),
    .Z(_01009_));
 MUX2_X1 _09944_ (.A(\samples_real[1][11] ),
    .B(\samples_real[3][11] ),
    .S(net59),
    .Z(_01010_));
 MUX2_X1 _09945_ (.A(_01009_),
    .B(_01010_),
    .S(_00886_),
    .Z(_01011_));
 MUX2_X1 _09946_ (.A(\samples_real[4][11] ),
    .B(\samples_real[6][11] ),
    .S(_00906_),
    .Z(_01012_));
 MUX2_X1 _09947_ (.A(\samples_real[5][11] ),
    .B(\samples_real[7][11] ),
    .S(_00906_),
    .Z(_01013_));
 MUX2_X1 _09948_ (.A(_01012_),
    .B(_01013_),
    .S(_00877_),
    .Z(_01014_));
 MUX2_X2 _09949_ (.A(_01011_),
    .B(_01014_),
    .S(_00882_),
    .Z(_08660_));
 MUX2_X1 _09950_ (.A(\samples_real[0][10] ),
    .B(\samples_real[2][10] ),
    .S(net129),
    .Z(_01015_));
 MUX2_X1 _09951_ (.A(\samples_real[1][10] ),
    .B(\samples_real[3][10] ),
    .S(net129),
    .Z(_01016_));
 MUX2_X1 _09952_ (.A(_01015_),
    .B(_01016_),
    .S(_00913_),
    .Z(_01017_));
 MUX2_X1 _09953_ (.A(\samples_real[4][10] ),
    .B(\samples_real[6][10] ),
    .S(net129),
    .Z(_01018_));
 MUX2_X1 _09954_ (.A(\samples_real[5][10] ),
    .B(\samples_real[7][10] ),
    .S(net129),
    .Z(_01019_));
 MUX2_X1 _09955_ (.A(_01018_),
    .B(_01019_),
    .S(_00913_),
    .Z(_01020_));
 MUX2_X2 _09956_ (.A(_01017_),
    .B(_01020_),
    .S(_00918_),
    .Z(_08665_));
 MUX2_X1 _09957_ (.A(\samples_real[0][9] ),
    .B(\samples_real[2][9] ),
    .S(net60),
    .Z(_01021_));
 MUX2_X1 _09958_ (.A(\samples_real[1][9] ),
    .B(\samples_real[3][9] ),
    .S(_00921_),
    .Z(_01022_));
 MUX2_X1 _09959_ (.A(_01021_),
    .B(_01022_),
    .S(_00923_),
    .Z(_01023_));
 MUX2_X1 _09960_ (.A(\samples_real[4][9] ),
    .B(\samples_real[6][9] ),
    .S(_00921_),
    .Z(_01024_));
 MUX2_X1 _09961_ (.A(\samples_real[5][9] ),
    .B(\samples_real[7][9] ),
    .S(_00921_),
    .Z(_01025_));
 MUX2_X1 _09962_ (.A(_01024_),
    .B(_01025_),
    .S(_00923_),
    .Z(_01026_));
 MUX2_X2 _09963_ (.A(_01023_),
    .B(_01026_),
    .S(_00918_),
    .Z(_08670_));
 MUX2_X1 _09964_ (.A(\samples_real[0][8] ),
    .B(\samples_real[2][8] ),
    .S(_00921_),
    .Z(_01027_));
 MUX2_X1 _09965_ (.A(\samples_real[1][8] ),
    .B(\samples_real[3][8] ),
    .S(_00921_),
    .Z(_01028_));
 MUX2_X1 _09966_ (.A(_01027_),
    .B(_01028_),
    .S(_00923_),
    .Z(_01029_));
 MUX2_X1 _09967_ (.A(\samples_real[4][8] ),
    .B(\samples_real[6][8] ),
    .S(net477),
    .Z(_01030_));
 MUX2_X1 _09968_ (.A(\samples_real[5][8] ),
    .B(\samples_real[7][8] ),
    .S(net477),
    .Z(_01031_));
 MUX2_X1 _09969_ (.A(_01030_),
    .B(_01031_),
    .S(_00913_),
    .Z(_01032_));
 MUX2_X2 _09970_ (.A(_01029_),
    .B(_01032_),
    .S(_00918_),
    .Z(_08675_));
 MUX2_X1 _09971_ (.A(\samples_real[0][7] ),
    .B(\samples_real[2][7] ),
    .S(_00935_),
    .Z(_01033_));
 MUX2_X1 _09972_ (.A(\samples_real[1][7] ),
    .B(\samples_real[3][7] ),
    .S(_00935_),
    .Z(_01034_));
 MUX2_X1 _09973_ (.A(_01033_),
    .B(_01034_),
    .S(_00899_),
    .Z(_01035_));
 MUX2_X1 _09974_ (.A(\samples_real[4][7] ),
    .B(\samples_real[6][7] ),
    .S(_00935_),
    .Z(_01036_));
 MUX2_X1 _09975_ (.A(\samples_real[5][7] ),
    .B(\samples_real[7][7] ),
    .S(_00935_),
    .Z(_01037_));
 MUX2_X1 _09976_ (.A(_01036_),
    .B(_01037_),
    .S(_00899_),
    .Z(_01038_));
 MUX2_X2 _09977_ (.A(_01035_),
    .B(_01038_),
    .S(_00901_),
    .Z(_08680_));
 MUX2_X1 _09978_ (.A(\samples_real[0][6] ),
    .B(\samples_real[2][6] ),
    .S(_00942_),
    .Z(_01039_));
 MUX2_X1 _09979_ (.A(\samples_real[1][6] ),
    .B(\samples_real[3][6] ),
    .S(_00891_),
    .Z(_01040_));
 MUX2_X1 _09980_ (.A(_01039_),
    .B(_01040_),
    .S(_00894_),
    .Z(_01041_));
 MUX2_X1 _09981_ (.A(\samples_real[4][6] ),
    .B(\samples_real[6][6] ),
    .S(_00891_),
    .Z(_01042_));
 MUX2_X1 _09982_ (.A(\samples_real[5][6] ),
    .B(\samples_real[7][6] ),
    .S(_00891_),
    .Z(_01043_));
 MUX2_X1 _09983_ (.A(_01042_),
    .B(_01043_),
    .S(_00894_),
    .Z(_01044_));
 MUX2_X2 _09984_ (.A(_01041_),
    .B(_01044_),
    .S(_00901_),
    .Z(_08685_));
 MUX2_X1 _09985_ (.A(\samples_real[0][5] ),
    .B(\samples_real[2][5] ),
    .S(_00906_),
    .Z(_01045_));
 MUX2_X1 _09986_ (.A(\samples_real[1][5] ),
    .B(\samples_real[3][5] ),
    .S(_00906_),
    .Z(_01046_));
 MUX2_X1 _09987_ (.A(_01045_),
    .B(_01046_),
    .S(_00877_),
    .Z(_01047_));
 MUX2_X1 _09988_ (.A(\samples_real[4][5] ),
    .B(\samples_real[6][5] ),
    .S(_00906_),
    .Z(_01048_));
 MUX2_X1 _09989_ (.A(\samples_real[5][5] ),
    .B(\samples_real[7][5] ),
    .S(_00874_),
    .Z(_01049_));
 MUX2_X1 _09990_ (.A(_01048_),
    .B(_01049_),
    .S(_00877_),
    .Z(_01050_));
 MUX2_X2 _09991_ (.A(_01047_),
    .B(_01050_),
    .S(_00882_),
    .Z(_08690_));
 MUX2_X1 _09992_ (.A(\samples_real[0][4] ),
    .B(\samples_real[2][4] ),
    .S(_00896_),
    .Z(_01051_));
 MUX2_X1 _09993_ (.A(\samples_real[1][4] ),
    .B(\samples_real[3][4] ),
    .S(_00896_),
    .Z(_01052_));
 MUX2_X1 _09994_ (.A(_01051_),
    .B(_01052_),
    .S(_00899_),
    .Z(_01053_));
 MUX2_X1 _09995_ (.A(\samples_real[4][4] ),
    .B(\samples_real[6][4] ),
    .S(_00896_),
    .Z(_01054_));
 MUX2_X1 _09996_ (.A(\samples_real[5][4] ),
    .B(\samples_real[7][4] ),
    .S(_00935_),
    .Z(_01055_));
 MUX2_X1 _09997_ (.A(_01054_),
    .B(_01055_),
    .S(_00899_),
    .Z(_01056_));
 MUX2_X2 _09998_ (.A(_01053_),
    .B(_01056_),
    .S(_00901_),
    .Z(_08695_));
 MUX2_X1 _09999_ (.A(\samples_real[0][3] ),
    .B(\samples_real[2][3] ),
    .S(_00942_),
    .Z(_01057_));
 MUX2_X1 _10000_ (.A(\samples_real[1][3] ),
    .B(\samples_real[3][3] ),
    .S(_00942_),
    .Z(_01058_));
 MUX2_X1 _10001_ (.A(_01057_),
    .B(_01058_),
    .S(_00894_),
    .Z(_01059_));
 MUX2_X1 _10002_ (.A(\samples_real[4][3] ),
    .B(\samples_real[6][3] ),
    .S(_00942_),
    .Z(_01060_));
 MUX2_X1 _10003_ (.A(\samples_real[5][3] ),
    .B(\samples_real[7][3] ),
    .S(_00942_),
    .Z(_01061_));
 MUX2_X1 _10004_ (.A(_01060_),
    .B(_01061_),
    .S(_00894_),
    .Z(_01062_));
 MUX2_X2 _10005_ (.A(_01059_),
    .B(_01062_),
    .S(_00901_),
    .Z(_08700_));
 MUX2_X1 _10006_ (.A(\samples_real[0][2] ),
    .B(\samples_real[2][2] ),
    .S(_00883_),
    .Z(_01063_));
 MUX2_X1 _10007_ (.A(\samples_real[1][2] ),
    .B(\samples_real[3][2] ),
    .S(_00902_),
    .Z(_01064_));
 MUX2_X1 _10008_ (.A(_01063_),
    .B(_01064_),
    .S(_00886_),
    .Z(_01065_));
 MUX2_X1 _10009_ (.A(\samples_real[4][2] ),
    .B(\samples_real[6][2] ),
    .S(net59),
    .Z(_01066_));
 MUX2_X1 _10010_ (.A(\samples_real[5][2] ),
    .B(\samples_real[7][2] ),
    .S(_00902_),
    .Z(_01067_));
 MUX2_X1 _10011_ (.A(_01066_),
    .B(_01067_),
    .S(_00886_),
    .Z(_01068_));
 MUX2_X2 _10012_ (.A(_01065_),
    .B(_01068_),
    .S(_00882_),
    .Z(_08705_));
 MUX2_X1 _10013_ (.A(\samples_real[0][1] ),
    .B(\samples_real[2][1] ),
    .S(net60),
    .Z(_01069_));
 MUX2_X1 _10014_ (.A(\samples_real[1][1] ),
    .B(\samples_real[3][1] ),
    .S(net60),
    .Z(_01070_));
 MUX2_X1 _10015_ (.A(_01069_),
    .B(_01070_),
    .S(_00923_),
    .Z(_01071_));
 MUX2_X1 _10016_ (.A(\samples_real[4][1] ),
    .B(\samples_real[6][1] ),
    .S(net60),
    .Z(_01072_));
 MUX2_X1 _10017_ (.A(\samples_real[5][1] ),
    .B(\samples_real[7][1] ),
    .S(_00919_),
    .Z(_01073_));
 MUX2_X1 _10018_ (.A(_01072_),
    .B(_01073_),
    .S(_00923_),
    .Z(_01074_));
 MUX2_X2 _10019_ (.A(_01071_),
    .B(_01074_),
    .S(_00918_),
    .Z(_08710_));
 MUX2_X1 _10020_ (.A(\samples_real[0][0] ),
    .B(\samples_real[2][0] ),
    .S(net130),
    .Z(_01075_));
 MUX2_X1 _10021_ (.A(\samples_real[1][0] ),
    .B(\samples_real[3][0] ),
    .S(_00931_),
    .Z(_01076_));
 MUX2_X1 _10022_ (.A(_01075_),
    .B(_01076_),
    .S(_00913_),
    .Z(_01077_));
 MUX2_X1 _10023_ (.A(\samples_real[4][0] ),
    .B(\samples_real[6][0] ),
    .S(_00931_),
    .Z(_01078_));
 MUX2_X1 _10024_ (.A(\samples_real[5][0] ),
    .B(\samples_real[7][0] ),
    .S(_00910_),
    .Z(_01079_));
 MUX2_X1 _10025_ (.A(_01078_),
    .B(_01079_),
    .S(_00913_),
    .Z(_01080_));
 MUX2_X2 _10026_ (.A(_01077_),
    .B(_01080_),
    .S(_00918_),
    .Z(_08640_));
 INV_X4 _10027_ (.A(_00847_),
    .ZN(_01081_));
 BUF_X4 _10028_ (.A(_09363_),
    .Z(_01082_));
 NAND2_X4 _10029_ (.A1(_01082_),
    .A2(_01081_),
    .ZN(_08715_));
 BUF_X4 _10030_ (.A(_09367_),
    .Z(_01083_));
 NAND2_X4 _10031_ (.A1(_00847_),
    .A2(_01083_),
    .ZN(_08777_));
 INV_X1 _10032_ (.A(_08777_),
    .ZN(_09313_));
 BUF_X4 _10033_ (.A(_09369_),
    .Z(_01084_));
 NAND2_X4 _10034_ (.A1(_00848_),
    .A2(_01084_),
    .ZN(_08764_));
 INV_X1 _10035_ (.A(_08764_),
    .ZN(_09317_));
 NAND2_X4 _10036_ (.A1(_00848_),
    .A2(_01082_),
    .ZN(_08743_));
 INV_X1 _10037_ (.A(_08743_),
    .ZN(_09321_));
 NAND2_X4 _10038_ (.A1(_09340_),
    .A2(_01083_),
    .ZN(_08721_));
 INV_X2 _10039_ (.A(_08721_),
    .ZN(_09329_));
 NAND2_X4 _10040_ (.A1(_09340_),
    .A2(_01084_),
    .ZN(_07367_));
 INV_X2 _10041_ (.A(_07367_),
    .ZN(_07363_));
 BUF_X4 _10042_ (.A(_09345_),
    .Z(_01085_));
 INV_X4 _10043_ (.A(_01085_),
    .ZN(_01086_));
 BUF_X4 _10044_ (.A(_01086_),
    .Z(_01087_));
 CLKBUF_X3 _10045_ (.A(_01087_),
    .Z(_01088_));
 CLKBUF_X3 _10046_ (.A(_01088_),
    .Z(_01089_));
 BUF_X4 _10047_ (.A(_01089_),
    .Z(_01090_));
 BUF_X4 _10048_ (.A(_01090_),
    .Z(_01091_));
 BUF_X8 _10049_ (.A(_01091_),
    .Z(_08819_));
 INV_X1 _10050_ (.A(_01082_),
    .ZN(_01092_));
 OAI22_X1 _10051_ (.A1(_00847_),
    .A2(_09340_),
    .B1(_01083_),
    .B2(_01084_),
    .ZN(_01093_));
 BUF_X2 _10052_ (.A(_09342_),
    .Z(_01094_));
 BUF_X4 _10053_ (.A(_00040_),
    .Z(_01095_));
 BUF_X4 _10054_ (.A(_09357_),
    .Z(_01096_));
 NAND2_X4 _10055_ (.A1(_01095_),
    .A2(_01096_),
    .ZN(_01097_));
 BUF_X4 _10056_ (.A(_09309_),
    .Z(_01098_));
 OR2_X4 _10057_ (.A1(_09325_),
    .A2(_01098_),
    .ZN(_01099_));
 OAI22_X4 _10058_ (.A1(_01094_),
    .A2(_01085_),
    .B1(_01099_),
    .B2(_01097_),
    .ZN(_01100_));
 AND4_X4 _10059_ (.A1(_01092_),
    .A2(_08717_),
    .A3(_01093_),
    .A4(_01100_),
    .ZN(_08718_));
 INV_X2 _10060_ (.A(net42),
    .ZN(_09286_));
 NOR3_X1 _10061_ (.A1(_01082_),
    .A2(_01083_),
    .A3(_01084_),
    .ZN(_01101_));
 OAI21_X2 _10062_ (.A(_01086_),
    .B1(_01101_),
    .B2(_01081_),
    .ZN(_01102_));
 AOI21_X4 _10063_ (.A(_01094_),
    .B1(_01083_),
    .B2(_09340_),
    .ZN(_01103_));
 INV_X1 _10064_ (.A(_01103_),
    .ZN(_01104_));
 OAI21_X2 _10065_ (.A(_08720_),
    .B1(_01092_),
    .B2(_00847_),
    .ZN(_01105_));
 NOR3_X2 clone22 (.A1(_04633_),
    .A2(_04647_),
    .A3(_04634_),
    .ZN(net22));
 INV_X2 _10067_ (.A(_08719_),
    .ZN(_01107_));
 AOI211_X2 _10068_ (.A(_01102_),
    .B(_01104_),
    .C1(_01107_),
    .C2(_01105_),
    .ZN(_01108_));
 BUF_X4 _10069_ (.A(\butterfly_count[2] ),
    .Z(_01109_));
 OR2_X2 _10070_ (.A1(_01095_),
    .A2(_01109_),
    .ZN(_01110_));
 INV_X2 _10071_ (.A(_01096_),
    .ZN(_01111_));
 AOI21_X2 _10072_ (.A(_01110_),
    .B1(_01111_),
    .B2(_01107_),
    .ZN(_01112_));
 MUX2_X1 _10073_ (.A(_01110_),
    .B(_01112_),
    .S(_08715_),
    .Z(_01113_));
 NAND2_X4 _10074_ (.A1(net383),
    .A2(_01113_),
    .ZN(_01114_));
 INV_X2 _10075_ (.A(_01114_),
    .ZN(_08725_));
 BUF_X4 _10076_ (.A(net31),
    .Z(_01115_));
 BUF_X4 _10077_ (.A(_01115_),
    .Z(_01116_));
 BUF_X4 _10078_ (.A(_01116_),
    .Z(_01117_));
 BUF_X4 _10079_ (.A(_01085_),
    .Z(_01118_));
 BUF_X4 _10080_ (.A(_01118_),
    .Z(_01119_));
 CLKBUF_X3 _10081_ (.A(_01119_),
    .Z(_01120_));
 BUF_X4 _10082_ (.A(_01120_),
    .Z(_01121_));
 CLKBUF_X3 _10083_ (.A(_01121_),
    .Z(_01122_));
 INV_X1 _10084_ (.A(_09002_),
    .ZN(_01123_));
 INV_X1 _10085_ (.A(_08996_),
    .ZN(_01124_));
 INV_X1 _10086_ (.A(_08990_),
    .ZN(_01125_));
 OAI21_X2 _10087_ (.A(_08991_),
    .B1(_08984_),
    .B2(_08985_),
    .ZN(_01126_));
 NAND2_X2 _10088_ (.A1(_01126_),
    .A2(_01125_),
    .ZN(_01127_));
 AND2_X4 _10089_ (.A1(_08988_),
    .A2(_01127_),
    .ZN(_01128_));
 OAI21_X4 _10090_ (.A(_08997_),
    .B1(_01128_),
    .B2(_08987_),
    .ZN(_01129_));
 NAND2_X4 _10091_ (.A1(_01124_),
    .A2(_01129_),
    .ZN(_01130_));
 AOI21_X4 _10092_ (.A(_08993_),
    .B1(_08994_),
    .B2(_01130_),
    .ZN(_01131_));
 INV_X1 _10093_ (.A(_09003_),
    .ZN(_01132_));
 OAI21_X4 _10094_ (.A(_01123_),
    .B1(_01131_),
    .B2(_01132_),
    .ZN(_01133_));
 AND2_X4 _10095_ (.A1(_09000_),
    .A2(_01133_),
    .ZN(_01134_));
 OR2_X4 _10096_ (.A1(_08999_),
    .A2(_01134_),
    .ZN(_01135_));
 NAND2_X1 _10097_ (.A1(_01122_),
    .A2(_01135_),
    .ZN(_01136_));
 NAND2_X1 _10098_ (.A1(_01117_),
    .A2(_01136_),
    .ZN(_01137_));
 AOI21_X4 clone6 (.A(_09201_),
    .B1(_03966_),
    .B2(_09202_),
    .ZN(net6));
 INV_X1 _10100_ (.A(_08967_),
    .ZN(_01139_));
 BUF_X2 _10101_ (.A(_08974_),
    .Z(_01140_));
 NAND2_X1 _10102_ (.A1(_01140_),
    .A2(_08977_),
    .ZN(_01141_));
 CLKBUF_X2 _10103_ (.A(_08983_),
    .Z(_01142_));
 INV_X1 _10104_ (.A(_01142_),
    .ZN(_01143_));
 OR3_X2 _10105_ (.A1(_01082_),
    .A2(_01083_),
    .A3(_01084_),
    .ZN(_01144_));
 AOI21_X4 _10106_ (.A(_01085_),
    .B1(_01144_),
    .B2(_00848_),
    .ZN(_01145_));
 INV_X1 _10107_ (.A(_08720_),
    .ZN(_01146_));
 AOI21_X2 _10108_ (.A(_01146_),
    .B1(_01082_),
    .B2(_01081_),
    .ZN(_01147_));
 OAI211_X4 _10109_ (.A(_01145_),
    .B(_01103_),
    .C1(_01147_),
    .C2(_08719_),
    .ZN(_01148_));
 AND2_X2 _10110_ (.A1(_01095_),
    .A2(_01109_),
    .ZN(_01149_));
 BUF_X4 _10111_ (.A(_01149_),
    .Z(_01150_));
 NAND2_X1 _10112_ (.A1(_01148_),
    .A2(_01150_),
    .ZN(_01151_));
 INV_X1 _10113_ (.A(_01098_),
    .ZN(_01152_));
 BUF_X4 _10114_ (.A(_01152_),
    .Z(_01153_));
 INV_X1 _10115_ (.A(_08733_),
    .ZN(_01154_));
 OR2_X1 _10116_ (.A1(_08742_),
    .A2(_08741_),
    .ZN(_01155_));
 AND2_X2 _10117_ (.A1(_08736_),
    .A2(_08739_),
    .ZN(_01156_));
 AOI221_X2 _10118_ (.A(_08735_),
    .B1(_01155_),
    .B2(_01156_),
    .C1(_08738_),
    .C2(_08736_),
    .ZN(_01157_));
 NOR2_X4 _10119_ (.A1(_01154_),
    .A2(_01157_),
    .ZN(_01158_));
 OAI21_X4 _10120_ (.A(_01145_),
    .B1(_01158_),
    .B2(_08732_),
    .ZN(_01159_));
 INV_X16 _10121_ (.A(_09325_),
    .ZN(_08730_));
 INV_X1 _10122_ (.A(_08724_),
    .ZN(_01160_));
 OAI21_X2 _10123_ (.A(_08727_),
    .B1(_08729_),
    .B2(_08728_),
    .ZN(_01161_));
 INV_X1 _10124_ (.A(_08726_),
    .ZN(_01162_));
 AOI21_X4 _10125_ (.A(_01160_),
    .B1(_01161_),
    .B2(_01162_),
    .ZN(_01163_));
 OAI211_X4 _10126_ (.A(_08730_),
    .B(_01145_),
    .C1(_01163_),
    .C2(_08723_),
    .ZN(_01164_));
 INV_X1 _10127_ (.A(_01164_),
    .ZN(_01165_));
 NOR2_X1 _10128_ (.A1(_08726_),
    .A2(_08724_),
    .ZN(_01166_));
 AOI21_X2 _10129_ (.A(_01163_),
    .B1(_01166_),
    .B2(_01161_),
    .ZN(_01167_));
 NAND3_X2 _10130_ (.A1(_01159_),
    .A2(_01165_),
    .A3(_01167_),
    .ZN(_01168_));
 INV_X2 _10131_ (.A(_01109_),
    .ZN(_01169_));
 NAND2_X4 _10132_ (.A1(_01169_),
    .A2(_01096_),
    .ZN(_01170_));
 NOR2_X2 _10133_ (.A1(_01098_),
    .A2(_01170_),
    .ZN(_01171_));
 NAND4_X1 _10134_ (.A1(_08724_),
    .A2(_08727_),
    .A3(_08730_),
    .A4(_08729_),
    .ZN(_01172_));
 AOI21_X2 _10135_ (.A(_01172_),
    .B1(_01144_),
    .B2(_00848_),
    .ZN(_01173_));
 NOR2_X4 _10136_ (.A1(_01112_),
    .A2(_01149_),
    .ZN(_01174_));
 OAI211_X4 _10137_ (.A(_01171_),
    .B(_01173_),
    .C1(_01148_),
    .C2(_01174_),
    .ZN(_01175_));
 XOR2_X1 _10138_ (.A(_08716_),
    .B(_08720_),
    .Z(_01176_));
 OR4_X4 _10139_ (.A1(_08719_),
    .A2(_01109_),
    .A3(_01095_),
    .A4(_01096_),
    .ZN(_01177_));
 NAND2_X2 _10140_ (.A1(_01177_),
    .A2(_01103_),
    .ZN(_01178_));
 AOI211_X4 _10141_ (.A(_01178_),
    .B(_01102_),
    .C1(_01105_),
    .C2(_01107_),
    .ZN(_01179_));
 MUX2_X2 _10142_ (.A(_08718_),
    .B(_01176_),
    .S(_01179_),
    .Z(_08722_));
 NAND4_X4 _10143_ (.A1(_01159_),
    .A2(_01164_),
    .A3(_01175_),
    .A4(_08722_),
    .ZN(_01180_));
 NOR2_X2 _10144_ (.A1(_01085_),
    .A2(_09313_),
    .ZN(_01181_));
 INV_X1 _10145_ (.A(_01181_),
    .ZN(_01182_));
 INV_X1 _10146_ (.A(_08767_),
    .ZN(_01183_));
 BUF_X2 _10147_ (.A(_08770_),
    .Z(_01184_));
 AOI21_X2 _10148_ (.A(_08769_),
    .B1(_08772_),
    .B2(_01184_),
    .ZN(_01185_));
 NAND3_X2 _10149_ (.A1(_08767_),
    .A2(_01184_),
    .A3(_08773_),
    .ZN(_01186_));
 BUF_X1 _10150_ (.A(_08760_),
    .Z(_01187_));
 NAND3_X4 clone8 (.A1(net12),
    .A2(_03926_),
    .A3(_03910_),
    .ZN(net8));
 BUF_X1 _10152_ (.A(_08763_),
    .Z(_01189_));
 OAI211_X2 _10153_ (.A(_08776_),
    .B(_01187_),
    .C1(_08762_),
    .C2(_01189_),
    .ZN(_01190_));
 AOI21_X2 _10154_ (.A(_08775_),
    .B1(_08776_),
    .B2(_08759_),
    .ZN(_01191_));
 AND2_X4 _10155_ (.A1(_01191_),
    .A2(_01190_),
    .ZN(_01192_));
 OAI22_X4 _10156_ (.A1(_01183_),
    .A2(_01185_),
    .B1(_01192_),
    .B2(_01186_),
    .ZN(_01193_));
 INV_X1 _10157_ (.A(_08773_),
    .ZN(_01194_));
 AOI21_X2 _10158_ (.A(_01194_),
    .B1(_01191_),
    .B2(_01190_),
    .ZN(_01195_));
 NOR4_X4 _10159_ (.A1(_08767_),
    .A2(_08769_),
    .A3(_08772_),
    .A4(_01195_),
    .ZN(_01196_));
 NOR3_X2 _10160_ (.A1(_08767_),
    .A2(_01184_),
    .A3(_08769_),
    .ZN(_01197_));
 NOR4_X4 _10161_ (.A1(_01196_),
    .A2(_01193_),
    .A3(_01182_),
    .A4(_01197_),
    .ZN(_01198_));
 NAND3_X1 _10162_ (.A1(_01189_),
    .A2(_01187_),
    .A3(_08776_),
    .ZN(_01199_));
 OR3_X4 _10163_ (.A1(_01186_),
    .A2(_01170_),
    .A3(_01199_),
    .ZN(_01200_));
 NOR2_X1 _10164_ (.A1(_01095_),
    .A2(_01109_),
    .ZN(_01201_));
 OAI21_X1 _10165_ (.A(_01201_),
    .B1(_01096_),
    .B2(_08719_),
    .ZN(_01202_));
 NAND2_X2 _10166_ (.A1(_01095_),
    .A2(_01109_),
    .ZN(_01203_));
 NAND2_X2 _10167_ (.A1(_01202_),
    .A2(_01203_),
    .ZN(_01204_));
 AOI21_X4 _10168_ (.A(_01200_),
    .B1(_01204_),
    .B2(net383),
    .ZN(_01205_));
 OAI21_X4 _10169_ (.A(_01198_),
    .B1(_08766_),
    .B2(_01205_),
    .ZN(_01206_));
 XNOR2_X1 _10170_ (.A(_08733_),
    .B(_01157_),
    .ZN(_01207_));
 NAND3_X2 _10171_ (.A1(_08732_),
    .A2(_01145_),
    .A3(_01207_),
    .ZN(_01208_));
 AOI21_X2 _10172_ (.A(_08751_),
    .B1(_08754_),
    .B2(_08752_),
    .ZN(_01209_));
 NAND2_X1 _10173_ (.A1(_08752_),
    .A2(_08755_),
    .ZN(_01210_));
 NOR2_X2 _10174_ (.A1(_08757_),
    .A2(_08756_),
    .ZN(_01211_));
 OAI21_X4 _10175_ (.A(_01209_),
    .B1(_01210_),
    .B2(_01211_),
    .ZN(_01212_));
 BUF_X2 _10176_ (.A(_08746_),
    .Z(_01213_));
 AND2_X2 _10177_ (.A1(_01213_),
    .A2(_08749_),
    .ZN(_01214_));
 AOI221_X2 _10178_ (.A(_08745_),
    .B1(_01212_),
    .B2(_01214_),
    .C1(_01213_),
    .C2(_08748_),
    .ZN(_01215_));
 OAI21_X2 _10179_ (.A(_00848_),
    .B1(_01083_),
    .B2(_01084_),
    .ZN(_01216_));
 NAND2_X2 _10180_ (.A1(_01086_),
    .A2(_01216_),
    .ZN(_01217_));
 OR2_X4 _10181_ (.A1(_01215_),
    .A2(_01217_),
    .ZN(_01218_));
 NAND3_X2 _10182_ (.A1(_01169_),
    .A2(_01152_),
    .A3(_01096_),
    .ZN(_01219_));
 AND2_X1 _10183_ (.A1(_08752_),
    .A2(_08755_),
    .ZN(_01220_));
 NAND4_X1 _10184_ (.A1(_08757_),
    .A2(_01220_),
    .A3(_01214_),
    .A4(_01216_),
    .ZN(_01221_));
 NOR2_X1 _10185_ (.A1(_01219_),
    .A2(_01221_),
    .ZN(_01222_));
 OAI21_X2 _10186_ (.A(_01222_),
    .B1(_01174_),
    .B2(_01148_),
    .ZN(_01223_));
 AND3_X1 _10187_ (.A1(_01208_),
    .A2(_01218_),
    .A3(_01223_),
    .ZN(_01224_));
 NAND4_X4 _10188_ (.A1(_01168_),
    .A2(_01180_),
    .A3(_01206_),
    .A4(_01224_),
    .ZN(_01225_));
 AOI21_X4 _10189_ (.A(_08748_),
    .B1(_08749_),
    .B2(_01212_),
    .ZN(_01226_));
 XNOR2_X2 _10190_ (.A(_01213_),
    .B(_01226_),
    .ZN(_01227_));
 AOI21_X4 _10191_ (.A(_01227_),
    .B1(_01223_),
    .B2(_01218_),
    .ZN(_01228_));
 OAI21_X4 _10192_ (.A(_01181_),
    .B1(_01193_),
    .B2(_08766_),
    .ZN(_01229_));
 INV_X4 _10193_ (.A(_01229_),
    .ZN(_01230_));
 OAI21_X4 _10194_ (.A(_01206_),
    .B1(_01228_),
    .B2(_01230_),
    .ZN(_01231_));
 NAND3_X4 _10195_ (.A1(_01153_),
    .A2(_01225_),
    .A3(_01231_),
    .ZN(_01232_));
 NAND3_X2 _10196_ (.A1(_08783_),
    .A2(_08789_),
    .A3(_08786_),
    .ZN(_01233_));
 BUF_X2 clone10 (.A(_01588_),
    .Z(net10));
 AOI21_X2 _10198_ (.A(_08791_),
    .B1(_08792_),
    .B2(_08794_),
    .ZN(_01235_));
 BUF_X1 _10199_ (.A(_08795_),
    .Z(_01236_));
 BUF_X4 _10200_ (.A(_08797_),
    .Z(_01237_));
 OAI211_X2 _10201_ (.A(_01236_),
    .B(_08792_),
    .C1(_08796_),
    .C2(_01237_),
    .ZN(_01238_));
 AOI21_X4 _10202_ (.A(_01233_),
    .B1(_01238_),
    .B2(_01235_),
    .ZN(_01239_));
 INV_X1 _10203_ (.A(_08783_),
    .ZN(_01240_));
 AOI21_X1 _10204_ (.A(_08785_),
    .B1(_08786_),
    .B2(_08788_),
    .ZN(_01241_));
 NOR2_X2 _10205_ (.A1(_01240_),
    .A2(_01241_),
    .ZN(_01242_));
 NOR4_X4 _10206_ (.A1(_01239_),
    .A2(_08779_),
    .A3(_01242_),
    .A4(_08782_),
    .ZN(_01243_));
 NAND3_X4 clone7 (.A1(_02124_),
    .A2(net15),
    .A3(_02125_),
    .ZN(net7));
 NOR2_X1 _10208_ (.A1(_08780_),
    .A2(_08779_),
    .ZN(_01245_));
 NOR3_X2 _10209_ (.A1(_01085_),
    .A2(_01243_),
    .A3(_01245_),
    .ZN(_01246_));
 AOI21_X2 _10210_ (.A(_01219_),
    .B1(_01204_),
    .B2(net383),
    .ZN(_01247_));
 INV_X1 _10211_ (.A(_01094_),
    .ZN(_01248_));
 NAND3_X1 _10212_ (.A1(_01248_),
    .A2(_08721_),
    .A3(_01149_),
    .ZN(_01249_));
 AOI211_X4 _10213_ (.A(_01102_),
    .B(_01249_),
    .C1(_01105_),
    .C2(_01107_),
    .ZN(_08740_));
 NAND4_X2 _10214_ (.A1(_01237_),
    .A2(_08780_),
    .A3(_08792_),
    .A4(_01236_),
    .ZN(_01250_));
 NOR3_X2 _10215_ (.A1(_01233_),
    .A2(_08740_),
    .A3(_01250_),
    .ZN(_01251_));
 AOI21_X4 _10216_ (.A(_01246_),
    .B1(_01247_),
    .B2(_01251_),
    .ZN(_01252_));
 INV_X1 _10217_ (.A(_08799_),
    .ZN(_01253_));
 INV_X1 _10218_ (.A(_08805_),
    .ZN(_01254_));
 AOI21_X2 _10219_ (.A(_08808_),
    .B1(_08811_),
    .B2(_08809_),
    .ZN(_01255_));
 INV_X1 _10220_ (.A(_08806_),
    .ZN(_01256_));
 OAI21_X4 _10221_ (.A(_01254_),
    .B1(_01256_),
    .B2(_01255_),
    .ZN(_01257_));
 INV_X4 _10222_ (.A(_01257_),
    .ZN(_01258_));
 AOI21_X1 _10223_ (.A(_08814_),
    .B1(_08817_),
    .B2(_08815_),
    .ZN(_01259_));
 NAND4_X2 _10224_ (.A1(_01148_),
    .A2(_01149_),
    .A3(_01258_),
    .A4(_01259_),
    .ZN(_01260_));
 INV_X1 _10225_ (.A(_08803_),
    .ZN(_01261_));
 AND2_X1 _10226_ (.A1(_08806_),
    .A2(_08809_),
    .ZN(_01262_));
 INV_X1 _10227_ (.A(_08812_),
    .ZN(_01263_));
 INV_X1 _10228_ (.A(_08814_),
    .ZN(_01264_));
 OAI21_X2 _10229_ (.A(_08815_),
    .B1(_08817_),
    .B2(_08818_),
    .ZN(_01265_));
 AOI21_X2 _10230_ (.A(_01263_),
    .B1(_01264_),
    .B2(_01265_),
    .ZN(_01266_));
 AOI21_X4 _10231_ (.A(_01257_),
    .B1(_01262_),
    .B2(_01266_),
    .ZN(_01267_));
 NOR2_X4 _10232_ (.A1(_01261_),
    .A2(_01267_),
    .ZN(_01268_));
 AOI21_X4 _10233_ (.A(_08802_),
    .B1(_01260_),
    .B2(_01268_),
    .ZN(_01269_));
 BUF_X1 _10234_ (.A(_08800_),
    .Z(_01270_));
 INV_X1 _10235_ (.A(_01270_),
    .ZN(_01271_));
 OAI21_X4 _10236_ (.A(_01253_),
    .B1(_01269_),
    .B2(_01271_),
    .ZN(_01272_));
 NAND2_X1 _10237_ (.A1(net31),
    .A2(_01206_),
    .ZN(_01273_));
 AND3_X4 _10238_ (.A1(_01252_),
    .A2(_01273_),
    .A3(_01272_),
    .ZN(_01274_));
 NAND2_X4 _10239_ (.A1(_01232_),
    .A2(_01274_),
    .ZN(_01275_));
 INV_X1 _10240_ (.A(_08780_),
    .ZN(_01276_));
 NOR3_X2 _10241_ (.A1(_08782_),
    .A2(_01239_),
    .A3(_01242_),
    .ZN(_01277_));
 NOR2_X1 _10242_ (.A1(_01276_),
    .A2(_01277_),
    .ZN(_01278_));
 AND2_X1 _10243_ (.A1(_01276_),
    .A2(_01277_),
    .ZN(_01279_));
 AND3_X2 _10244_ (.A1(net3),
    .A2(_01165_),
    .A3(_01167_),
    .ZN(_01280_));
 AND4_X2 _10245_ (.A1(net3),
    .A2(_01164_),
    .A3(_01175_),
    .A4(_08722_),
    .ZN(_01281_));
 OR4_X2 _10246_ (.A1(_01182_),
    .A2(_01193_),
    .A3(_01196_),
    .A4(_01197_),
    .ZN(_01282_));
 NOR3_X1 _10247_ (.A1(_01170_),
    .A2(_01186_),
    .A3(_01199_),
    .ZN(_01283_));
 OAI21_X2 _10248_ (.A(_01283_),
    .B1(_01174_),
    .B2(_01148_),
    .ZN(_01284_));
 INV_X1 _10249_ (.A(_08766_),
    .ZN(_01285_));
 AOI21_X4 _10250_ (.A(_01282_),
    .B1(_01284_),
    .B2(_01285_),
    .ZN(_01286_));
 NAND3_X4 _10251_ (.A1(_01208_),
    .A2(_01218_),
    .A3(_01223_),
    .ZN(_01287_));
 NOR4_X4 _10252_ (.A1(_01280_),
    .A2(_01281_),
    .A3(_01286_),
    .A4(_01287_),
    .ZN(_01288_));
 XOR2_X2 _10253_ (.A(_01213_),
    .B(_01226_),
    .Z(_01289_));
 OR2_X1 _10254_ (.A1(_01219_),
    .A2(_01221_),
    .ZN(_01290_));
 AOI21_X4 _10255_ (.A(_01290_),
    .B1(_01204_),
    .B2(net383),
    .ZN(_01291_));
 NOR2_X4 _10256_ (.A1(_01215_),
    .A2(_01217_),
    .ZN(_01292_));
 OAI21_X2 _10257_ (.A(_01289_),
    .B1(_01291_),
    .B2(_01292_),
    .ZN(_01293_));
 AOI21_X4 _10258_ (.A(_01286_),
    .B1(_01293_),
    .B2(_01229_),
    .ZN(_01294_));
 NAND2_X1 _10259_ (.A1(_01086_),
    .A2(_01252_),
    .ZN(_01295_));
 OAI33_X1 _10260_ (.A1(_01278_),
    .A2(_01252_),
    .A3(_01279_),
    .B1(_01288_),
    .B2(_01294_),
    .B3(_01295_),
    .ZN(_01296_));
 OR3_X4 _10261_ (.A1(_01243_),
    .A2(_01085_),
    .A3(_01245_),
    .ZN(_01297_));
 OAI21_X2 _10262_ (.A(_01171_),
    .B1(_01174_),
    .B2(_01148_),
    .ZN(_01298_));
 OR3_X4 _10263_ (.A1(_01233_),
    .A2(_01250_),
    .A3(_08740_),
    .ZN(_01299_));
 OAI21_X4 _10264_ (.A(_01297_),
    .B1(_01298_),
    .B2(_01299_),
    .ZN(_01300_));
 XNOR2_X1 _10265_ (.A(_08780_),
    .B(_01277_),
    .ZN(_01301_));
 XNOR2_X1 _10266_ (.A(_01098_),
    .B(_01301_),
    .ZN(_01302_));
 NAND2_X1 _10267_ (.A1(_01300_),
    .A2(_01302_),
    .ZN(_01303_));
 NAND4_X2 _10268_ (.A1(_01098_),
    .A2(_01252_),
    .A3(_01229_),
    .A4(_01293_),
    .ZN(_01304_));
 NOR3_X4 _10269_ (.A1(_01287_),
    .A2(_01281_),
    .A3(_01280_),
    .ZN(_01305_));
 OAI21_X4 _10270_ (.A(_01303_),
    .B1(_01304_),
    .B2(_01305_),
    .ZN(_01306_));
 AOI21_X4 _10271_ (.A(_01296_),
    .B1(_01272_),
    .B2(_01306_),
    .ZN(_01307_));
 NAND2_X4 _10272_ (.A1(_01275_),
    .A2(_01307_),
    .ZN(_01308_));
 BUF_X8 _10273_ (.A(_01308_),
    .Z(_01309_));
 NOR2_X2 _10274_ (.A1(_01151_),
    .A2(net36),
    .ZN(_01310_));
 INV_X2 _10275_ (.A(_01095_),
    .ZN(_01311_));
 BUF_X2 _10276_ (.A(_08822_),
    .Z(_01312_));
 INV_X1 _10277_ (.A(_08824_),
    .ZN(_01313_));
 BUF_X2 _10278_ (.A(_08827_),
    .Z(_01314_));
 BUF_X2 clone9 (.A(_01720_),
    .Z(net9));
 AOI21_X2 _10280_ (.A(_01314_),
    .B1(_08828_),
    .B2(_08830_),
    .ZN(_01316_));
 INV_X1 _10281_ (.A(_08825_),
    .ZN(_01317_));
 OAI21_X1 _10282_ (.A(_01313_),
    .B1(_01316_),
    .B2(_01317_),
    .ZN(_01318_));
 AOI21_X2 _10283_ (.A(_08821_),
    .B1(_01318_),
    .B2(_01312_),
    .ZN(_01319_));
 CLKBUF_X2 _10284_ (.A(_08831_),
    .Z(_01320_));
 NAND4_X2 _10285_ (.A1(_01312_),
    .A2(_08825_),
    .A3(_08828_),
    .A4(_01320_),
    .ZN(_01321_));
 INV_X1 _10286_ (.A(_08836_),
    .ZN(_01322_));
 OAI21_X2 _10287_ (.A(_08837_),
    .B1(_08839_),
    .B2(_08838_),
    .ZN(_01323_));
 NAND2_X2 _10288_ (.A1(_01322_),
    .A2(_01323_),
    .ZN(_01324_));
 AOI21_X4 _10289_ (.A(_08833_),
    .B1(_01324_),
    .B2(_08834_),
    .ZN(_01325_));
 OR2_X4 _10290_ (.A1(_01325_),
    .A2(_01094_),
    .ZN(_01326_));
 OAI21_X4 _10291_ (.A(_01319_),
    .B1(_01321_),
    .B2(_01326_),
    .ZN(_01327_));
 INV_X1 _10292_ (.A(_01327_),
    .ZN(_01328_));
 BUF_X8 _10293_ (.A(_01300_),
    .Z(_01329_));
 INV_X1 _10294_ (.A(_01301_),
    .ZN(_01330_));
 OAI21_X1 _10295_ (.A(net25),
    .B1(_01330_),
    .B2(_01085_),
    .ZN(_01331_));
 AOI21_X1 _10296_ (.A(_08799_),
    .B1(_08802_),
    .B2(_01270_),
    .ZN(_01332_));
 NAND2_X1 _10297_ (.A1(_01270_),
    .A2(_08803_),
    .ZN(_01333_));
 OAI21_X1 _10298_ (.A(_01332_),
    .B1(_01333_),
    .B2(_01267_),
    .ZN(_01334_));
 XNOR2_X1 _10299_ (.A(net31),
    .B(_01334_),
    .ZN(_01335_));
 NAND2_X1 _10300_ (.A1(_01086_),
    .A2(_01335_),
    .ZN(_01336_));
 NAND2_X2 _10301_ (.A1(_01331_),
    .A2(_01336_),
    .ZN(_01337_));
 AOI21_X4 _10302_ (.A(net25),
    .B1(_01225_),
    .B2(_01231_),
    .ZN(_01338_));
 OAI21_X2 _10303_ (.A(_01328_),
    .B1(_01337_),
    .B2(_01338_),
    .ZN(_01339_));
 OAI21_X4 _10304_ (.A(_09325_),
    .B1(_01248_),
    .B2(_01325_),
    .ZN(_01340_));
 INV_X4 _10305_ (.A(_01340_),
    .ZN(_01341_));
 OAI21_X4 _10306_ (.A(_01319_),
    .B1(_01341_),
    .B2(_01321_),
    .ZN(_01342_));
 INV_X1 _10307_ (.A(_01342_),
    .ZN(_01343_));
 OAI21_X4 _10308_ (.A(_01343_),
    .B1(_01337_),
    .B2(_01338_),
    .ZN(_01344_));
 NAND2_X1 _10309_ (.A1(_01264_),
    .A2(_01265_),
    .ZN(_01345_));
 OR3_X1 _10310_ (.A1(_08814_),
    .A2(_08817_),
    .A3(_01203_),
    .ZN(_01346_));
 OAI21_X2 _10311_ (.A(_01345_),
    .B1(_01346_),
    .B2(_01108_),
    .ZN(_01347_));
 XNOR2_X2 _10312_ (.A(_08812_),
    .B(_01347_),
    .ZN(_01348_));
 NAND2_X1 _10313_ (.A1(_01296_),
    .A2(_01348_),
    .ZN(_01349_));
 AND2_X1 _10314_ (.A1(_01272_),
    .A2(_01348_),
    .ZN(_01350_));
 AND4_X1 _10315_ (.A1(_01252_),
    .A2(_01272_),
    .A3(_01273_),
    .A4(_01348_),
    .ZN(_01351_));
 AOI22_X4 _10316_ (.A1(_01306_),
    .A2(_01350_),
    .B1(_01351_),
    .B2(_01232_),
    .ZN(_01352_));
 NAND2_X2 _10317_ (.A1(_01225_),
    .A2(_01231_),
    .ZN(_01353_));
 INV_X1 _10318_ (.A(_01272_),
    .ZN(_01354_));
 NAND3_X1 _10319_ (.A1(_01168_),
    .A2(_01180_),
    .A3(_01224_),
    .ZN(_01355_));
 NOR4_X2 _10320_ (.A1(_01153_),
    .A2(_01300_),
    .A3(_01230_),
    .A4(_01228_),
    .ZN(_01356_));
 AOI22_X2 _10321_ (.A1(_01355_),
    .A2(_01356_),
    .B1(_01302_),
    .B2(net25),
    .ZN(_01357_));
 OAI222_X2 _10322_ (.A1(_01252_),
    .A2(_01330_),
    .B1(_01353_),
    .B2(_01295_),
    .C1(_01354_),
    .C2(_01357_),
    .ZN(_01358_));
 INV_X1 _10323_ (.A(_01189_),
    .ZN(_01359_));
 NOR2_X1 _10324_ (.A1(_01148_),
    .A2(_01202_),
    .ZN(_08761_));
 MUX2_X1 _10325_ (.A(_01359_),
    .B(_08761_),
    .S(_01229_),
    .Z(_08793_));
 OAI21_X1 _10326_ (.A(_01236_),
    .B1(_08796_),
    .B2(_01237_),
    .ZN(_01360_));
 OR3_X1 _10327_ (.A1(_01237_),
    .A2(_01236_),
    .A3(_08796_),
    .ZN(_01361_));
 AND2_X1 _10328_ (.A1(_01360_),
    .A2(_01361_),
    .ZN(_01362_));
 MUX2_X2 _10329_ (.A(_08793_),
    .B(_01362_),
    .S(_01300_),
    .Z(_08810_));
 NOR3_X4 _10330_ (.A1(net31),
    .A2(_01288_),
    .A3(_01294_),
    .ZN(_01363_));
 NAND3_X2 _10331_ (.A1(_01252_),
    .A2(_01272_),
    .A3(_01273_),
    .ZN(_01364_));
 OAI21_X2 _10332_ (.A(_08810_),
    .B1(_01363_),
    .B2(_01364_),
    .ZN(_01365_));
 OAI211_X4 _10333_ (.A(_01349_),
    .B(_01352_),
    .C1(_01358_),
    .C2(_01365_),
    .ZN(_01366_));
 MUX2_X2 _10334_ (.A(_01339_),
    .B(_01344_),
    .S(_01366_),
    .Z(_01367_));
 BUF_X8 _10335_ (.A(_01367_),
    .Z(_01368_));
 OAI21_X2 _10336_ (.A(_01311_),
    .B1(_01179_),
    .B2(_01368_),
    .ZN(_01369_));
 BUF_X2 _10337_ (.A(_08871_),
    .Z(_01370_));
 NAND4_X1 _10338_ (.A1(_08877_),
    .A2(_08863_),
    .A3(_08874_),
    .A4(_08880_),
    .ZN(_01371_));
 NOR2_X2 _10339_ (.A1(_01170_),
    .A2(_01371_),
    .ZN(_01372_));
 NAND4_X4 _10340_ (.A1(_08868_),
    .A2(_08866_),
    .A3(_01370_),
    .A4(_01372_),
    .ZN(_01373_));
 INV_X4 _10341_ (.A(_01373_),
    .ZN(_01374_));
 AND3_X1 _10342_ (.A1(_01118_),
    .A2(_01369_),
    .A3(_01374_),
    .ZN(_01375_));
 NAND2_X1 _10343_ (.A1(_01312_),
    .A2(_01313_),
    .ZN(_01376_));
 OR2_X1 _10344_ (.A1(_01314_),
    .A2(_01376_),
    .ZN(_01377_));
 INV_X1 _10345_ (.A(_08830_),
    .ZN(_01378_));
 INV_X1 _10346_ (.A(_08833_),
    .ZN(_01379_));
 INV_X1 _10347_ (.A(_08838_),
    .ZN(_01380_));
 OAI21_X1 _10348_ (.A(_08839_),
    .B1(_01110_),
    .B2(_01179_),
    .ZN(_01381_));
 NAND2_X1 _10349_ (.A1(_01380_),
    .A2(_01381_),
    .ZN(_01382_));
 AOI21_X1 _10350_ (.A(_08836_),
    .B1(_01382_),
    .B2(_08837_),
    .ZN(_01383_));
 INV_X1 _10351_ (.A(_08834_),
    .ZN(_01384_));
 OAI21_X1 _10352_ (.A(_01379_),
    .B1(_01383_),
    .B2(_01384_),
    .ZN(_01385_));
 NAND2_X1 _10353_ (.A1(_01320_),
    .A2(_01385_),
    .ZN(_01386_));
 OR2_X1 _10354_ (.A1(_01248_),
    .A2(_08810_),
    .ZN(_01387_));
 NAND2_X1 _10355_ (.A1(_01248_),
    .A2(_08810_),
    .ZN(_01388_));
 AOI221_X2 _10356_ (.A(_08830_),
    .B1(_01232_),
    .B2(_01274_),
    .C1(_01387_),
    .C2(_01388_),
    .ZN(_01389_));
 AOI22_X4 _10357_ (.A1(_01378_),
    .A2(_01386_),
    .B1(_01389_),
    .B2(_01307_),
    .ZN(_01390_));
 XNOR2_X1 _10358_ (.A(_01094_),
    .B(_01348_),
    .ZN(_01391_));
 NOR2_X2 _10359_ (.A1(_08830_),
    .A2(_01391_),
    .ZN(_01392_));
 NOR2_X4 _10360_ (.A1(_01363_),
    .A2(_01364_),
    .ZN(_01393_));
 OAI21_X4 _10361_ (.A(_01392_),
    .B1(_01358_),
    .B2(_01393_),
    .ZN(_01394_));
 INV_X1 _10362_ (.A(_01320_),
    .ZN(_01395_));
 NOR2_X2 _10363_ (.A1(_09325_),
    .A2(_01395_),
    .ZN(_01396_));
 AOI221_X2 _10364_ (.A(_01377_),
    .B1(_01390_),
    .B2(_01394_),
    .C1(_01366_),
    .C2(_01396_),
    .ZN(_01397_));
 INV_X1 _10365_ (.A(_01312_),
    .ZN(_01398_));
 NAND2_X1 _10366_ (.A1(_01398_),
    .A2(_08824_),
    .ZN(_01399_));
 OAI21_X1 _10367_ (.A(_08825_),
    .B1(_08828_),
    .B2(_01314_),
    .ZN(_01400_));
 NAND3_X1 _10368_ (.A1(_01312_),
    .A2(_01313_),
    .A3(_01400_),
    .ZN(_01401_));
 NAND2_X1 _10369_ (.A1(_01399_),
    .A2(_01401_),
    .ZN(_01402_));
 OAI21_X4 _10370_ (.A(_01367_),
    .B1(_01397_),
    .B2(_01402_),
    .ZN(_01403_));
 NOR2_X4 _10371_ (.A1(_01338_),
    .A2(_01337_),
    .ZN(_01404_));
 NOR2_X2 _10372_ (.A1(_01327_),
    .A2(_01404_),
    .ZN(_01405_));
 NOR2_X2 _10373_ (.A1(_01342_),
    .A2(_01404_),
    .ZN(_01406_));
 MUX2_X2 _10374_ (.A(_01405_),
    .B(_01406_),
    .S(_01366_),
    .Z(_01407_));
 AOI221_X2 _10375_ (.A(_01314_),
    .B1(_01394_),
    .B2(_01390_),
    .C1(_01396_),
    .C2(_01366_),
    .ZN(_01408_));
 OR2_X1 _10376_ (.A1(_01312_),
    .A2(_01400_),
    .ZN(_01409_));
 OR3_X4 _10377_ (.A1(_01407_),
    .A2(_01408_),
    .A3(_01409_),
    .ZN(_01410_));
 BUF_X4 _10378_ (.A(_01407_),
    .Z(_01411_));
 INV_X1 _10379_ (.A(_08785_),
    .ZN(_01412_));
 NAND2_X1 _10380_ (.A1(_01238_),
    .A2(_01235_),
    .ZN(_01413_));
 AOI21_X1 _10381_ (.A(_08788_),
    .B1(_01413_),
    .B2(_08789_),
    .ZN(_01414_));
 INV_X1 _10382_ (.A(_08786_),
    .ZN(_01415_));
 OAI21_X1 _10383_ (.A(_01412_),
    .B1(_01414_),
    .B2(_01415_),
    .ZN(_01416_));
 XNOR2_X1 _10384_ (.A(_01240_),
    .B(_01416_),
    .ZN(_01417_));
 NAND2_X1 _10385_ (.A1(net25),
    .A2(_01417_),
    .ZN(_01418_));
 NOR2_X4 _10386_ (.A1(_01292_),
    .A2(_01291_),
    .ZN(_01419_));
 INV_X2 _10387_ (.A(_01419_),
    .ZN(_01420_));
 INV_X1 _10388_ (.A(_08738_),
    .ZN(_01421_));
 NAND2_X1 _10389_ (.A1(_08739_),
    .A2(_01155_),
    .ZN(_01422_));
 NAND2_X1 _10390_ (.A1(_01421_),
    .A2(_01422_),
    .ZN(_01423_));
 XOR2_X1 _10391_ (.A(_08736_),
    .B(_01423_),
    .Z(_01424_));
 NOR2_X1 _10392_ (.A1(_01159_),
    .A2(_01424_),
    .ZN(_01425_));
 OR3_X1 _10393_ (.A1(_08727_),
    .A2(_08729_),
    .A3(_08728_),
    .ZN(_01426_));
 NAND2_X1 _10394_ (.A1(_01161_),
    .A2(_01426_),
    .ZN(_01427_));
 NAND2_X2 _10395_ (.A1(_01164_),
    .A2(_01175_),
    .ZN(_01428_));
 MUX2_X2 _10396_ (.A(_01114_),
    .B(_01427_),
    .S(_01428_),
    .Z(_01429_));
 AOI211_X2 _10397_ (.A(_01420_),
    .B(_01425_),
    .C1(_01429_),
    .C2(net3),
    .ZN(_01430_));
 XOR2_X1 _10398_ (.A(_08749_),
    .B(_01212_),
    .Z(_01431_));
 OAI21_X1 _10399_ (.A(_01431_),
    .B1(_01291_),
    .B2(_01292_),
    .ZN(_01432_));
 NAND2_X1 _10400_ (.A1(_01229_),
    .A2(_01432_),
    .ZN(_01433_));
 NOR2_X1 _10401_ (.A1(_08772_),
    .A2(_01195_),
    .ZN(_01434_));
 XNOR2_X2 _10402_ (.A(_01184_),
    .B(_01434_),
    .ZN(_01435_));
 OAI22_X4 _10403_ (.A1(_01430_),
    .A2(_01433_),
    .B1(_01435_),
    .B2(_01229_),
    .ZN(_01436_));
 OAI21_X2 _10404_ (.A(_01418_),
    .B1(_01436_),
    .B2(net25),
    .ZN(_08798_));
 XNOR2_X1 _10405_ (.A(_01270_),
    .B(_01269_),
    .ZN(_01437_));
 MUX2_X2 _10406_ (.A(_08798_),
    .B(_01437_),
    .S(_01308_),
    .Z(_08820_));
 NAND2_X2 _10407_ (.A1(_01411_),
    .A2(_08820_),
    .ZN(_01438_));
 AND3_X1 _10408_ (.A1(_01403_),
    .A2(_01410_),
    .A3(_01438_),
    .ZN(_01439_));
 BUF_X4 _10409_ (.A(_01439_),
    .Z(_01440_));
 INV_X1 _10410_ (.A(_08841_),
    .ZN(_01441_));
 INV_X1 _10411_ (.A(_08845_),
    .ZN(_01442_));
 INV_X1 _10412_ (.A(_08859_),
    .ZN(_01443_));
 INV_X1 _10413_ (.A(_08853_),
    .ZN(_01444_));
 OAI21_X2 _10414_ (.A(_08854_),
    .B1(_08857_),
    .B2(_08856_),
    .ZN(_01445_));
 NAND2_X2 _10415_ (.A1(_01444_),
    .A2(_01445_),
    .ZN(_01446_));
 AND2_X4 _10416_ (.A1(_08848_),
    .A2(_01446_),
    .ZN(_01447_));
 OAI21_X4 _10417_ (.A(_08860_),
    .B1(_08847_),
    .B2(_01447_),
    .ZN(_01448_));
 AOI21_X4 _10418_ (.A(_01442_),
    .B1(_01443_),
    .B2(_01448_),
    .ZN(_01449_));
 OAI21_X4 _10419_ (.A(_08842_),
    .B1(_08844_),
    .B2(_01449_),
    .ZN(_01450_));
 NAND2_X2 _10420_ (.A1(_01441_),
    .A2(_01450_),
    .ZN(_01451_));
 XNOR2_X2 _10421_ (.A(_08851_),
    .B(_01451_),
    .ZN(_01452_));
 NOR2_X1 _10422_ (.A1(_01440_),
    .A2(_01452_),
    .ZN(_01453_));
 INV_X1 _10423_ (.A(_08851_),
    .ZN(_01454_));
 AOI21_X4 _10424_ (.A(_01454_),
    .B1(_01441_),
    .B2(_01450_),
    .ZN(_01455_));
 OR2_X4 _10425_ (.A1(_01455_),
    .A2(_08850_),
    .ZN(_01456_));
 NAND2_X4 _10426_ (.A1(_01086_),
    .A2(_01456_),
    .ZN(_01457_));
 NAND2_X1 _10427_ (.A1(_01272_),
    .A2(_01348_),
    .ZN(_01458_));
 NAND4_X1 _10428_ (.A1(_01252_),
    .A2(_01272_),
    .A3(_01273_),
    .A4(_01348_),
    .ZN(_01459_));
 OAI22_X1 _10429_ (.A1(_01357_),
    .A2(_01458_),
    .B1(_01459_),
    .B2(_01363_),
    .ZN(_01460_));
 INV_X1 _10430_ (.A(_08810_),
    .ZN(_01461_));
 AOI21_X1 _10431_ (.A(_01461_),
    .B1(_01232_),
    .B2(_01274_),
    .ZN(_01462_));
 AOI221_X4 _10432_ (.A(_01460_),
    .B1(_01462_),
    .B2(_01307_),
    .C1(_01296_),
    .C2(_01348_),
    .ZN(_01463_));
 XNOR2_X2 _10433_ (.A(_01261_),
    .B(_01267_),
    .ZN(_01464_));
 AND2_X1 _10434_ (.A1(_01331_),
    .A2(_01336_),
    .ZN(_01465_));
 OAI21_X1 _10435_ (.A(_01252_),
    .B1(_01288_),
    .B2(_01294_),
    .ZN(_01466_));
 AOI211_X2 _10436_ (.A(_01327_),
    .B(_01464_),
    .C1(_01465_),
    .C2(_01466_),
    .ZN(_01467_));
 OAI21_X2 _10437_ (.A(_01467_),
    .B1(_01358_),
    .B2(_01393_),
    .ZN(_01468_));
 XNOR2_X1 _10438_ (.A(_01415_),
    .B(_01414_),
    .ZN(_01469_));
 NAND2_X1 _10439_ (.A1(_01329_),
    .A2(_01469_),
    .ZN(_01470_));
 OR2_X1 _10440_ (.A1(_08757_),
    .A2(_08756_),
    .ZN(_01471_));
 AOI21_X1 _10441_ (.A(_08754_),
    .B1(_01471_),
    .B2(_08755_),
    .ZN(_01472_));
 XNOR2_X1 _10442_ (.A(_08752_),
    .B(_01472_),
    .ZN(_01473_));
 XOR2_X1 _10443_ (.A(_08739_),
    .B(_01155_),
    .Z(_01474_));
 NOR2_X1 _10444_ (.A1(_08729_),
    .A2(_01164_),
    .ZN(_08737_));
 MUX2_X1 _10445_ (.A(_01474_),
    .B(_08737_),
    .S(_01159_),
    .Z(_08750_));
 MUX2_X1 _10446_ (.A(_01473_),
    .B(_08750_),
    .S(_01419_),
    .Z(_08771_));
 XNOR2_X1 _10447_ (.A(_08773_),
    .B(_01192_),
    .ZN(_01475_));
 MUX2_X2 _10448_ (.A(_08771_),
    .B(_01475_),
    .S(_01230_),
    .Z(_08784_));
 OAI21_X4 _10449_ (.A(_01470_),
    .B1(_08784_),
    .B2(_01329_),
    .ZN(_01476_));
 OR4_X2 _10450_ (.A1(_01393_),
    .A2(_01358_),
    .A3(_01339_),
    .A4(_01476_),
    .ZN(_01477_));
 NAND2_X1 _10451_ (.A1(_08828_),
    .A2(_01320_),
    .ZN(_01478_));
 OAI21_X1 _10452_ (.A(_01316_),
    .B1(_01478_),
    .B2(_01326_),
    .ZN(_01479_));
 XNOR2_X1 _10453_ (.A(_01317_),
    .B(_01479_),
    .ZN(_01480_));
 NAND2_X2 _10454_ (.A1(_01339_),
    .A2(_01480_),
    .ZN(_01481_));
 NAND4_X4 _10455_ (.A1(_01463_),
    .A2(_01468_),
    .A3(_01477_),
    .A4(_01481_),
    .ZN(_01482_));
 AOI211_X2 _10456_ (.A(_01344_),
    .B(_01464_),
    .C1(_01275_),
    .C2(_01307_),
    .ZN(_01483_));
 NOR4_X4 _10457_ (.A1(_01393_),
    .A2(_01358_),
    .A3(_01344_),
    .A4(_01476_),
    .ZN(_01484_));
 OAI21_X1 _10458_ (.A(_01316_),
    .B1(_01478_),
    .B2(_01341_),
    .ZN(_01485_));
 XNOR2_X1 _10459_ (.A(_01317_),
    .B(_01485_),
    .ZN(_01486_));
 AND2_X1 _10460_ (.A1(_01344_),
    .A2(_01486_),
    .ZN(_01487_));
 OR4_X1 _10461_ (.A1(_01463_),
    .A2(_01483_),
    .A3(_01484_),
    .A4(_01487_),
    .ZN(_01488_));
 BUF_X4 _10462_ (.A(_01488_),
    .Z(_01489_));
 AOI21_X4 _10463_ (.A(_01457_),
    .B1(_01482_),
    .B2(_01489_),
    .ZN(_01490_));
 NAND2_X4 _10464_ (.A1(_01456_),
    .A2(_01085_),
    .ZN(_01491_));
 NAND2_X4 _10465_ (.A1(_01491_),
    .A2(_01115_),
    .ZN(_01492_));
 AND3_X4 _10466_ (.A1(_01492_),
    .A2(_01482_),
    .A3(_01489_),
    .ZN(_01493_));
 NOR2_X4 _10467_ (.A1(_01493_),
    .A2(_01490_),
    .ZN(_01494_));
 NAND2_X1 _10468_ (.A1(_08740_),
    .A2(_01159_),
    .ZN(_01495_));
 OAI21_X1 _10469_ (.A(_01495_),
    .B1(net3),
    .B2(_08742_),
    .ZN(_08753_));
 XNOR2_X1 _10470_ (.A(_08755_),
    .B(_01211_),
    .ZN(_01496_));
 MUX2_X1 _10471_ (.A(_08753_),
    .B(_01496_),
    .S(_01420_),
    .Z(_08774_));
 OR2_X1 _10472_ (.A1(_01189_),
    .A2(_08762_),
    .ZN(_01497_));
 AOI21_X1 _10473_ (.A(_08759_),
    .B1(_01497_),
    .B2(_01187_),
    .ZN(_01498_));
 XNOR2_X1 _10474_ (.A(_08776_),
    .B(_01498_),
    .ZN(_01499_));
 MUX2_X1 _10475_ (.A(_08774_),
    .B(_01499_),
    .S(_01230_),
    .Z(_08787_));
 XOR2_X1 _10476_ (.A(_08789_),
    .B(_01413_),
    .Z(_01500_));
 MUX2_X1 _10477_ (.A(_08787_),
    .B(_01500_),
    .S(_01329_),
    .Z(_08804_));
 INV_X1 _10478_ (.A(_08811_),
    .ZN(_01501_));
 OAI21_X1 _10479_ (.A(_01501_),
    .B1(_01347_),
    .B2(_01263_),
    .ZN(_01502_));
 AOI21_X1 _10480_ (.A(_08808_),
    .B1(_01502_),
    .B2(_08809_),
    .ZN(_01503_));
 XNOR2_X1 _10481_ (.A(_08806_),
    .B(_01503_),
    .ZN(_01504_));
 MUX2_X2 _10482_ (.A(_08804_),
    .B(_01504_),
    .S(_01308_),
    .Z(_08826_));
 NOR2_X1 _10483_ (.A1(_01368_),
    .A2(_08826_),
    .ZN(_01505_));
 AOI22_X4 _10484_ (.A1(_01394_),
    .A2(_01390_),
    .B1(_01396_),
    .B2(_01366_),
    .ZN(_01506_));
 XOR2_X2 _10485_ (.A(_08828_),
    .B(_01506_),
    .Z(_01507_));
 AOI21_X4 _10486_ (.A(_01505_),
    .B1(_01507_),
    .B2(_01368_),
    .ZN(_08849_));
 AND3_X1 _10487_ (.A1(_01440_),
    .A2(_01494_),
    .A3(_08849_),
    .ZN(_01508_));
 OAI21_X2 _10488_ (.A(_01375_),
    .B1(_01453_),
    .B2(_01508_),
    .ZN(_01509_));
 MUX2_X2 _10489_ (.A(_01327_),
    .B(_01342_),
    .S(_01366_),
    .Z(_01510_));
 AND2_X1 _10490_ (.A1(_01404_),
    .A2(_01510_),
    .ZN(_01511_));
 NOR2_X4 _10491_ (.A1(_08850_),
    .A2(_01455_),
    .ZN(_01512_));
 NOR2_X2 _10492_ (.A1(_01118_),
    .A2(_01512_),
    .ZN(_01513_));
 AND4_X4 _10493_ (.A1(_01463_),
    .A2(_01468_),
    .A3(_01477_),
    .A4(_01481_),
    .ZN(_01514_));
 NOR4_X4 _10494_ (.A1(_01463_),
    .A2(_01483_),
    .A3(_01484_),
    .A4(_01487_),
    .ZN(_01515_));
 OAI21_X4 _10495_ (.A(_01513_),
    .B1(_01514_),
    .B2(_01515_),
    .ZN(_01516_));
 NAND3_X4 _10496_ (.A1(_01489_),
    .A2(_01482_),
    .A3(_01492_),
    .ZN(_01517_));
 NAND2_X4 _10497_ (.A1(_01516_),
    .A2(_01517_),
    .ZN(_01518_));
 NAND2_X4 _10498_ (.A1(net383),
    .A2(_01177_),
    .ZN(_01519_));
 NAND3_X1 _10499_ (.A1(_01086_),
    .A2(_01519_),
    .A3(_01374_),
    .ZN(_01520_));
 NAND2_X1 _10500_ (.A1(_01095_),
    .A2(_01086_),
    .ZN(_01521_));
 OAI22_X2 _10501_ (.A1(_01367_),
    .A2(_01520_),
    .B1(_01521_),
    .B2(_01373_),
    .ZN(_01522_));
 OAI21_X2 _10502_ (.A(_01149_),
    .B1(_01179_),
    .B2(_01308_),
    .ZN(_01523_));
 NAND4_X1 _10503_ (.A1(_08842_),
    .A2(_08854_),
    .A3(_08860_),
    .A4(_08851_),
    .ZN(_01524_));
 NAND3_X1 _10504_ (.A1(_08857_),
    .A2(_08845_),
    .A3(_08848_),
    .ZN(_01525_));
 NOR3_X1 _10505_ (.A1(_01097_),
    .A2(_01524_),
    .A3(_01525_),
    .ZN(_01526_));
 NAND2_X1 _10506_ (.A1(_01523_),
    .A2(_01526_),
    .ZN(_01527_));
 NOR2_X4 _10507_ (.A1(_01515_),
    .A2(_01514_),
    .ZN(_01528_));
 OAI221_X2 _10508_ (.A(_01522_),
    .B1(_01507_),
    .B2(net11),
    .C1(_01527_),
    .C2(_01528_),
    .ZN(_01529_));
 NOR3_X2 _10509_ (.A1(_01368_),
    .A2(_08820_),
    .A3(_08826_),
    .ZN(_01530_));
 NAND3_X1 _10510_ (.A1(_01398_),
    .A2(_08825_),
    .A3(_01314_),
    .ZN(_01531_));
 NAND3_X1 _10511_ (.A1(_01399_),
    .A2(_01401_),
    .A3(_01531_),
    .ZN(_01532_));
 NOR2_X1 _10512_ (.A1(net11),
    .A2(_01532_),
    .ZN(_01533_));
 MUX2_X1 _10513_ (.A(_01409_),
    .B(_01377_),
    .S(_01506_),
    .Z(_01534_));
 AOI21_X1 _10514_ (.A(_01530_),
    .B1(_01533_),
    .B2(_01534_),
    .ZN(_01535_));
 NOR3_X2 _10515_ (.A1(_01518_),
    .A2(_01529_),
    .A3(_01535_),
    .ZN(_01536_));
 OAI211_X2 _10516_ (.A(_01369_),
    .B(_01374_),
    .C1(_01490_),
    .C2(_01493_),
    .ZN(_01537_));
 XNOR2_X2 _10517_ (.A(_01454_),
    .B(_01451_),
    .ZN(_01538_));
 XNOR2_X2 _10518_ (.A(_01118_),
    .B(_01538_),
    .ZN(_01539_));
 INV_X1 _10519_ (.A(_01539_),
    .ZN(_01540_));
 OAI21_X1 _10520_ (.A(_01440_),
    .B1(_01537_),
    .B2(_01540_),
    .ZN(_01541_));
 AND2_X1 _10521_ (.A1(_01452_),
    .A2(_01522_),
    .ZN(_01542_));
 OR2_X1 _10522_ (.A1(_01518_),
    .A2(_01542_),
    .ZN(_01543_));
 AOI211_X4 _10523_ (.A(_01511_),
    .B(_01536_),
    .C1(_01541_),
    .C2(_01543_),
    .ZN(_01544_));
 NAND2_X1 _10524_ (.A1(_01118_),
    .A2(_01512_),
    .ZN(_01545_));
 AOI22_X2 _10525_ (.A1(_01489_),
    .A2(_01482_),
    .B1(_01457_),
    .B2(_01545_),
    .ZN(_01546_));
 NOR2_X2 _10526_ (.A1(_01115_),
    .A2(_01118_),
    .ZN(_01547_));
 NAND2_X1 _10527_ (.A1(_01547_),
    .A2(_01512_),
    .ZN(_01548_));
 AOI211_X2 _10528_ (.A(_01515_),
    .B(_01514_),
    .C1(_01491_),
    .C2(_01548_),
    .ZN(_01549_));
 NOR2_X1 _10529_ (.A1(_01118_),
    .A2(_01456_),
    .ZN(_01550_));
 AND4_X1 _10530_ (.A1(_01404_),
    .A2(_01489_),
    .A3(_01482_),
    .A4(_01510_),
    .ZN(_01551_));
 AOI211_X2 _10531_ (.A(_01546_),
    .B(_01549_),
    .C1(_01550_),
    .C2(_01551_),
    .ZN(_01552_));
 NAND2_X1 _10532_ (.A1(_01528_),
    .A2(_01550_),
    .ZN(_01553_));
 NAND2_X4 _10533_ (.A1(_01404_),
    .A2(_01510_),
    .ZN(_01554_));
 NAND4_X4 _10534_ (.A1(_01403_),
    .A2(_01410_),
    .A3(_01438_),
    .A4(_01554_),
    .ZN(_01555_));
 OAI221_X2 _10535_ (.A(_01552_),
    .B1(_01553_),
    .B2(_01440_),
    .C1(_01528_),
    .C2(_01555_),
    .ZN(_01556_));
 OR3_X1 _10536_ (.A1(_01367_),
    .A2(_08820_),
    .A3(_08826_),
    .ZN(_01557_));
 OR2_X1 _10537_ (.A1(_01411_),
    .A2(_01532_),
    .ZN(_01558_));
 NAND2_X1 _10538_ (.A1(net43),
    .A2(_01409_),
    .ZN(_01559_));
 NOR2_X1 _10539_ (.A1(_01314_),
    .A2(_01376_),
    .ZN(_01560_));
 OR2_X1 _10540_ (.A1(net43),
    .A2(_01560_),
    .ZN(_01561_));
 MUX2_X1 _10541_ (.A(_01559_),
    .B(_01561_),
    .S(_01506_),
    .Z(_01562_));
 OAI21_X4 _10542_ (.A(_01557_),
    .B1(_01558_),
    .B2(_01562_),
    .ZN(_01563_));
 INV_X1 _10543_ (.A(_08873_),
    .ZN(_01564_));
 INV_X1 _10544_ (.A(_08879_),
    .ZN(_01565_));
 INV_X1 _10545_ (.A(_08865_),
    .ZN(_01566_));
 OAI21_X1 _10546_ (.A(_08866_),
    .B1(_08867_),
    .B2(_08868_),
    .ZN(_01567_));
 NAND2_X1 _10547_ (.A1(_01566_),
    .A2(_01567_),
    .ZN(_01568_));
 AND2_X4 _10548_ (.A1(_01568_),
    .A2(_08863_),
    .ZN(_01569_));
 OAI21_X4 _10549_ (.A(_08880_),
    .B1(_01569_),
    .B2(_08862_),
    .ZN(_01570_));
 NAND2_X4 _10550_ (.A1(_01565_),
    .A2(_01570_),
    .ZN(_01571_));
 AOI21_X4 _10551_ (.A(_08876_),
    .B1(_01571_),
    .B2(_08877_),
    .ZN(_01572_));
 INV_X1 _10552_ (.A(_08874_),
    .ZN(_01573_));
 OAI21_X4 _10553_ (.A(_01564_),
    .B1(_01573_),
    .B2(_01572_),
    .ZN(_01574_));
 AND2_X4 _10554_ (.A1(_01574_),
    .A2(_01370_),
    .ZN(_01575_));
 NOR2_X4 _10555_ (.A1(_08870_),
    .A2(_01575_),
    .ZN(_01576_));
 NOR2_X4 _10556_ (.A1(_01576_),
    .A2(_01118_),
    .ZN(_01577_));
 AND4_X2 _10557_ (.A1(_01494_),
    .A2(_01554_),
    .A3(_01563_),
    .A4(_01577_),
    .ZN(_01578_));
 NAND2_X1 _10558_ (.A1(_01452_),
    .A2(_01577_),
    .ZN(_01579_));
 AND4_X4 _10559_ (.A1(_01403_),
    .A2(_01410_),
    .A3(_01438_),
    .A4(_01554_),
    .ZN(_01580_));
 AOI21_X1 _10560_ (.A(_01579_),
    .B1(_01580_),
    .B2(_01494_),
    .ZN(_01581_));
 NOR3_X2 _10561_ (.A1(_01490_),
    .A2(_01493_),
    .A3(_01511_),
    .ZN(_01582_));
 OR2_X2 _10562_ (.A1(_08870_),
    .A2(_01575_),
    .ZN(_01583_));
 NAND2_X2 _10563_ (.A1(_01118_),
    .A2(_01583_),
    .ZN(_01584_));
 AOI22_X2 _10564_ (.A1(_01582_),
    .A2(_01563_),
    .B1(_01584_),
    .B2(_01115_),
    .ZN(_01585_));
 OAI21_X4 _10565_ (.A(_01452_),
    .B1(_01555_),
    .B2(_01518_),
    .ZN(_01586_));
 AOI211_X2 _10566_ (.A(_01578_),
    .B(_01581_),
    .C1(_01585_),
    .C2(_01586_),
    .ZN(_01587_));
 NAND4_X2 _10567_ (.A1(_01509_),
    .A2(_01544_),
    .A3(_01556_),
    .A4(_01587_),
    .ZN(_01588_));
 BUF_X4 _10568_ (.A(_01588_),
    .Z(_01589_));
 XOR2_X2 _10569_ (.A(_01370_),
    .B(_01574_),
    .Z(_01590_));
 NOR3_X2 _10570_ (.A1(_08894_),
    .A2(_08897_),
    .A3(_08900_),
    .ZN(_01591_));
 OAI21_X2 _10571_ (.A(_08901_),
    .B1(_08882_),
    .B2(_08883_),
    .ZN(_01592_));
 OR2_X1 _10572_ (.A1(_08882_),
    .A2(_08885_),
    .ZN(_01593_));
 INV_X1 _10573_ (.A(_08888_),
    .ZN(_01594_));
 NOR2_X4 _10574_ (.A1(_01108_),
    .A2(_01203_),
    .ZN(_01595_));
 NAND3_X2 _10575_ (.A1(_01595_),
    .A2(_01275_),
    .A3(_01307_),
    .ZN(_01596_));
 BUF_X1 _10576_ (.A(_08892_),
    .Z(_01597_));
 AOI21_X1 _10577_ (.A(_08891_),
    .B1(_01596_),
    .B2(_01597_),
    .ZN(_01598_));
 INV_X1 _10578_ (.A(_08889_),
    .ZN(_01599_));
 OAI21_X2 _10579_ (.A(_01594_),
    .B1(_01598_),
    .B2(_01599_),
    .ZN(_01600_));
 OAI21_X4 clone3 (.A(_01145_),
    .B1(_08732_),
    .B2(_01158_),
    .ZN(net3));
 AOI21_X4 _10581_ (.A(_01593_),
    .B1(_01600_),
    .B2(_08886_),
    .ZN(_01602_));
 OAI21_X4 _10582_ (.A(_01591_),
    .B1(_01602_),
    .B2(_01592_),
    .ZN(_01603_));
 NOR2_X4 clone4 (.A1(_01493_),
    .A2(_01490_),
    .ZN(net4));
 NOR3_X2 _10584_ (.A1(_08898_),
    .A2(_08894_),
    .A3(_08897_),
    .ZN(_01605_));
 NOR2_X2 _10585_ (.A1(_08895_),
    .A2(_08894_),
    .ZN(_01606_));
 NOR2_X4 _10586_ (.A1(_01606_),
    .A2(_01605_),
    .ZN(_01607_));
 NAND2_X2 _10587_ (.A1(_01603_),
    .A2(_01607_),
    .ZN(_01608_));
 NOR3_X4 _10588_ (.A1(_01608_),
    .A2(_01590_),
    .A3(_01119_),
    .ZN(_01609_));
 XNOR2_X1 _10589_ (.A(_01370_),
    .B(_01574_),
    .ZN(_01610_));
 NAND3_X4 _10590_ (.A1(_01603_),
    .A2(_01119_),
    .A3(_01607_),
    .ZN(_01611_));
 AOI21_X4 _10591_ (.A(_01610_),
    .B1(_01611_),
    .B2(_01115_),
    .ZN(_01612_));
 OAI21_X2 _10592_ (.A(net10),
    .B1(_01609_),
    .B2(_01612_),
    .ZN(_01613_));
 NAND3_X1 _10593_ (.A1(_01119_),
    .A2(_01369_),
    .A3(_01374_),
    .ZN(_01614_));
 NAND3_X2 _10594_ (.A1(_01403_),
    .A2(_01410_),
    .A3(_01438_),
    .ZN(_01615_));
 NAND2_X1 _10595_ (.A1(_01615_),
    .A2(_01538_),
    .ZN(_01616_));
 NAND3_X2 _10596_ (.A1(_01440_),
    .A2(_01494_),
    .A3(_08849_),
    .ZN(_01617_));
 AOI21_X4 _10597_ (.A(_01614_),
    .B1(_01616_),
    .B2(_01617_),
    .ZN(_01618_));
 OR3_X1 _10598_ (.A1(_01518_),
    .A2(_01529_),
    .A3(_01535_),
    .ZN(_01619_));
 NAND2_X4 _10599_ (.A1(_01411_),
    .A2(_01519_),
    .ZN(_01620_));
 AOI221_X2 _10600_ (.A(_01373_),
    .B1(_01517_),
    .B2(_01516_),
    .C1(_01311_),
    .C2(_01620_),
    .ZN(_01621_));
 AOI21_X2 _10601_ (.A(_01615_),
    .B1(_01621_),
    .B2(_01539_),
    .ZN(_01622_));
 NOR2_X1 _10602_ (.A1(_01518_),
    .A2(_01542_),
    .ZN(_01623_));
 OAI211_X4 _10603_ (.A(_01554_),
    .B(_01619_),
    .C1(_01622_),
    .C2(_01623_),
    .ZN(_01624_));
 NOR2_X1 _10604_ (.A1(_01086_),
    .A2(_01456_),
    .ZN(_01625_));
 OAI22_X2 _10605_ (.A1(_01515_),
    .A2(_01514_),
    .B1(_01513_),
    .B2(_01625_),
    .ZN(_01626_));
 INV_X1 _10606_ (.A(_01491_),
    .ZN(_01627_));
 AND2_X1 _10607_ (.A1(_01547_),
    .A2(_01512_),
    .ZN(_01628_));
 OAI211_X2 _10608_ (.A(_01489_),
    .B(_01482_),
    .C1(_01627_),
    .C2(_01628_),
    .ZN(_01629_));
 INV_X1 _10609_ (.A(_01550_),
    .ZN(_01630_));
 NAND4_X1 _10610_ (.A1(_01404_),
    .A2(_01489_),
    .A3(_01482_),
    .A4(_01510_),
    .ZN(_01631_));
 OAI211_X2 _10611_ (.A(_01626_),
    .B(_01629_),
    .C1(_01630_),
    .C2(_01631_),
    .ZN(_01632_));
 NAND2_X2 _10612_ (.A1(_01489_),
    .A2(_01482_),
    .ZN(_01633_));
 NOR2_X1 _10613_ (.A1(_01633_),
    .A2(_01630_),
    .ZN(_01634_));
 AOI221_X2 _10614_ (.A(_01632_),
    .B1(_01634_),
    .B2(_01615_),
    .C1(_01633_),
    .C2(_01580_),
    .ZN(_01635_));
 CLKBUF_X3 _10615_ (.A(_01635_),
    .Z(_01636_));
 NAND4_X2 _10616_ (.A1(net4),
    .A2(_01554_),
    .A3(_01563_),
    .A4(_01577_),
    .ZN(_01637_));
 NOR3_X1 _10617_ (.A1(_01119_),
    .A2(_01538_),
    .A3(_01576_),
    .ZN(_01638_));
 OAI21_X2 _10618_ (.A(_01638_),
    .B1(_01555_),
    .B2(_01518_),
    .ZN(_01639_));
 NAND2_X1 _10619_ (.A1(_01115_),
    .A2(_01584_),
    .ZN(_01640_));
 AND2_X1 _10620_ (.A1(net43),
    .A2(_01409_),
    .ZN(_01641_));
 NOR2_X1 _10621_ (.A1(net43),
    .A2(_01560_),
    .ZN(_01642_));
 MUX2_X1 _10622_ (.A(_01641_),
    .B(_01642_),
    .S(_01506_),
    .Z(_01643_));
 AOI21_X2 _10623_ (.A(_01530_),
    .B1(_01533_),
    .B2(_01643_),
    .ZN(_01644_));
 NAND3_X2 _10624_ (.A1(_01516_),
    .A2(_01517_),
    .A3(_01554_),
    .ZN(_01645_));
 OAI21_X2 _10625_ (.A(_01640_),
    .B1(_01644_),
    .B2(_01645_),
    .ZN(_01646_));
 AOI21_X4 _10626_ (.A(_01538_),
    .B1(_01580_),
    .B2(net4),
    .ZN(_01647_));
 OAI211_X4 _10627_ (.A(_01637_),
    .B(_01639_),
    .C1(_01646_),
    .C2(_01647_),
    .ZN(_01648_));
 NOR4_X4 _10628_ (.A1(_01618_),
    .A2(_01624_),
    .A3(_01636_),
    .A4(_01648_),
    .ZN(_01649_));
 XOR2_X1 _10629_ (.A(_01187_),
    .B(_01497_),
    .Z(_01650_));
 NOR3_X2 _10630_ (.A1(_08757_),
    .A2(_01215_),
    .A3(_01217_),
    .ZN(_08758_));
 MUX2_X1 _10631_ (.A(_01650_),
    .B(_08758_),
    .S(_01229_),
    .Z(_08790_));
 NOR2_X1 _10632_ (.A1(_01329_),
    .A2(_08790_),
    .ZN(_01651_));
 INV_X1 _10633_ (.A(_08794_),
    .ZN(_01652_));
 NAND2_X1 _10634_ (.A1(_01652_),
    .A2(_01360_),
    .ZN(_01653_));
 XNOR2_X1 _10635_ (.A(_08792_),
    .B(_01653_),
    .ZN(_01654_));
 AOI21_X2 _10636_ (.A(_01651_),
    .B1(_01654_),
    .B2(_01329_),
    .ZN(_08807_));
 NOR2_X1 _10637_ (.A1(_08811_),
    .A2(_01266_),
    .ZN(_01655_));
 XNOR2_X1 _10638_ (.A(_08809_),
    .B(_01655_),
    .ZN(_01656_));
 MUX2_X1 _10639_ (.A(_08807_),
    .B(_01656_),
    .S(_01308_),
    .Z(_08829_));
 MUX2_X1 _10640_ (.A(_01326_),
    .B(_01341_),
    .S(_01366_),
    .Z(_01657_));
 XNOR2_X1 _10641_ (.A(_01320_),
    .B(_01657_),
    .ZN(_01658_));
 MUX2_X2 _10642_ (.A(_08829_),
    .B(_01658_),
    .S(_01368_),
    .Z(_08840_));
 NAND3_X2 _10643_ (.A1(net4),
    .A2(_01580_),
    .A3(_08840_),
    .ZN(_01659_));
 NAND2_X4 _10644_ (.A1(_01494_),
    .A2(_01580_),
    .ZN(_01660_));
 OR3_X1 _10645_ (.A1(_08842_),
    .A2(_08844_),
    .A3(_01449_),
    .ZN(_01661_));
 AND2_X1 _10646_ (.A1(_01450_),
    .A2(_01661_),
    .ZN(_01662_));
 NAND2_X1 _10647_ (.A1(_01660_),
    .A2(_01662_),
    .ZN(_01663_));
 AOI22_X4 _10648_ (.A1(_01659_),
    .A2(_01663_),
    .B1(_01115_),
    .B2(_01611_),
    .ZN(_01664_));
 MUX2_X2 _10649_ (.A(_08840_),
    .B(_01662_),
    .S(_01660_),
    .Z(_08869_));
 NOR3_X4 _10650_ (.A1(_01608_),
    .A2(_08869_),
    .A3(_01119_),
    .ZN(_01665_));
 OAI21_X4 _10651_ (.A(_01649_),
    .B1(_01664_),
    .B2(_01665_),
    .ZN(_01666_));
 NAND2_X1 _10652_ (.A1(_01118_),
    .A2(_01576_),
    .ZN(_01667_));
 NOR3_X1 _10653_ (.A1(_01528_),
    .A2(_01512_),
    .A3(_01667_),
    .ZN(_01668_));
 NOR2_X1 _10654_ (.A1(_01456_),
    .A2(_01667_),
    .ZN(_01669_));
 AOI22_X2 _10655_ (.A1(_01555_),
    .A2(_01668_),
    .B1(_01669_),
    .B2(_01528_),
    .ZN(_01670_));
 NOR2_X2 _10656_ (.A1(_01645_),
    .A2(_01644_),
    .ZN(_01671_));
 OAI21_X2 _10657_ (.A(_01670_),
    .B1(_01671_),
    .B2(_01647_),
    .ZN(_01672_));
 AOI221_X2 _10658_ (.A(_01672_),
    .B1(_01544_),
    .B2(_01509_),
    .C1(_01087_),
    .C2(_01583_),
    .ZN(_01673_));
 NAND2_X2 _10659_ (.A1(_01582_),
    .A2(_01563_),
    .ZN(_01674_));
 AOI22_X1 _10660_ (.A1(_01586_),
    .A2(_01674_),
    .B1(_01636_),
    .B2(_01670_),
    .ZN(_01675_));
 NAND2_X2 _10661_ (.A1(_01087_),
    .A2(_01576_),
    .ZN(_01676_));
 NAND3_X1 _10662_ (.A1(_01153_),
    .A2(_01633_),
    .A3(_01512_),
    .ZN(_01677_));
 NAND3_X1 _10663_ (.A1(_01115_),
    .A2(_01528_),
    .A3(_01512_),
    .ZN(_01678_));
 AOI21_X1 _10664_ (.A(_01580_),
    .B1(_01677_),
    .B2(_01678_),
    .ZN(_01679_));
 NAND3_X1 _10665_ (.A1(_01115_),
    .A2(_01633_),
    .A3(_01456_),
    .ZN(_01680_));
 NAND2_X1 _10666_ (.A1(_01153_),
    .A2(_01456_),
    .ZN(_01681_));
 OAI21_X1 _10667_ (.A(_01680_),
    .B1(_01681_),
    .B2(_01633_),
    .ZN(_01682_));
 NOR3_X1 _10668_ (.A1(_01153_),
    .A2(_01528_),
    .A3(_01555_),
    .ZN(_01683_));
 NOR4_X2 _10669_ (.A1(_01676_),
    .A2(_01679_),
    .A3(_01682_),
    .A4(_01683_),
    .ZN(_01684_));
 NOR2_X2 _10670_ (.A1(_01647_),
    .A2(_01671_),
    .ZN(_01685_));
 AOI21_X2 _10671_ (.A(_01675_),
    .B1(_01684_),
    .B2(_01685_),
    .ZN(_01686_));
 OR2_X1 _10672_ (.A1(_01584_),
    .A2(_01636_),
    .ZN(_01687_));
 AOI21_X2 _10673_ (.A(_01672_),
    .B1(_01544_),
    .B2(_01509_),
    .ZN(_01688_));
 OAI22_X4 _10674_ (.A1(_01673_),
    .A2(_01686_),
    .B1(_01687_),
    .B2(_01688_),
    .ZN(_01689_));
 NOR3_X1 _10675_ (.A1(_01490_),
    .A2(_01493_),
    .A3(_01554_),
    .ZN(_01690_));
 MUX2_X2 _10676_ (.A(_01518_),
    .B(_01690_),
    .S(_01440_),
    .Z(_01691_));
 AOI21_X4 _10677_ (.A(_01554_),
    .B1(net4),
    .B2(_01440_),
    .ZN(_01692_));
 NAND2_X2 _10678_ (.A1(_01556_),
    .A2(_01587_),
    .ZN(_01693_));
 AOI21_X4 _10679_ (.A(_01691_),
    .B1(_01692_),
    .B2(_01693_),
    .ZN(_01694_));
 AND4_X1 _10680_ (.A1(_01613_),
    .A2(_01666_),
    .A3(_01689_),
    .A4(_01694_),
    .ZN(_01695_));
 BUF_X4 _10681_ (.A(_01695_),
    .Z(_01696_));
 AOI21_X1 _10682_ (.A(_01143_),
    .B1(_01310_),
    .B2(_01696_),
    .ZN(_01697_));
 OAI21_X1 _10683_ (.A(_08980_),
    .B1(_08982_),
    .B2(_01697_),
    .ZN(_01698_));
 INV_X1 _10684_ (.A(_08979_),
    .ZN(_01699_));
 AOI21_X1 _10685_ (.A(_01141_),
    .B1(_01698_),
    .B2(_01699_),
    .ZN(_01700_));
 AOI21_X1 _10686_ (.A(_08973_),
    .B1(_08976_),
    .B2(_01140_),
    .ZN(_01701_));
 INV_X1 _10687_ (.A(_01701_),
    .ZN(_01702_));
 OR2_X1 _10688_ (.A1(_01700_),
    .A2(_01702_),
    .ZN(_01703_));
 AOI21_X1 _10689_ (.A(_08970_),
    .B1(_01703_),
    .B2(_08971_),
    .ZN(_01704_));
 BUF_X1 _10690_ (.A(_08968_),
    .Z(_01705_));
 INV_X1 _10691_ (.A(_01705_),
    .ZN(_01706_));
 OAI21_X1 _10692_ (.A(_01139_),
    .B1(_01704_),
    .B2(_01706_),
    .ZN(_01707_));
 XOR2_X2 _10693_ (.A(_08965_),
    .B(_01707_),
    .Z(_01708_));
 NAND2_X1 _10694_ (.A1(_01137_),
    .A2(_01708_),
    .ZN(_01709_));
 BUF_X4 _10695_ (.A(_01201_),
    .Z(_01710_));
 AOI22_X4 _10696_ (.A1(_01595_),
    .A2(_01309_),
    .B1(_01620_),
    .B2(_01710_),
    .ZN(_01711_));
 INV_X4 _10697_ (.A(_01711_),
    .ZN(_08855_));
 NOR2_X4 _10698_ (.A1(_01660_),
    .A2(_08855_),
    .ZN(_01712_));
 AOI21_X2 _10699_ (.A(_01712_),
    .B1(_01660_),
    .B2(_08857_),
    .ZN(_08864_));
 OR3_X1 _10700_ (.A1(_08868_),
    .A2(_08866_),
    .A3(_08867_),
    .ZN(_01713_));
 AND2_X1 _10701_ (.A1(_01567_),
    .A2(_01713_),
    .ZN(_01714_));
 MUX2_X1 _10702_ (.A(_08864_),
    .B(_01714_),
    .S(_01589_),
    .Z(_08884_));
 INV_X1 _10703_ (.A(_08891_),
    .ZN(_01715_));
 INV_X1 _10704_ (.A(_01597_),
    .ZN(_01716_));
 OAI21_X1 _10705_ (.A(_01715_),
    .B1(_01310_),
    .B2(_01716_),
    .ZN(_01717_));
 AOI21_X1 _10706_ (.A(_08888_),
    .B1(_01717_),
    .B2(_08889_),
    .ZN(_01718_));
 XNOR2_X1 _10707_ (.A(_08886_),
    .B(_01718_),
    .ZN(_01719_));
 NAND4_X4 _10708_ (.A1(_01666_),
    .A2(_01613_),
    .A3(_01689_),
    .A4(_01694_),
    .ZN(_01720_));
 BUF_X4 _10709_ (.A(_01720_),
    .Z(_01721_));
 MUX2_X1 _10710_ (.A(_08884_),
    .B(_01719_),
    .S(_01721_),
    .Z(_08911_));
 AOI21_X2 _10711_ (.A(_08903_),
    .B1(_08906_),
    .B2(_08904_),
    .ZN(_01722_));
 OR2_X1 _10712_ (.A1(_08915_),
    .A2(_08914_),
    .ZN(_01723_));
 NAND3_X1 _10713_ (.A1(_08907_),
    .A2(_08904_),
    .A3(_01723_),
    .ZN(_01724_));
 OR3_X1 _10714_ (.A1(_08914_),
    .A2(_01110_),
    .A3(_01368_),
    .ZN(_01725_));
 AOI221_X2 _10715_ (.A(_01725_),
    .B1(_01308_),
    .B2(_01595_),
    .C1(_01710_),
    .C2(_01620_),
    .ZN(_01726_));
 OAI21_X4 _10716_ (.A(_01722_),
    .B1(_01724_),
    .B2(_01726_),
    .ZN(_01727_));
 XOR2_X1 _10717_ (.A(_08913_),
    .B(_01727_),
    .Z(_01728_));
 OAI211_X4 _10718_ (.A(_01556_),
    .B(_01587_),
    .C1(_01618_),
    .C2(_01624_),
    .ZN(_01729_));
 NOR3_X1 _10719_ (.A1(_01647_),
    .A2(_01671_),
    .A3(_01576_),
    .ZN(_01730_));
 AOI21_X1 _10720_ (.A(_01556_),
    .B1(_01674_),
    .B2(_01586_),
    .ZN(_01731_));
 AOI221_X2 _10721_ (.A(_01087_),
    .B1(_01556_),
    .B2(_01730_),
    .C1(_01731_),
    .C2(_01576_),
    .ZN(_01732_));
 NOR3_X1 _10722_ (.A1(_01647_),
    .A2(_01671_),
    .A3(_01583_),
    .ZN(_01733_));
 XNOR2_X1 _10723_ (.A(_01115_),
    .B(_01636_),
    .ZN(_01734_));
 AOI21_X1 _10724_ (.A(_01636_),
    .B1(_01674_),
    .B2(_01586_),
    .ZN(_01735_));
 AOI221_X2 _10725_ (.A(_01119_),
    .B1(_01733_),
    .B2(_01734_),
    .C1(_01735_),
    .C2(_01583_),
    .ZN(_01736_));
 NOR3_X2 _10726_ (.A1(_01691_),
    .A2(_01732_),
    .A3(_01736_),
    .ZN(_01737_));
 NOR3_X2 _10727_ (.A1(_01685_),
    .A2(_01577_),
    .A3(_01636_),
    .ZN(_01738_));
 NOR2_X2 _10728_ (.A1(_01618_),
    .A2(_01624_),
    .ZN(_01739_));
 AOI21_X4 _10729_ (.A(_01737_),
    .B1(_01738_),
    .B2(_01739_),
    .ZN(_01740_));
 INV_X1 _10730_ (.A(_08897_),
    .ZN(_01741_));
 INV_X1 _10731_ (.A(_08882_),
    .ZN(_01742_));
 OAI21_X1 _10732_ (.A(_08889_),
    .B1(_08891_),
    .B2(_01597_),
    .ZN(_01743_));
 NAND2_X1 _10733_ (.A1(_01594_),
    .A2(_01743_),
    .ZN(_01744_));
 AOI21_X1 _10734_ (.A(_08885_),
    .B1(_01744_),
    .B2(_08886_),
    .ZN(_01745_));
 INV_X1 _10735_ (.A(_08883_),
    .ZN(_01746_));
 OAI21_X1 _10736_ (.A(_01742_),
    .B1(_01745_),
    .B2(_01746_),
    .ZN(_01747_));
 AOI21_X2 _10737_ (.A(_08900_),
    .B1(_01747_),
    .B2(_08901_),
    .ZN(_01748_));
 INV_X1 _10738_ (.A(_08898_),
    .ZN(_01749_));
 OAI21_X1 _10739_ (.A(_01741_),
    .B1(_01748_),
    .B2(_01749_),
    .ZN(_01750_));
 AOI21_X2 _10740_ (.A(_08894_),
    .B1(_01750_),
    .B2(_08895_),
    .ZN(_01751_));
 NOR2_X1 _10741_ (.A1(_01119_),
    .A2(_01751_),
    .ZN(_01752_));
 OAI21_X1 _10742_ (.A(_01116_),
    .B1(_01087_),
    .B2(_01751_),
    .ZN(_01753_));
 MUX2_X1 _10743_ (.A(_08869_),
    .B(_01590_),
    .S(_01588_),
    .Z(_01754_));
 MUX2_X1 _10744_ (.A(_01752_),
    .B(_01753_),
    .S(_01754_),
    .Z(_01755_));
 OAI221_X2 _10745_ (.A(_01692_),
    .B1(_01729_),
    .B2(_01691_),
    .C1(_01740_),
    .C2(_01755_),
    .ZN(_01756_));
 OR3_X1 _10746_ (.A1(net10),
    .A2(_01664_),
    .A3(_01665_),
    .ZN(_01757_));
 OR3_X1 _10747_ (.A1(_01649_),
    .A2(_01609_),
    .A3(_01612_),
    .ZN(_01758_));
 NAND2_X1 _10748_ (.A1(_01757_),
    .A2(_01758_),
    .ZN(_01759_));
 AOI221_X2 _10749_ (.A(_01691_),
    .B1(_01676_),
    .B2(_01584_),
    .C1(_01674_),
    .C2(_01586_),
    .ZN(_01760_));
 NAND2_X1 _10750_ (.A1(_01584_),
    .A2(_01676_),
    .ZN(_01761_));
 NOR4_X1 _10751_ (.A1(_01647_),
    .A2(_01671_),
    .A3(_01691_),
    .A4(_01761_),
    .ZN(_01762_));
 OAI22_X1 _10752_ (.A1(_01636_),
    .A2(_01648_),
    .B1(_01760_),
    .B2(_01762_),
    .ZN(_01763_));
 NAND2_X1 _10753_ (.A1(_01586_),
    .A2(_01674_),
    .ZN(_01764_));
 NAND3_X1 _10754_ (.A1(_01764_),
    .A2(_01691_),
    .A3(_01761_),
    .ZN(_01765_));
 OAI21_X1 _10755_ (.A(_01763_),
    .B1(_01765_),
    .B2(_01729_),
    .ZN(_01766_));
 NOR2_X1 _10756_ (.A1(_01440_),
    .A2(net4),
    .ZN(_01767_));
 AOI21_X1 _10757_ (.A(_01767_),
    .B1(_01690_),
    .B2(_01440_),
    .ZN(_01768_));
 OR3_X1 _10758_ (.A1(_01764_),
    .A2(_01768_),
    .A3(_01761_),
    .ZN(_01769_));
 OAI22_X2 _10759_ (.A1(_01764_),
    .A2(net10),
    .B1(_01769_),
    .B2(_01693_),
    .ZN(_01770_));
 AOI211_X2 _10760_ (.A(_01766_),
    .B(_01770_),
    .C1(_01689_),
    .C2(_01694_),
    .ZN(_01771_));
 NAND2_X1 _10761_ (.A1(_01636_),
    .A2(_01648_),
    .ZN(_01772_));
 AND2_X1 _10762_ (.A1(_01729_),
    .A2(_01772_),
    .ZN(_01773_));
 NOR3_X2 _10763_ (.A1(_01649_),
    .A2(_01609_),
    .A3(_01612_),
    .ZN(_01774_));
 NOR3_X2 _10764_ (.A1(net10),
    .A2(_01664_),
    .A3(_01665_),
    .ZN(_01775_));
 OAI21_X2 _10765_ (.A(_01773_),
    .B1(_01774_),
    .B2(_01775_),
    .ZN(_01776_));
 OAI22_X4 _10766_ (.A1(_01740_),
    .A2(_01759_),
    .B1(_01771_),
    .B2(_01776_),
    .ZN(_01777_));
 XNOR2_X1 _10767_ (.A(_01119_),
    .B(_01751_),
    .ZN(_01778_));
 AND2_X1 _10768_ (.A1(_01754_),
    .A2(_01778_),
    .ZN(_01779_));
 AOI211_X2 _10769_ (.A(_01754_),
    .B(_01778_),
    .C1(_01694_),
    .C2(_01689_),
    .ZN(_01780_));
 AOI21_X1 _10770_ (.A(_01153_),
    .B1(_01603_),
    .B2(_01607_),
    .ZN(_01781_));
 AND4_X1 _10771_ (.A1(_01754_),
    .A2(_01689_),
    .A3(_01694_),
    .A4(_01781_),
    .ZN(_01782_));
 NOR3_X4 _10772_ (.A1(_01779_),
    .A2(_01780_),
    .A3(_01782_),
    .ZN(_01783_));
 INV_X1 _10773_ (.A(_08909_),
    .ZN(_01784_));
 NAND2_X1 _10774_ (.A1(_01724_),
    .A2(_01722_),
    .ZN(_01785_));
 AOI21_X2 _10775_ (.A(_08912_),
    .B1(_08913_),
    .B2(_01785_),
    .ZN(_01786_));
 INV_X1 _10776_ (.A(_08910_),
    .ZN(_01787_));
 OAI21_X2 _10777_ (.A(_01784_),
    .B1(_01787_),
    .B2(_01786_),
    .ZN(_01788_));
 AOI21_X4 _10778_ (.A(_08920_),
    .B1(_08921_),
    .B2(_01788_),
    .ZN(_01789_));
 INV_X4 _10779_ (.A(_01789_),
    .ZN(_01790_));
 AOI21_X2 _10780_ (.A(_08917_),
    .B1(_08918_),
    .B2(_01790_),
    .ZN(_01791_));
 INV_X2 _10781_ (.A(_01791_),
    .ZN(_01792_));
 NAND2_X1 _10782_ (.A1(_01792_),
    .A2(_01087_),
    .ZN(_01793_));
 AND4_X1 _10783_ (.A1(_08918_),
    .A2(_08910_),
    .A3(_08913_),
    .A4(_08921_),
    .ZN(_01794_));
 INV_X1 _10784_ (.A(_08920_),
    .ZN(_01795_));
 AOI21_X1 _10785_ (.A(_08909_),
    .B1(_08912_),
    .B2(_08910_),
    .ZN(_01796_));
 INV_X1 _10786_ (.A(_08921_),
    .ZN(_01797_));
 OAI21_X1 _10787_ (.A(_01795_),
    .B1(_01796_),
    .B2(_01797_),
    .ZN(_01798_));
 AOI221_X2 _10788_ (.A(_08917_),
    .B1(_01794_),
    .B2(_01727_),
    .C1(_01798_),
    .C2(_08918_),
    .ZN(_01799_));
 OAI21_X2 _10789_ (.A(_01116_),
    .B1(_01087_),
    .B2(_01799_),
    .ZN(_01800_));
 INV_X1 _10790_ (.A(_01800_),
    .ZN(_01801_));
 XNOR2_X1 _10791_ (.A(_01248_),
    .B(_01385_),
    .ZN(_01802_));
 NOR2_X1 _10792_ (.A1(_01411_),
    .A2(_01802_),
    .ZN(_01803_));
 XNOR2_X1 _10793_ (.A(_01463_),
    .B(_01803_),
    .ZN(_08843_));
 NAND2_X1 _10794_ (.A1(_01443_),
    .A2(_01448_),
    .ZN(_01804_));
 XNOR2_X1 _10795_ (.A(_01442_),
    .B(_01804_),
    .ZN(_01805_));
 MUX2_X1 _10796_ (.A(_08843_),
    .B(_01805_),
    .S(_01660_),
    .Z(_08872_));
 INV_X1 _10797_ (.A(_08872_),
    .ZN(_01806_));
 XNOR2_X1 _10798_ (.A(_01573_),
    .B(_01572_),
    .ZN(_01807_));
 MUX2_X2 _10799_ (.A(_01806_),
    .B(_01807_),
    .S(_01589_),
    .Z(_01808_));
 INV_X4 _10800_ (.A(_01808_),
    .ZN(_08893_));
 MUX2_X1 _10801_ (.A(_01793_),
    .B(_01801_),
    .S(_08893_),
    .Z(_01809_));
 INV_X1 _10802_ (.A(_08900_),
    .ZN(_01810_));
 OAI21_X1 _10803_ (.A(_01810_),
    .B1(_01602_),
    .B2(_01592_),
    .ZN(_01811_));
 AOI21_X2 _10804_ (.A(_08897_),
    .B1(_01811_),
    .B2(_08898_),
    .ZN(_01812_));
 XOR2_X2 _10805_ (.A(_08895_),
    .B(_01812_),
    .Z(_01813_));
 INV_X1 _10806_ (.A(_01813_),
    .ZN(_01814_));
 XNOR2_X1 _10807_ (.A(_01087_),
    .B(_01813_),
    .ZN(_01815_));
 AOI22_X1 _10808_ (.A1(_01153_),
    .A2(_01814_),
    .B1(_01792_),
    .B2(_01815_),
    .ZN(_01816_));
 MUX2_X2 _10809_ (.A(_01809_),
    .B(_01816_),
    .S(_01720_),
    .Z(_01817_));
 NAND4_X4 _10810_ (.A1(_01756_),
    .A2(_01777_),
    .A3(_01783_),
    .A4(_01817_),
    .ZN(_01818_));
 BUF_X4 _10811_ (.A(_01818_),
    .Z(_01819_));
 MUX2_X1 _10812_ (.A(_08911_),
    .B(_01728_),
    .S(_01819_),
    .Z(_08928_));
 INV_X1 _10813_ (.A(_08932_),
    .ZN(_01820_));
 INV_X1 _10814_ (.A(_08938_),
    .ZN(_01821_));
 OAI21_X2 _10815_ (.A(_08939_),
    .B1(_08942_),
    .B2(_08941_),
    .ZN(_01822_));
 NAND2_X2 _10816_ (.A1(_01822_),
    .A2(_01821_),
    .ZN(_01823_));
 AND2_X4 _10817_ (.A1(_08936_),
    .A2(_01823_),
    .ZN(_01824_));
 OAI21_X4 _10818_ (.A(_08933_),
    .B1(_01824_),
    .B2(_08935_),
    .ZN(_01825_));
 NAND2_X4 _10819_ (.A1(_01820_),
    .A2(_01825_),
    .ZN(_01826_));
 XOR2_X1 _10820_ (.A(_08930_),
    .B(_01826_),
    .Z(_01827_));
 OR3_X2 _10821_ (.A1(_01779_),
    .A2(_01780_),
    .A3(_01782_),
    .ZN(_01828_));
 NOR2_X1 _10822_ (.A1(_01120_),
    .A2(_01791_),
    .ZN(_01829_));
 MUX2_X1 _10823_ (.A(_01829_),
    .B(_01800_),
    .S(_08893_),
    .Z(_01830_));
 XNOR2_X1 _10824_ (.A(_01119_),
    .B(_01813_),
    .ZN(_01831_));
 OAI22_X1 _10825_ (.A1(_01116_),
    .A2(_01813_),
    .B1(_01791_),
    .B2(_01831_),
    .ZN(_01832_));
 MUX2_X2 _10826_ (.A(_01830_),
    .B(_01832_),
    .S(_01720_),
    .Z(_01833_));
 NOR2_X4 _10827_ (.A1(_01828_),
    .A2(_01833_),
    .ZN(_01834_));
 NOR2_X1 _10828_ (.A1(_01311_),
    .A2(_01111_),
    .ZN(_01835_));
 OAI21_X1 _10829_ (.A(_01109_),
    .B1(_01179_),
    .B2(net36),
    .ZN(_01836_));
 AND3_X1 _10830_ (.A1(_08907_),
    .A2(_08904_),
    .A3(_08915_),
    .ZN(_01837_));
 AND4_X1 _10831_ (.A1(_01835_),
    .A2(_01836_),
    .A3(_01794_),
    .A4(_01837_),
    .ZN(_01838_));
 NAND2_X1 _10832_ (.A1(_01120_),
    .A2(_01808_),
    .ZN(_01839_));
 OAI21_X1 _10833_ (.A(_01838_),
    .B1(_01839_),
    .B2(net9),
    .ZN(_01840_));
 NAND2_X1 _10834_ (.A1(_01120_),
    .A2(_01813_),
    .ZN(_01841_));
 XNOR2_X2 _10835_ (.A(_01179_),
    .B(net36),
    .ZN(_01842_));
 NAND2_X1 _10836_ (.A1(_01150_),
    .A2(_01842_),
    .ZN(_01843_));
 AOI21_X1 _10837_ (.A(_01696_),
    .B1(_01841_),
    .B2(_01843_),
    .ZN(_01844_));
 MUX2_X2 _10838_ (.A(_01814_),
    .B(_08893_),
    .S(_01696_),
    .Z(_01845_));
 AOI211_X2 _10839_ (.A(_01840_),
    .B(_01844_),
    .C1(_01088_),
    .C2(_01845_),
    .ZN(_01846_));
 NAND2_X1 _10840_ (.A1(_01756_),
    .A2(_01777_),
    .ZN(_01847_));
 OAI21_X2 _10841_ (.A(_01834_),
    .B1(_01846_),
    .B2(_01847_),
    .ZN(_01848_));
 XNOR2_X2 _10842_ (.A(_08918_),
    .B(_01789_),
    .ZN(_01849_));
 INV_X1 _10843_ (.A(_01849_),
    .ZN(_01850_));
 XNOR2_X1 _10844_ (.A(_01087_),
    .B(_01849_),
    .ZN(_01851_));
 INV_X1 _10845_ (.A(_08926_),
    .ZN(_01852_));
 AOI21_X4 _10846_ (.A(_08929_),
    .B1(_08930_),
    .B2(_01826_),
    .ZN(_01853_));
 INV_X1 _10847_ (.A(_08927_),
    .ZN(_01854_));
 OAI21_X4 _10848_ (.A(_01852_),
    .B1(_01853_),
    .B2(_01854_),
    .ZN(_01855_));
 AND2_X4 _10849_ (.A1(_08924_),
    .A2(_01855_),
    .ZN(_01856_));
 NOR2_X4 _10850_ (.A1(_08923_),
    .A2(_01856_),
    .ZN(_01857_));
 OAI22_X2 _10851_ (.A1(_01116_),
    .A2(_01850_),
    .B1(_01851_),
    .B2(_01857_),
    .ZN(_01858_));
 INV_X1 _10852_ (.A(_01858_),
    .ZN(_01859_));
 MUX2_X2 _10853_ (.A(_01813_),
    .B(_01808_),
    .S(_01696_),
    .Z(_01860_));
 XNOR2_X2 _10854_ (.A(_01120_),
    .B(_01799_),
    .ZN(_01861_));
 XNOR2_X1 _10855_ (.A(_01860_),
    .B(_01861_),
    .ZN(_01862_));
 AND3_X1 _10856_ (.A1(_01818_),
    .A2(_01859_),
    .A3(_01862_),
    .ZN(_01863_));
 NOR2_X2 _10857_ (.A1(_01120_),
    .A2(_01857_),
    .ZN(_01864_));
 OAI21_X1 _10858_ (.A(_01116_),
    .B1(_01857_),
    .B2(_01087_),
    .ZN(_01865_));
 NOR2_X2 _10859_ (.A1(_01237_),
    .A2(_01297_),
    .ZN(_08813_));
 NOR2_X1 _10860_ (.A1(_01309_),
    .A2(_08813_),
    .ZN(_01866_));
 INV_X1 _10861_ (.A(_01308_),
    .ZN(_01867_));
 OR3_X1 _10862_ (.A1(_08818_),
    .A2(_08815_),
    .A3(_08817_),
    .ZN(_01868_));
 AOI21_X1 _10863_ (.A(_01867_),
    .B1(_01868_),
    .B2(_01265_),
    .ZN(_01869_));
 NOR2_X1 _10864_ (.A1(_01866_),
    .A2(_01869_),
    .ZN(_08832_));
 XOR2_X1 _10865_ (.A(_08834_),
    .B(_01324_),
    .Z(_01870_));
 MUX2_X1 _10866_ (.A(_08832_),
    .B(_01870_),
    .S(_01368_),
    .Z(_08858_));
 OR3_X1 _10867_ (.A1(_08860_),
    .A2(_08847_),
    .A3(_01447_),
    .ZN(_01871_));
 AND2_X1 _10868_ (.A1(_01448_),
    .A2(_01871_),
    .ZN(_01872_));
 MUX2_X1 _10869_ (.A(_08858_),
    .B(_01872_),
    .S(_01660_),
    .Z(_08875_));
 XOR2_X1 _10870_ (.A(_08877_),
    .B(_01571_),
    .Z(_01873_));
 MUX2_X1 _10871_ (.A(_08875_),
    .B(_01873_),
    .S(_01589_),
    .Z(_08896_));
 XNOR2_X1 _10872_ (.A(_08898_),
    .B(_01748_),
    .ZN(_01874_));
 MUX2_X2 _10873_ (.A(_08896_),
    .B(_01874_),
    .S(_01720_),
    .Z(_08916_));
 MUX2_X1 _10874_ (.A(_01864_),
    .B(_01865_),
    .S(_08916_),
    .Z(_01875_));
 NOR3_X4 _10875_ (.A1(_01818_),
    .A2(_01875_),
    .A3(_01845_),
    .ZN(_01876_));
 OAI221_X2 _10876_ (.A(_01848_),
    .B1(_01863_),
    .B2(_01876_),
    .C1(_01817_),
    .C2(_01783_),
    .ZN(_01877_));
 AND4_X1 _10877_ (.A1(_08939_),
    .A2(_08942_),
    .A3(_08924_),
    .A4(_08936_),
    .ZN(_01878_));
 NAND4_X2 _10878_ (.A1(_08927_),
    .A2(_08930_),
    .A3(_08933_),
    .A4(_01878_),
    .ZN(_01879_));
 AND4_X4 _10879_ (.A1(_01756_),
    .A2(_01777_),
    .A3(_01783_),
    .A4(_01817_),
    .ZN(_01880_));
 NAND2_X1 _10880_ (.A1(_01710_),
    .A2(_01519_),
    .ZN(_01881_));
 OR2_X2 _10881_ (.A1(_01368_),
    .A2(_01881_),
    .ZN(_01882_));
 OAI21_X4 _10882_ (.A(_01711_),
    .B1(_01880_),
    .B2(_01882_),
    .ZN(_01883_));
 XNOR2_X1 _10883_ (.A(_01088_),
    .B(_08916_),
    .ZN(_01884_));
 MUX2_X1 _10884_ (.A(_01851_),
    .B(_01884_),
    .S(_01880_),
    .Z(_01885_));
 NOR4_X4 _10885_ (.A1(_01170_),
    .A2(_01879_),
    .A3(_01883_),
    .A4(_01885_),
    .ZN(_01886_));
 NAND2_X1 _10886_ (.A1(_01729_),
    .A2(_01772_),
    .ZN(_01887_));
 NAND2_X1 _10887_ (.A1(net10),
    .A2(_01761_),
    .ZN(_01888_));
 XNOR2_X2 _10888_ (.A(_01685_),
    .B(_01888_),
    .ZN(_01889_));
 NOR3_X2 _10889_ (.A1(_01755_),
    .A2(_01889_),
    .A3(_01696_),
    .ZN(_01890_));
 XNOR2_X1 _10890_ (.A(_01887_),
    .B(_01890_),
    .ZN(_01891_));
 NOR2_X1 _10891_ (.A1(_01691_),
    .A2(_01729_),
    .ZN(_01892_));
 AND2_X1 _10892_ (.A1(_01768_),
    .A2(_01692_),
    .ZN(_01893_));
 OAI21_X1 _10893_ (.A(_01689_),
    .B1(_01774_),
    .B2(_01775_),
    .ZN(_01894_));
 MUX2_X1 _10894_ (.A(_01893_),
    .B(_01691_),
    .S(_01894_),
    .Z(_01895_));
 AOI21_X2 _10895_ (.A(_01892_),
    .B1(_01895_),
    .B2(_01693_),
    .ZN(_01896_));
 NAND2_X1 _10896_ (.A1(_01891_),
    .A2(_01896_),
    .ZN(_01897_));
 AOI22_X2 _10897_ (.A1(_01757_),
    .A2(_01758_),
    .B1(_01689_),
    .B2(_01694_),
    .ZN(_01898_));
 XNOR2_X2 _10898_ (.A(_01889_),
    .B(_01898_),
    .ZN(_01899_));
 NOR2_X1 _10899_ (.A1(_01120_),
    .A2(_01799_),
    .ZN(_01900_));
 NAND2_X1 _10900_ (.A1(_01813_),
    .A2(_01900_),
    .ZN(_01901_));
 NAND2_X1 _10901_ (.A1(_01808_),
    .A2(_01900_),
    .ZN(_01902_));
 MUX2_X1 _10902_ (.A(_01901_),
    .B(_01902_),
    .S(_01696_),
    .Z(_01903_));
 NAND2_X1 _10903_ (.A1(_08893_),
    .A2(_01800_),
    .ZN(_01904_));
 NAND2_X1 _10904_ (.A1(_01814_),
    .A2(_01800_),
    .ZN(_01905_));
 MUX2_X1 _10905_ (.A(_01904_),
    .B(_01905_),
    .S(_01720_),
    .Z(_01906_));
 AND3_X1 _10906_ (.A1(_01783_),
    .A2(_01903_),
    .A3(_01906_),
    .ZN(_01907_));
 AOI21_X4 _10907_ (.A(_01899_),
    .B1(_01818_),
    .B2(_01907_),
    .ZN(_01908_));
 INV_X1 _10908_ (.A(_01899_),
    .ZN(_01909_));
 NAND3_X2 _10909_ (.A1(_01783_),
    .A2(_01903_),
    .A3(_01906_),
    .ZN(_01910_));
 NOR3_X4 _10910_ (.A1(_01909_),
    .A2(_01880_),
    .A3(_01910_),
    .ZN(_01911_));
 AOI21_X4 _10911_ (.A(_01756_),
    .B1(_01777_),
    .B2(_01834_),
    .ZN(_01912_));
 OR4_X4 _10912_ (.A1(_01897_),
    .A2(_01908_),
    .A3(_01911_),
    .A4(_01912_),
    .ZN(_01913_));
 OR3_X4 _10913_ (.A1(_01877_),
    .A2(_01886_),
    .A3(_01913_),
    .ZN(_01914_));
 BUF_X4 clone33 (.A(_01914_),
    .Z(net33));
 BUF_X8 _10915_ (.A(_01914_),
    .Z(_01916_));
 MUX2_X1 _10916_ (.A(_08928_),
    .B(_01827_),
    .S(net33),
    .Z(_08946_));
 BUF_X1 _10917_ (.A(_08948_),
    .Z(_01917_));
 INV_X1 _10918_ (.A(_08953_),
    .ZN(_01918_));
 INV_X1 _10919_ (.A(_08959_),
    .ZN(_01919_));
 BUF_X1 _10920_ (.A(_08962_),
    .Z(_01920_));
 OAI21_X2 _10921_ (.A(_08960_),
    .B1(_01920_),
    .B2(_08961_),
    .ZN(_01921_));
 NAND2_X2 _10922_ (.A1(_01921_),
    .A2(_01919_),
    .ZN(_01922_));
 AND2_X4 _10923_ (.A1(_08957_),
    .A2(_01922_),
    .ZN(_01923_));
 OAI21_X4 _10924_ (.A(_08954_),
    .B1(_01923_),
    .B2(_08956_),
    .ZN(_01924_));
 NAND2_X4 _10925_ (.A1(_01918_),
    .A2(_01924_),
    .ZN(_01925_));
 BUF_X1 _10926_ (.A(_08951_),
    .Z(_01926_));
 AOI21_X4 _10927_ (.A(_08950_),
    .B1(_01926_),
    .B2(_01925_),
    .ZN(_01927_));
 XNOR2_X1 _10928_ (.A(_01917_),
    .B(_01927_),
    .ZN(_01928_));
 BUF_X4 _10929_ (.A(_01203_),
    .Z(_01929_));
 AND3_X2 _10930_ (.A1(_08818_),
    .A2(_01519_),
    .A3(_01309_),
    .ZN(_01930_));
 AOI21_X2 _10931_ (.A(_01930_),
    .B1(_01867_),
    .B2(_01179_),
    .ZN(_01931_));
 AOI21_X1 _10932_ (.A(_08740_),
    .B1(_01309_),
    .B2(_01929_),
    .ZN(_01932_));
 OAI22_X2 _10933_ (.A1(_01929_),
    .A2(_01931_),
    .B1(_01932_),
    .B2(_08818_),
    .ZN(_08835_));
 INV_X1 _10934_ (.A(_08837_),
    .ZN(_01933_));
 XNOR2_X1 _10935_ (.A(_01933_),
    .B(_01382_),
    .ZN(_01934_));
 MUX2_X1 _10936_ (.A(_08835_),
    .B(_01934_),
    .S(_01368_),
    .Z(_08846_));
 XOR2_X1 _10937_ (.A(_08848_),
    .B(_01446_),
    .Z(_01935_));
 MUX2_X1 _10938_ (.A(_08846_),
    .B(_01935_),
    .S(_01660_),
    .Z(_08878_));
 OR3_X1 _10939_ (.A1(_08880_),
    .A2(_08862_),
    .A3(_01569_),
    .ZN(_01936_));
 AND2_X1 _10940_ (.A1(_01570_),
    .A2(_01936_),
    .ZN(_01937_));
 MUX2_X1 _10941_ (.A(_08878_),
    .B(_01937_),
    .S(_01589_),
    .Z(_08899_));
 AOI21_X1 _10942_ (.A(_08885_),
    .B1(_01600_),
    .B2(_08886_),
    .ZN(_01938_));
 OAI21_X1 _10943_ (.A(_01742_),
    .B1(_01938_),
    .B2(_01746_),
    .ZN(_01939_));
 XOR2_X1 _10944_ (.A(_08901_),
    .B(_01939_),
    .Z(_01940_));
 MUX2_X1 _10945_ (.A(_08899_),
    .B(_01940_),
    .S(_01721_),
    .Z(_08919_));
 AOI21_X1 _10946_ (.A(_08912_),
    .B1(_01727_),
    .B2(_08913_),
    .ZN(_01941_));
 OAI21_X1 _10947_ (.A(_01784_),
    .B1(_01941_),
    .B2(_01787_),
    .ZN(_01942_));
 XNOR2_X1 _10948_ (.A(_01797_),
    .B(_01942_),
    .ZN(_01943_));
 MUX2_X1 _10949_ (.A(_08919_),
    .B(_01943_),
    .S(_01819_),
    .Z(_01944_));
 BUF_X2 _10950_ (.A(_01944_),
    .Z(_08922_));
 XNOR2_X1 _10951_ (.A(_01121_),
    .B(_08922_),
    .ZN(_01945_));
 BUF_X2 _10952_ (.A(_08945_),
    .Z(_01946_));
 INV_X1 _10953_ (.A(_08947_),
    .ZN(_01947_));
 INV_X1 _10954_ (.A(_01917_),
    .ZN(_01948_));
 OAI21_X4 _10955_ (.A(_01947_),
    .B1(_01927_),
    .B2(_01948_),
    .ZN(_01949_));
 AND2_X4 _10956_ (.A1(_01949_),
    .A2(_01946_),
    .ZN(_01950_));
 OR2_X2 _10957_ (.A1(_01950_),
    .A2(_08944_),
    .ZN(_01951_));
 AOI22_X2 _10958_ (.A1(_01153_),
    .A2(_08922_),
    .B1(_01951_),
    .B2(_01945_),
    .ZN(_01952_));
 NOR2_X4 _10959_ (.A1(_01950_),
    .A2(_08944_),
    .ZN(_01953_));
 XOR2_X2 _10960_ (.A(_08924_),
    .B(_01855_),
    .Z(_01954_));
 NOR2_X1 _10961_ (.A1(_01121_),
    .A2(_01954_),
    .ZN(_01955_));
 INV_X1 _10962_ (.A(_01954_),
    .ZN(_01956_));
 NOR2_X1 _10963_ (.A1(_01088_),
    .A2(_01956_),
    .ZN(_01957_));
 NOR2_X1 _10964_ (.A1(_01955_),
    .A2(_01957_),
    .ZN(_01958_));
 NOR2_X1 _10965_ (.A1(_01953_),
    .A2(_01958_),
    .ZN(_01959_));
 BUF_X4 _10966_ (.A(_01153_),
    .Z(_01960_));
 AOI21_X1 _10967_ (.A(_01959_),
    .B1(_01954_),
    .B2(_01960_),
    .ZN(_01961_));
 MUX2_X2 _10968_ (.A(_01952_),
    .B(_01961_),
    .S(_01914_),
    .Z(_01962_));
 NOR3_X1 _10969_ (.A1(_08923_),
    .A2(_01120_),
    .A3(_01856_),
    .ZN(_01963_));
 XNOR2_X1 _10970_ (.A(_01153_),
    .B(_01845_),
    .ZN(_01964_));
 BUF_X4 _10971_ (.A(_01880_),
    .Z(_01965_));
 OAI21_X1 _10972_ (.A(_01964_),
    .B1(_01861_),
    .B2(_01965_),
    .ZN(_01966_));
 OR3_X1 _10973_ (.A1(_01965_),
    .A2(_01861_),
    .A3(_01964_),
    .ZN(_01967_));
 MUX2_X2 _10974_ (.A(_01849_),
    .B(_08916_),
    .S(_01965_),
    .Z(_01968_));
 NAND4_X2 _10975_ (.A1(_01963_),
    .A2(_01966_),
    .A3(_01967_),
    .A4(_01968_),
    .ZN(_01969_));
 OAI21_X2 _10976_ (.A(_01845_),
    .B1(_01965_),
    .B2(_01861_),
    .ZN(_01970_));
 XNOR2_X2 _10977_ (.A(_01088_),
    .B(_01799_),
    .ZN(_01971_));
 NAND3_X2 _10978_ (.A1(_01860_),
    .A2(_01819_),
    .A3(_01971_),
    .ZN(_01972_));
 INV_X1 _10979_ (.A(_08916_),
    .ZN(_01973_));
 MUX2_X2 _10980_ (.A(_01850_),
    .B(_01973_),
    .S(_01965_),
    .Z(_01974_));
 NAND4_X2 _10981_ (.A1(_01864_),
    .A2(_01970_),
    .A3(_01972_),
    .A4(_01974_),
    .ZN(_01975_));
 AOI21_X1 _10982_ (.A(_01845_),
    .B1(_01819_),
    .B2(_01971_),
    .ZN(_01976_));
 NOR3_X1 _10983_ (.A1(_01860_),
    .A2(_01965_),
    .A3(_01861_),
    .ZN(_01977_));
 NAND2_X1 _10984_ (.A1(_01120_),
    .A2(_01857_),
    .ZN(_01978_));
 OR4_X1 _10985_ (.A1(_01976_),
    .A2(_01977_),
    .A3(_01968_),
    .A4(_01978_),
    .ZN(_01979_));
 NOR2_X1 _10986_ (.A1(_01088_),
    .A2(_01857_),
    .ZN(_01980_));
 NAND4_X2 _10987_ (.A1(_01980_),
    .A2(_01970_),
    .A3(_01972_),
    .A4(_01968_),
    .ZN(_01981_));
 NAND4_X4 _10988_ (.A1(_01969_),
    .A2(_01975_),
    .A3(_01979_),
    .A4(_01981_),
    .ZN(_01982_));
 OR2_X1 _10989_ (.A1(_01864_),
    .A2(_01968_),
    .ZN(_01983_));
 NOR4_X4 _10990_ (.A1(_01877_),
    .A2(_01886_),
    .A3(_01913_),
    .A4(_01983_),
    .ZN(_01984_));
 OR2_X4 _10991_ (.A1(_01982_),
    .A2(_01984_),
    .ZN(_01985_));
 NOR2_X2 _10992_ (.A1(_01863_),
    .A2(_01876_),
    .ZN(_01986_));
 NOR2_X1 _10993_ (.A1(_01818_),
    .A2(_01875_),
    .ZN(_01987_));
 NAND2_X2 _10994_ (.A1(_01828_),
    .A2(_01833_),
    .ZN(_01988_));
 AOI221_X2 _10995_ (.A(_01863_),
    .B1(_01987_),
    .B2(_01860_),
    .C1(_01848_),
    .C2(_01988_),
    .ZN(_01989_));
 OR2_X2 _10996_ (.A1(_01908_),
    .A2(_01911_),
    .ZN(_01990_));
 INV_X1 _10997_ (.A(_01988_),
    .ZN(_01991_));
 NAND3_X1 _10998_ (.A1(_01818_),
    .A2(_01859_),
    .A3(_01862_),
    .ZN(_01992_));
 OR3_X1 _10999_ (.A1(_01845_),
    .A2(_01818_),
    .A3(_01875_),
    .ZN(_01993_));
 AND2_X1 _11000_ (.A1(_01756_),
    .A2(_01777_),
    .ZN(_01994_));
 NAND4_X1 _11001_ (.A1(_01835_),
    .A2(_01836_),
    .A3(_01794_),
    .A4(_01837_),
    .ZN(_01995_));
 NOR2_X1 _11002_ (.A1(_01088_),
    .A2(_08893_),
    .ZN(_01996_));
 AOI21_X1 _11003_ (.A(_01995_),
    .B1(_01996_),
    .B2(_01696_),
    .ZN(_01997_));
 NOR2_X1 _11004_ (.A1(_01088_),
    .A2(_01814_),
    .ZN(_01998_));
 AND2_X1 _11005_ (.A1(_01150_),
    .A2(_01842_),
    .ZN(_01999_));
 OAI21_X1 _11006_ (.A(net9),
    .B1(_01998_),
    .B2(_01999_),
    .ZN(_02000_));
 OAI211_X2 _11007_ (.A(_01997_),
    .B(_02000_),
    .C1(_01120_),
    .C2(_01860_),
    .ZN(_02001_));
 NAND2_X1 _11008_ (.A1(_01994_),
    .A2(_02001_),
    .ZN(_02002_));
 AOI221_X2 _11009_ (.A(_01991_),
    .B1(_01992_),
    .B2(_01993_),
    .C1(_01834_),
    .C2(_02002_),
    .ZN(_02003_));
 OAI33_X1 _11010_ (.A1(_01986_),
    .A2(_01886_),
    .A3(_01913_),
    .B1(_01989_),
    .B2(_01990_),
    .B3(_02003_),
    .ZN(_02004_));
 NOR4_X2 _11011_ (.A1(_01887_),
    .A2(_01909_),
    .A3(_01965_),
    .A4(_01910_),
    .ZN(_02005_));
 XNOR2_X2 _11012_ (.A(_01896_),
    .B(_02005_),
    .ZN(_02006_));
 XNOR2_X2 _11013_ (.A(_01773_),
    .B(_01890_),
    .ZN(_02007_));
 OR3_X2 _11014_ (.A1(_02007_),
    .A2(_01908_),
    .A3(_01911_),
    .ZN(_02008_));
 OAI21_X4 _11015_ (.A(_02006_),
    .B1(_02008_),
    .B2(_01877_),
    .ZN(_02009_));
 INV_X1 _11016_ (.A(_01912_),
    .ZN(_02010_));
 NAND3_X1 _11017_ (.A1(_01899_),
    .A2(_01783_),
    .A3(_01817_),
    .ZN(_02011_));
 AOI21_X2 _11018_ (.A(_02011_),
    .B1(_02001_),
    .B2(_01994_),
    .ZN(_02012_));
 XNOR2_X2 _11019_ (.A(_02007_),
    .B(_02012_),
    .ZN(_02013_));
 AND2_X2 _11020_ (.A1(_02010_),
    .A2(_02013_),
    .ZN(_02014_));
 AND3_X2 _11021_ (.A1(net381),
    .A2(_02009_),
    .A3(_02014_),
    .ZN(_02015_));
 NAND3_X4 _11022_ (.A1(_02015_),
    .A2(_01962_),
    .A3(_01985_),
    .ZN(_02016_));
 BUF_X8 _11023_ (.A(_02016_),
    .Z(_02017_));
 MUX2_X2 _11024_ (.A(_08946_),
    .B(_01928_),
    .S(_02017_),
    .Z(_08963_));
 NAND2_X1 _11025_ (.A1(_01137_),
    .A2(_08963_),
    .ZN(_02018_));
 OR2_X2 _11026_ (.A1(_01886_),
    .A2(_01913_),
    .ZN(_02019_));
 NOR2_X2 _11027_ (.A1(_01986_),
    .A2(_02019_),
    .ZN(_02020_));
 NOR3_X2 _11028_ (.A1(_02003_),
    .A2(_01990_),
    .A3(_01989_),
    .ZN(_02021_));
 NOR2_X4 _11029_ (.A1(_02020_),
    .A2(_02021_),
    .ZN(_02022_));
 NAND3_X4 _11030_ (.A1(net381),
    .A2(_02009_),
    .A3(_02014_),
    .ZN(_02023_));
 INV_X1 _11031_ (.A(_08922_),
    .ZN(_02024_));
 NOR2_X1 _11032_ (.A1(_01088_),
    .A2(_02024_),
    .ZN(_02025_));
 MUX2_X2 _11033_ (.A(_02025_),
    .B(_01957_),
    .S(_01914_),
    .Z(_02026_));
 NOR2_X1 _11034_ (.A1(_01121_),
    .A2(_08922_),
    .ZN(_02027_));
 MUX2_X2 _11035_ (.A(_02027_),
    .B(_01955_),
    .S(_01914_),
    .Z(_02028_));
 NOR3_X4 _11036_ (.A1(_02023_),
    .A2(_02026_),
    .A3(_02028_),
    .ZN(_02029_));
 NOR2_X1 _11037_ (.A1(_01170_),
    .A2(_01883_),
    .ZN(_02030_));
 NAND4_X1 _11038_ (.A1(_08960_),
    .A2(_01920_),
    .A3(_01946_),
    .A4(_08957_),
    .ZN(_02031_));
 NAND3_X1 _11039_ (.A1(_01917_),
    .A2(_01926_),
    .A3(_08954_),
    .ZN(_02032_));
 NOR2_X1 _11040_ (.A1(_02031_),
    .A2(_02032_),
    .ZN(_02033_));
 AND3_X1 _11041_ (.A1(_02030_),
    .A2(_02004_),
    .A3(_02033_),
    .ZN(_02034_));
 OAI221_X2 _11042_ (.A(_01962_),
    .B1(_01982_),
    .B2(_01984_),
    .C1(_02023_),
    .C2(_02034_),
    .ZN(_02035_));
 NOR2_X4 _11043_ (.A1(_02029_),
    .A2(_02035_),
    .ZN(_02036_));
 XNOR2_X1 _11044_ (.A(_01088_),
    .B(_08922_),
    .ZN(_02037_));
 OAI22_X1 _11045_ (.A1(_01116_),
    .A2(_02024_),
    .B1(_02037_),
    .B2(_01953_),
    .ZN(_02038_));
 OAI22_X1 _11046_ (.A1(_01116_),
    .A2(_01956_),
    .B1(_01958_),
    .B2(_01953_),
    .ZN(_02039_));
 MUX2_X2 _11047_ (.A(_02038_),
    .B(_02039_),
    .S(_01914_),
    .Z(_02040_));
 OR2_X1 _11048_ (.A1(_01980_),
    .A2(_01963_),
    .ZN(_02041_));
 INV_X1 _11049_ (.A(_02041_),
    .ZN(_02042_));
 NOR3_X2 _11050_ (.A1(_01877_),
    .A2(_01886_),
    .A3(_01913_),
    .ZN(_02043_));
 OAI21_X2 _11051_ (.A(_01974_),
    .B1(_02042_),
    .B2(_02043_),
    .ZN(_02044_));
 NAND3_X2 _11052_ (.A1(net33),
    .A2(_01968_),
    .A3(_02041_),
    .ZN(_02045_));
 AOI21_X4 _11053_ (.A(_02040_),
    .B1(_02044_),
    .B2(_02045_),
    .ZN(_02046_));
 INV_X1 _11054_ (.A(_01986_),
    .ZN(_02047_));
 NAND2_X2 _11055_ (.A1(_01848_),
    .A2(_01988_),
    .ZN(_02048_));
 OAI21_X1 _11056_ (.A(_02047_),
    .B1(_02019_),
    .B2(_02048_),
    .ZN(_02049_));
 NOR2_X1 _11057_ (.A1(_01965_),
    .A2(_01858_),
    .ZN(_02050_));
 OR4_X1 _11058_ (.A1(_01987_),
    .A2(_01976_),
    .A3(_01977_),
    .A4(_02050_),
    .ZN(_02051_));
 AND2_X1 _11059_ (.A1(_02049_),
    .A2(_02051_),
    .ZN(_02052_));
 NOR2_X4 _11060_ (.A1(_02046_),
    .A2(_02052_),
    .ZN(_02053_));
 OR3_X4 _11061_ (.A1(_02022_),
    .A2(_02036_),
    .A3(_02053_),
    .ZN(_02054_));
 MUX2_X2 _11062_ (.A(_02024_),
    .B(_01956_),
    .S(net33),
    .Z(_02055_));
 XNOR2_X2 _11063_ (.A(_01121_),
    .B(_01953_),
    .ZN(_02056_));
 NAND2_X1 _11064_ (.A1(_02055_),
    .A2(_02056_),
    .ZN(_02057_));
 NAND2_X1 _11065_ (.A1(_01985_),
    .A2(_02055_),
    .ZN(_02058_));
 NAND2_X1 _11066_ (.A1(_01962_),
    .A2(_02015_),
    .ZN(_02059_));
 MUX2_X1 _11067_ (.A(_08922_),
    .B(_01954_),
    .S(net33),
    .Z(_02060_));
 XNOR2_X1 _11068_ (.A(_01089_),
    .B(_01953_),
    .ZN(_02061_));
 NAND2_X1 _11069_ (.A1(_02060_),
    .A2(_02061_),
    .ZN(_02062_));
 NOR2_X4 _11070_ (.A1(_01982_),
    .A2(_01984_),
    .ZN(_02063_));
 NOR3_X4 _11071_ (.A1(_02040_),
    .A2(_02063_),
    .A3(_02023_),
    .ZN(_02064_));
 OAI221_X2 _11072_ (.A(_02057_),
    .B1(_02058_),
    .B2(_02059_),
    .C1(_02062_),
    .C2(_02064_),
    .ZN(_02065_));
 AOI21_X2 _11073_ (.A(_01968_),
    .B1(_02041_),
    .B2(net33),
    .ZN(_02066_));
 NOR3_X2 _11074_ (.A1(_02043_),
    .A2(_01974_),
    .A3(_02042_),
    .ZN(_02067_));
 NOR3_X2 _11075_ (.A1(_01962_),
    .A2(_02066_),
    .A3(_02067_),
    .ZN(_02068_));
 OAI21_X4 _11076_ (.A(net28),
    .B1(_02068_),
    .B2(_02046_),
    .ZN(_02069_));
 NOR2_X1 _11077_ (.A1(_08839_),
    .A2(_01411_),
    .ZN(_08852_));
 OR3_X1 _11078_ (.A1(_08854_),
    .A2(_08857_),
    .A3(_08856_),
    .ZN(_02070_));
 AND2_X1 _11079_ (.A1(_01445_),
    .A2(_02070_),
    .ZN(_02071_));
 MUX2_X1 _11080_ (.A(_08852_),
    .B(_02071_),
    .S(_01660_),
    .Z(_08861_));
 XOR2_X1 _11081_ (.A(_08863_),
    .B(_01568_),
    .Z(_02072_));
 MUX2_X1 _11082_ (.A(_08861_),
    .B(_02072_),
    .S(_01589_),
    .Z(_08881_));
 XNOR2_X1 _11083_ (.A(_08883_),
    .B(_01745_),
    .ZN(_02073_));
 MUX2_X1 _11084_ (.A(_08881_),
    .B(_02073_),
    .S(_01721_),
    .Z(_08908_));
 XNOR2_X1 _11085_ (.A(_08910_),
    .B(_01786_),
    .ZN(_02074_));
 MUX2_X1 _11086_ (.A(_08908_),
    .B(_02074_),
    .S(_01819_),
    .Z(_08925_));
 INV_X1 _11087_ (.A(_08925_),
    .ZN(_02075_));
 XNOR2_X1 _11088_ (.A(_01854_),
    .B(_01853_),
    .ZN(_02076_));
 MUX2_X2 _11089_ (.A(_02075_),
    .B(_02076_),
    .S(_01914_),
    .Z(_02077_));
 NAND4_X2 _11090_ (.A1(_01962_),
    .A2(_01985_),
    .A3(_02015_),
    .A4(_02077_),
    .ZN(_02078_));
 XOR2_X2 _11091_ (.A(_01946_),
    .B(_01949_),
    .Z(_02079_));
 BUF_X2 _11092_ (.A(_08964_),
    .Z(_02080_));
 OAI21_X1 _11093_ (.A(_08965_),
    .B1(_01705_),
    .B2(_08967_),
    .ZN(_02081_));
 NOR2_X1 _11094_ (.A1(_08967_),
    .A2(_08970_),
    .ZN(_02082_));
 OAI21_X1 _11095_ (.A(_08971_),
    .B1(_01700_),
    .B2(_01702_),
    .ZN(_02083_));
 AOI21_X2 _11096_ (.A(_02081_),
    .B1(_02082_),
    .B2(_02083_),
    .ZN(_02084_));
 NOR2_X1 _11097_ (.A1(_02080_),
    .A2(_02084_),
    .ZN(_02085_));
 NOR2_X1 _11098_ (.A1(_01089_),
    .A2(_02085_),
    .ZN(_02086_));
 OAI221_X2 _11099_ (.A(_02078_),
    .B1(_02079_),
    .B2(_02064_),
    .C1(_02086_),
    .C2(_01960_),
    .ZN(_02087_));
 INV_X2 _11100_ (.A(_02077_),
    .ZN(_08943_));
 NAND4_X2 _11101_ (.A1(_01962_),
    .A2(_01985_),
    .A3(_02015_),
    .A4(_08943_),
    .ZN(_02088_));
 NOR2_X1 _11102_ (.A1(_01121_),
    .A2(_02085_),
    .ZN(_02089_));
 XNOR2_X2 _11103_ (.A(_01946_),
    .B(_01949_),
    .ZN(_02090_));
 OAI211_X4 _11104_ (.A(_02088_),
    .B(_02089_),
    .C1(_02064_),
    .C2(_02090_),
    .ZN(_02091_));
 NAND4_X4 _11105_ (.A1(_02065_),
    .A2(_02069_),
    .A3(_02087_),
    .A4(_02091_),
    .ZN(_02092_));
 OR2_X1 _11106_ (.A1(_01877_),
    .A2(_02008_),
    .ZN(_02093_));
 OAI21_X1 _11107_ (.A(_01912_),
    .B1(_02006_),
    .B2(_02093_),
    .ZN(_02094_));
 AND3_X1 _11108_ (.A1(net381),
    .A2(_02013_),
    .A3(_02094_),
    .ZN(_02095_));
 NOR2_X2 _11109_ (.A1(_02040_),
    .A2(_02063_),
    .ZN(_02096_));
 AOI22_X4 _11110_ (.A1(_02009_),
    .A2(_02014_),
    .B1(_02095_),
    .B2(_02096_),
    .ZN(_02097_));
 OAI21_X1 _11111_ (.A(net9),
    .B1(net36),
    .B2(_01519_),
    .ZN(_02098_));
 INV_X1 _11112_ (.A(_02098_),
    .ZN(_02099_));
 AOI21_X2 _11113_ (.A(_02099_),
    .B1(net36),
    .B2(_01519_),
    .ZN(_02100_));
 OAI21_X1 _11114_ (.A(_01179_),
    .B1(_01368_),
    .B2(_01819_),
    .ZN(_02101_));
 OAI21_X2 _11115_ (.A(_02101_),
    .B1(_01819_),
    .B2(_01620_),
    .ZN(_02102_));
 BUF_X4 _11116_ (.A(_01110_),
    .Z(_02103_));
 OAI22_X4 _11117_ (.A1(_01929_),
    .A2(_02100_),
    .B1(_02102_),
    .B2(_02103_),
    .ZN(_02104_));
 INV_X1 _11118_ (.A(_08971_),
    .ZN(_02105_));
 NAND4_X1 _11119_ (.A1(_08980_),
    .A2(_01142_),
    .A3(_08965_),
    .A4(_01705_),
    .ZN(_02106_));
 OR4_X4 _11120_ (.A1(_02106_),
    .A2(_01170_),
    .A3(_01141_),
    .A4(_02105_),
    .ZN(_02107_));
 XNOR2_X1 _11121_ (.A(_01696_),
    .B(_01842_),
    .ZN(_02108_));
 OAI22_X2 _11122_ (.A1(_02103_),
    .A2(net11),
    .B1(_02108_),
    .B2(_01929_),
    .ZN(_02109_));
 NAND2_X1 _11123_ (.A1(_01710_),
    .A2(_01819_),
    .ZN(_02110_));
 MUX2_X1 _11124_ (.A(net11),
    .B(_02109_),
    .S(_02110_),
    .Z(_02111_));
 BUF_X4 _11125_ (.A(_02111_),
    .Z(_02112_));
 OR3_X4 _11126_ (.A1(_02107_),
    .A2(_02104_),
    .A3(_02112_),
    .ZN(_02113_));
 NAND2_X1 _11127_ (.A1(_01121_),
    .A2(_02079_),
    .ZN(_02114_));
 NAND2_X1 _11128_ (.A1(_01089_),
    .A2(_02090_),
    .ZN(_02115_));
 AOI221_X2 _11129_ (.A(_02113_),
    .B1(_02114_),
    .B2(_02115_),
    .C1(_02096_),
    .C2(_02015_),
    .ZN(_02116_));
 NOR3_X2 _11130_ (.A1(_02104_),
    .A2(_02107_),
    .A3(_02112_),
    .ZN(_02117_));
 NAND3_X2 _11131_ (.A1(_01121_),
    .A2(_08943_),
    .A3(_02117_),
    .ZN(_02118_));
 NAND3_X2 _11132_ (.A1(_01089_),
    .A2(_02077_),
    .A3(_02117_),
    .ZN(_02119_));
 AOI21_X4 _11133_ (.A(_02016_),
    .B1(_02118_),
    .B2(_02119_),
    .ZN(_02120_));
 OR3_X4 _11134_ (.A1(_02097_),
    .A2(_02116_),
    .A3(_02120_),
    .ZN(_02121_));
 NOR3_X4 _11135_ (.A1(_02054_),
    .A2(_02092_),
    .A3(_02121_),
    .ZN(_02122_));
 MUX2_X2 _11136_ (.A(_01709_),
    .B(_02018_),
    .S(_02122_),
    .Z(_02123_));
 NOR3_X4 _11137_ (.A1(_02022_),
    .A2(_02036_),
    .A3(_02053_),
    .ZN(_02124_));
 AND4_X2 _11138_ (.A1(_02065_),
    .A2(_02069_),
    .A3(_02087_),
    .A4(_02091_),
    .ZN(_02125_));
 BUF_X4 _11139_ (.A(_02125_),
    .Z(_02126_));
 NOR3_X4 _11140_ (.A1(_02097_),
    .A2(_02116_),
    .A3(_02120_),
    .ZN(_02127_));
 NAND2_X4 _11141_ (.A1(_01089_),
    .A2(_01135_),
    .ZN(_02128_));
 NOR2_X1 _11142_ (.A1(_08963_),
    .A2(_02128_),
    .ZN(_02129_));
 AND4_X1 _11143_ (.A1(_02124_),
    .A2(_02126_),
    .A3(_02127_),
    .A4(_02129_),
    .ZN(_02130_));
 NOR2_X4 _11144_ (.A1(_01708_),
    .A2(_02128_),
    .ZN(_02131_));
 NAND3_X4 _11145_ (.A1(_02124_),
    .A2(_02125_),
    .A3(_02127_),
    .ZN(_02132_));
 AOI21_X4 _11146_ (.A(_02130_),
    .B1(_02131_),
    .B2(net7),
    .ZN(_02133_));
 NOR2_X1 _11147_ (.A1(_02060_),
    .A2(_02061_),
    .ZN(_02134_));
 NOR2_X1 _11148_ (.A1(_02063_),
    .A2(_02060_),
    .ZN(_02135_));
 NOR2_X1 _11149_ (.A1(_02040_),
    .A2(_02023_),
    .ZN(_02136_));
 NOR2_X1 _11150_ (.A1(_02055_),
    .A2(_02056_),
    .ZN(_02137_));
 AOI221_X2 _11151_ (.A(_02134_),
    .B1(_02135_),
    .B2(_02136_),
    .C1(_02137_),
    .C2(net28),
    .ZN(_02138_));
 NOR4_X2 _11152_ (.A1(_02040_),
    .A2(_02063_),
    .A3(_02023_),
    .A4(_02077_),
    .ZN(_02139_));
 INV_X1 _11153_ (.A(_08973_),
    .ZN(_02140_));
 OAI21_X1 _11154_ (.A(_08980_),
    .B1(_01142_),
    .B2(_08982_),
    .ZN(_02141_));
 NAND2_X1 _11155_ (.A1(_01699_),
    .A2(_02141_),
    .ZN(_02142_));
 AOI21_X1 _11156_ (.A(_08976_),
    .B1(_02142_),
    .B2(_08977_),
    .ZN(_02143_));
 INV_X1 _11157_ (.A(_01140_),
    .ZN(_02144_));
 OAI21_X1 _11158_ (.A(_02140_),
    .B1(_02143_),
    .B2(_02144_),
    .ZN(_02145_));
 AOI21_X2 _11159_ (.A(_08970_),
    .B1(_02145_),
    .B2(_08971_),
    .ZN(_02146_));
 OAI21_X1 _11160_ (.A(_01139_),
    .B1(_02146_),
    .B2(_01706_),
    .ZN(_02147_));
 AOI21_X2 _11161_ (.A(_02080_),
    .B1(_02147_),
    .B2(_08965_),
    .ZN(_02148_));
 OR2_X1 _11162_ (.A1(_01121_),
    .A2(_02148_),
    .ZN(_02149_));
 AOI211_X2 _11163_ (.A(_02139_),
    .B(_02149_),
    .C1(net28),
    .C2(_02079_),
    .ZN(_02150_));
 NOR4_X4 _11164_ (.A1(_02040_),
    .A2(_02063_),
    .A3(_02023_),
    .A4(_08943_),
    .ZN(_02151_));
 OR2_X1 _11165_ (.A1(_01089_),
    .A2(_02148_),
    .ZN(_02152_));
 AOI221_X2 _11166_ (.A(_02151_),
    .B1(_02090_),
    .B2(_02016_),
    .C1(_02152_),
    .C2(_01116_),
    .ZN(_02153_));
 NOR3_X2 _11167_ (.A1(_02138_),
    .A2(_02150_),
    .A3(_02153_),
    .ZN(_02154_));
 XNOR2_X1 _11168_ (.A(_02069_),
    .B(_02154_),
    .ZN(_02155_));
 AND2_X2 _11169_ (.A1(_02087_),
    .A2(_02091_),
    .ZN(_02156_));
 XNOR2_X1 _11170_ (.A(_02065_),
    .B(_02156_),
    .ZN(_02157_));
 OAI21_X2 _11171_ (.A(_02132_),
    .B1(_02155_),
    .B2(_02157_),
    .ZN(_02158_));
 AOI21_X4 _11172_ (.A(_02151_),
    .B1(_02090_),
    .B2(net28),
    .ZN(_02159_));
 XNOR2_X2 _11173_ (.A(_01121_),
    .B(_02148_),
    .ZN(_02160_));
 AND2_X1 _11174_ (.A1(_02159_),
    .A2(_02160_),
    .ZN(_02161_));
 NAND3_X2 _11175_ (.A1(_02040_),
    .A2(_02044_),
    .A3(_02045_),
    .ZN(_02162_));
 OAI21_X2 _11176_ (.A(_01962_),
    .B1(_02066_),
    .B2(_02067_),
    .ZN(_02163_));
 AOI21_X4 _11177_ (.A(_02064_),
    .B1(_02162_),
    .B2(_02163_),
    .ZN(_02164_));
 NAND2_X1 _11178_ (.A1(net28),
    .A2(_02137_),
    .ZN(_02165_));
 OAI21_X2 _11179_ (.A(_02055_),
    .B1(_02064_),
    .B2(_02056_),
    .ZN(_02166_));
 AOI221_X2 _11180_ (.A(_02164_),
    .B1(_02165_),
    .B2(_02166_),
    .C1(_01960_),
    .C2(_02159_),
    .ZN(_02167_));
 OAI21_X1 _11181_ (.A(_02078_),
    .B1(_02079_),
    .B2(_02064_),
    .ZN(_02168_));
 OR2_X1 _11182_ (.A1(_02080_),
    .A2(_02084_),
    .ZN(_02169_));
 AOI21_X1 _11183_ (.A(_02168_),
    .B1(_02169_),
    .B2(_01122_),
    .ZN(_02170_));
 AND4_X1 _11184_ (.A1(_02124_),
    .A2(_02167_),
    .A3(_02127_),
    .A4(_02170_),
    .ZN(_02171_));
 NOR2_X1 _11185_ (.A1(_02159_),
    .A2(_02160_),
    .ZN(_02172_));
 AOI211_X2 _11186_ (.A(_02161_),
    .B(_02171_),
    .C1(_02132_),
    .C2(_02172_),
    .ZN(_02173_));
 NAND4_X4 _11187_ (.A1(_02123_),
    .A2(_02133_),
    .A3(_02158_),
    .A4(_02173_),
    .ZN(_02174_));
 NAND2_X2 _11188_ (.A1(net382),
    .A2(_02036_),
    .ZN(_02175_));
 INV_X1 _11189_ (.A(_02013_),
    .ZN(_02176_));
 NOR2_X2 _11190_ (.A1(_01908_),
    .A2(_01911_),
    .ZN(_02177_));
 NAND3_X1 _11191_ (.A1(_02003_),
    .A2(_02177_),
    .A3(_02019_),
    .ZN(_02178_));
 XNOR2_X2 _11192_ (.A(_02176_),
    .B(_02178_),
    .ZN(_02179_));
 XNOR2_X2 _11193_ (.A(_02175_),
    .B(_02179_),
    .ZN(_02180_));
 NOR4_X2 _11194_ (.A1(_02138_),
    .A2(_02164_),
    .A3(_02150_),
    .A4(_02153_),
    .ZN(_02181_));
 NAND2_X1 _11195_ (.A1(_02124_),
    .A2(_02181_),
    .ZN(_02182_));
 NAND4_X2 _11196_ (.A1(_01962_),
    .A2(_01985_),
    .A3(net382),
    .A4(_02013_),
    .ZN(_02183_));
 NAND4_X1 _11197_ (.A1(_08960_),
    .A2(_01926_),
    .A3(_08954_),
    .A4(_08957_),
    .ZN(_02184_));
 NAND3_X1 _11198_ (.A1(_01920_),
    .A2(_01946_),
    .A3(_01917_),
    .ZN(_02185_));
 NOR4_X2 _11199_ (.A1(_01170_),
    .A2(_01883_),
    .A3(_02184_),
    .A4(_02185_),
    .ZN(_02186_));
 OAI221_X1 _11200_ (.A(_02186_),
    .B1(_02028_),
    .B2(_02026_),
    .C1(_02020_),
    .C2(_02021_),
    .ZN(_02187_));
 AOI21_X1 _11201_ (.A(_02183_),
    .B1(_02094_),
    .B2(_02187_),
    .ZN(_02188_));
 NOR2_X1 _11202_ (.A1(_01886_),
    .A2(_01912_),
    .ZN(_02189_));
 NOR2_X1 _11203_ (.A1(_02093_),
    .A2(_02189_),
    .ZN(_02190_));
 MUX2_X1 _11204_ (.A(_02190_),
    .B(_02093_),
    .S(_02006_),
    .Z(_02191_));
 MUX2_X2 _11205_ (.A(_02188_),
    .B(_02183_),
    .S(_02191_),
    .Z(_02192_));
 NOR4_X4 _11206_ (.A1(_02180_),
    .A2(_02122_),
    .A3(_02182_),
    .A4(_02192_),
    .ZN(_02193_));
 OAI221_X2 _11207_ (.A(_01912_),
    .B1(_02006_),
    .B2(_02093_),
    .C1(_02183_),
    .C2(_02191_),
    .ZN(_02194_));
 OR2_X1 _11208_ (.A1(_02193_),
    .A2(_02194_),
    .ZN(_02195_));
 BUF_X4 _11209_ (.A(_02195_),
    .Z(_02196_));
 XOR2_X2 _11210_ (.A(_02175_),
    .B(_02179_),
    .Z(_02197_));
 NAND2_X2 _11211_ (.A1(_02047_),
    .A2(_02019_),
    .ZN(_02198_));
 NOR2_X1 _11212_ (.A1(_02048_),
    .A2(_02198_),
    .ZN(_02199_));
 NOR4_X4 _11213_ (.A1(_01989_),
    .A2(_02036_),
    .A3(_02053_),
    .A4(_02199_),
    .ZN(_02200_));
 AOI21_X1 _11214_ (.A(_01990_),
    .B1(_02019_),
    .B2(_02047_),
    .ZN(_02201_));
 OAI21_X2 _11215_ (.A(_02201_),
    .B1(_02035_),
    .B2(_02029_),
    .ZN(_02202_));
 INV_X2 _11216_ (.A(_02048_),
    .ZN(_02203_));
 NAND2_X1 _11217_ (.A1(_02203_),
    .A2(_01990_),
    .ZN(_02204_));
 NOR2_X1 _11218_ (.A1(_02198_),
    .A2(_02204_),
    .ZN(_02205_));
 AOI21_X2 _11219_ (.A(_02205_),
    .B1(_02177_),
    .B2(_02048_),
    .ZN(_02206_));
 OR2_X4 _11220_ (.A1(_02029_),
    .A2(_02035_),
    .ZN(_02207_));
 OAI211_X4 _11221_ (.A(_02202_),
    .B(_02206_),
    .C1(_02204_),
    .C2(_02207_),
    .ZN(_02208_));
 AND4_X2 _11222_ (.A1(_02200_),
    .A2(_02208_),
    .A3(_02126_),
    .A4(_02121_),
    .ZN(_02209_));
 AOI21_X4 _11223_ (.A(_02054_),
    .B1(_02126_),
    .B2(_02121_),
    .ZN(_02210_));
 OAI21_X4 _11224_ (.A(_02198_),
    .B1(_02035_),
    .B2(_02029_),
    .ZN(_02211_));
 OR3_X1 _11225_ (.A1(_01989_),
    .A2(_02046_),
    .A3(_02052_),
    .ZN(_02212_));
 AOI22_X4 _11226_ (.A1(_02203_),
    .A2(_02211_),
    .B1(_02212_),
    .B2(_02207_),
    .ZN(_02213_));
 AND3_X1 _11227_ (.A1(_02177_),
    .A2(_02126_),
    .A3(_02213_),
    .ZN(_02214_));
 OAI22_X4 _11228_ (.A1(_02197_),
    .A2(_02209_),
    .B1(_02210_),
    .B2(_02214_),
    .ZN(_02215_));
 AND3_X1 _11229_ (.A1(_02208_),
    .A2(_02156_),
    .A3(net15),
    .ZN(_02216_));
 AOI221_X2 _11230_ (.A(_02176_),
    .B1(_02166_),
    .B2(_02165_),
    .C1(_02159_),
    .C2(_01960_),
    .ZN(_02217_));
 NOR4_X2 _11231_ (.A1(_02022_),
    .A2(_02036_),
    .A3(_02053_),
    .A4(_02164_),
    .ZN(_02218_));
 AOI21_X2 _11232_ (.A(_02192_),
    .B1(_02217_),
    .B2(_02218_),
    .ZN(_02219_));
 NAND3_X1 _11233_ (.A1(_02084_),
    .A2(_02065_),
    .A3(_02069_),
    .ZN(_02220_));
 INV_X1 _11234_ (.A(_02080_),
    .ZN(_02221_));
 NAND2_X1 _11235_ (.A1(_01122_),
    .A2(_02159_),
    .ZN(_02222_));
 NAND2_X1 _11236_ (.A1(_01089_),
    .A2(_02168_),
    .ZN(_02223_));
 AOI221_X2 _11237_ (.A(_02192_),
    .B1(_02220_),
    .B2(_02221_),
    .C1(_02222_),
    .C2(_02223_),
    .ZN(_02224_));
 NOR3_X4 _11238_ (.A1(_02216_),
    .A2(_02219_),
    .A3(_02224_),
    .ZN(_02225_));
 NAND3_X2 _11239_ (.A1(_02208_),
    .A2(_02156_),
    .A3(_02127_),
    .ZN(_02226_));
 AND2_X1 _11240_ (.A1(_02218_),
    .A2(_02217_),
    .ZN(_02227_));
 XNOR2_X1 _11241_ (.A(_01122_),
    .B(_02159_),
    .ZN(_02228_));
 AND3_X1 _11242_ (.A1(_02084_),
    .A2(_02065_),
    .A3(_02069_),
    .ZN(_02229_));
 OAI21_X2 _11243_ (.A(_02228_),
    .B1(_02229_),
    .B2(_02080_),
    .ZN(_02230_));
 NAND4_X4 _11244_ (.A1(_02192_),
    .A2(_02226_),
    .A3(_02227_),
    .A4(_02230_),
    .ZN(_02231_));
 AOI21_X4 _11245_ (.A(_02215_),
    .B1(_02225_),
    .B2(_02231_),
    .ZN(_02232_));
 AOI21_X4 _11246_ (.A(_02174_),
    .B1(_02196_),
    .B2(_02232_),
    .ZN(_02233_));
 XNOR2_X2 _11247_ (.A(_02164_),
    .B(_02154_),
    .ZN(_02234_));
 NOR4_X4 _11248_ (.A1(_02054_),
    .A2(_02092_),
    .A3(_02121_),
    .A4(_08963_),
    .ZN(_02235_));
 INV_X2 _11249_ (.A(_01708_),
    .ZN(_02236_));
 AOI221_X2 _11250_ (.A(_02235_),
    .B1(_02236_),
    .B2(_02132_),
    .C1(_01136_),
    .C2(_01116_),
    .ZN(_02237_));
 MUX2_X2 _11251_ (.A(_02131_),
    .B(_02129_),
    .S(_02122_),
    .Z(_02238_));
 NAND2_X1 _11252_ (.A1(_02159_),
    .A2(_02160_),
    .ZN(_02239_));
 NAND2_X1 _11253_ (.A1(_02167_),
    .A2(_02170_),
    .ZN(_02240_));
 NAND2_X1 _11254_ (.A1(_02124_),
    .A2(_02127_),
    .ZN(_02241_));
 OR2_X1 _11255_ (.A1(_02159_),
    .A2(_02160_),
    .ZN(_02242_));
 OAI221_X2 _11256_ (.A(_02239_),
    .B1(_02240_),
    .B2(_02241_),
    .C1(_02122_),
    .C2(_02242_),
    .ZN(_02243_));
 BUF_X4 _11257_ (.A(_02243_),
    .Z(_02244_));
 OR2_X1 _11258_ (.A1(_02065_),
    .A2(_02156_),
    .ZN(_02245_));
 AND4_X1 _11259_ (.A1(_02200_),
    .A2(_02208_),
    .A3(_02069_),
    .A4(net15),
    .ZN(_02246_));
 NAND2_X1 _11260_ (.A1(_02065_),
    .A2(_02156_),
    .ZN(_02247_));
 OAI21_X2 _11261_ (.A(_02245_),
    .B1(_02246_),
    .B2(_02247_),
    .ZN(_02248_));
 NOR4_X4 _11262_ (.A1(_02237_),
    .A2(_02238_),
    .A3(_02244_),
    .A4(_02248_),
    .ZN(_02249_));
 NOR3_X2 _11263_ (.A1(_02122_),
    .A2(_02234_),
    .A3(_02249_),
    .ZN(_02250_));
 NAND3_X1 _11264_ (.A1(_02123_),
    .A2(_02133_),
    .A3(_02173_),
    .ZN(_02251_));
 AND2_X1 _11265_ (.A1(_02251_),
    .A2(_02248_),
    .ZN(_02252_));
 XNOR2_X2 _11266_ (.A(_02138_),
    .B(_02156_),
    .ZN(_02253_));
 AOI21_X4 _11267_ (.A(_02122_),
    .B1(_02234_),
    .B2(_02253_),
    .ZN(_02254_));
 AND2_X1 _11268_ (.A1(_02254_),
    .A2(_02249_),
    .ZN(_02255_));
 NOR4_X4 _11269_ (.A1(_02233_),
    .A2(_02250_),
    .A3(_02252_),
    .A4(_02255_),
    .ZN(_02256_));
 NAND2_X2 _11270_ (.A1(_02126_),
    .A2(_02241_),
    .ZN(_02257_));
 OAI22_X4 _11271_ (.A1(_02200_),
    .A2(_02126_),
    .B1(_02213_),
    .B2(_02257_),
    .ZN(_02258_));
 NOR4_X4 _11272_ (.A1(_02237_),
    .A2(_02238_),
    .A3(_02254_),
    .A4(_02244_),
    .ZN(_02259_));
 AND2_X1 _11273_ (.A1(_02200_),
    .A2(_02126_),
    .ZN(_02260_));
 NOR2_X1 _11274_ (.A1(_02208_),
    .A2(_02260_),
    .ZN(_02261_));
 NOR2_X1 _11275_ (.A1(_02209_),
    .A2(_02261_),
    .ZN(_02262_));
 NOR2_X1 _11276_ (.A1(_02259_),
    .A2(_02262_),
    .ZN(_02263_));
 NOR2_X4 _11277_ (.A1(_02258_),
    .A2(_02263_),
    .ZN(_02264_));
 AND2_X2 _11278_ (.A1(_02256_),
    .A2(_02264_),
    .ZN(_02265_));
 NOR2_X4 _11279_ (.A1(_02193_),
    .A2(_02194_),
    .ZN(_02266_));
 OR3_X2 _11280_ (.A1(_02216_),
    .A2(_02219_),
    .A3(_02224_),
    .ZN(_02267_));
 AND4_X2 _11281_ (.A1(_02192_),
    .A2(_02226_),
    .A3(_02227_),
    .A4(_02230_),
    .ZN(_02268_));
 NOR2_X4 _11282_ (.A1(_02267_),
    .A2(_02268_),
    .ZN(_02269_));
 NAND4_X2 _11283_ (.A1(_02200_),
    .A2(_02208_),
    .A3(_02126_),
    .A4(_02121_),
    .ZN(_02270_));
 OAI21_X2 _11284_ (.A(_02124_),
    .B1(_02092_),
    .B2(net15),
    .ZN(_02271_));
 NAND3_X2 _11285_ (.A1(_02177_),
    .A2(_02126_),
    .A3(_02213_),
    .ZN(_02272_));
 AOI22_X4 _11286_ (.A1(_02180_),
    .A2(_02270_),
    .B1(_02271_),
    .B2(_02272_),
    .ZN(_02273_));
 NAND2_X2 _11287_ (.A1(_02259_),
    .A2(_02273_),
    .ZN(_02274_));
 AOI21_X4 _11288_ (.A(_02266_),
    .B1(_02269_),
    .B2(_02274_),
    .ZN(_02275_));
 XNOR2_X2 _11289_ (.A(_02180_),
    .B(_02209_),
    .ZN(_02276_));
 INV_X1 _11290_ (.A(_02276_),
    .ZN(_02277_));
 NAND3_X4 _11291_ (.A1(_02259_),
    .A2(_02196_),
    .A3(_02232_),
    .ZN(_02278_));
 AOI21_X4 _11292_ (.A(_02235_),
    .B1(_02236_),
    .B2(net7),
    .ZN(_02279_));
 NOR2_X1 _11293_ (.A1(_08999_),
    .A2(_01134_),
    .ZN(_02280_));
 NAND2_X1 _11294_ (.A1(_01122_),
    .A2(_02280_),
    .ZN(_02281_));
 OAI21_X1 _11295_ (.A(_02128_),
    .B1(_02173_),
    .B2(_02281_),
    .ZN(_02282_));
 NOR2_X1 _11296_ (.A1(_02279_),
    .A2(_02282_),
    .ZN(_02283_));
 AOI21_X1 _11297_ (.A(_02279_),
    .B1(_02244_),
    .B2(_01090_),
    .ZN(_02284_));
 OAI22_X1 _11298_ (.A1(_01135_),
    .A2(_02279_),
    .B1(_02244_),
    .B2(_01136_),
    .ZN(_02285_));
 NOR2_X1 _11299_ (.A1(_02284_),
    .A2(_02285_),
    .ZN(_02286_));
 XNOR2_X1 _11300_ (.A(_01960_),
    .B(_02244_),
    .ZN(_02287_));
 OR3_X1 _11301_ (.A1(_01122_),
    .A2(_01135_),
    .A3(_02287_),
    .ZN(_02288_));
 AOI221_X2 _11302_ (.A(_02277_),
    .B1(_02278_),
    .B2(_02283_),
    .C1(_02286_),
    .C2(_02288_),
    .ZN(_02289_));
 BUF_X4 _11303_ (.A(_02289_),
    .Z(_02290_));
 NOR2_X1 _11304_ (.A1(_08868_),
    .A2(_01649_),
    .ZN(_08887_));
 NAND3_X1 _11305_ (.A1(_01716_),
    .A2(_01599_),
    .A3(_01715_),
    .ZN(_02291_));
 AND2_X1 _11306_ (.A1(_01743_),
    .A2(_02291_),
    .ZN(_02292_));
 MUX2_X1 _11307_ (.A(_08887_),
    .B(_02292_),
    .S(_01721_),
    .Z(_08902_));
 AOI21_X1 _11308_ (.A(_08906_),
    .B1(_01723_),
    .B2(_08907_),
    .ZN(_02293_));
 XNOR2_X1 _11309_ (.A(_08904_),
    .B(_02293_),
    .ZN(_02294_));
 MUX2_X1 _11310_ (.A(_08902_),
    .B(_02294_),
    .S(_01819_),
    .Z(_08931_));
 OR3_X1 _11311_ (.A1(_08933_),
    .A2(_08935_),
    .A3(_01824_),
    .ZN(_02295_));
 AND2_X1 _11312_ (.A1(_01825_),
    .A2(_02295_),
    .ZN(_02296_));
 MUX2_X1 _11313_ (.A(_08931_),
    .B(_02296_),
    .S(_01916_),
    .Z(_08949_));
 XOR2_X1 _11314_ (.A(_01926_),
    .B(_01925_),
    .Z(_02297_));
 MUX2_X1 _11315_ (.A(_08949_),
    .B(_02297_),
    .S(_02017_),
    .Z(_08966_));
 XNOR2_X1 _11316_ (.A(_01705_),
    .B(_02146_),
    .ZN(_02298_));
 MUX2_X1 _11317_ (.A(_08966_),
    .B(_02298_),
    .S(_02132_),
    .Z(_02299_));
 CLKBUF_X3 _11318_ (.A(_02299_),
    .Z(_08998_));
 AND2_X1 _11319_ (.A1(_01960_),
    .A2(_08998_),
    .ZN(_02300_));
 INV_X2 _11320_ (.A(_09011_),
    .ZN(_02301_));
 INV_X1 _11321_ (.A(_09012_),
    .ZN(_02302_));
 INV_X1 _11322_ (.A(_09017_),
    .ZN(_02303_));
 INV_X1 _11323_ (.A(_09023_),
    .ZN(_02304_));
 INV_X1 _11324_ (.A(_09008_),
    .ZN(_02305_));
 AOI21_X4 _11325_ (.A(_01883_),
    .B1(net9),
    .B2(_01310_),
    .ZN(_02306_));
 INV_X4 _11326_ (.A(_02306_),
    .ZN(_08940_));
 NOR2_X1 _11327_ (.A1(_01696_),
    .A2(_01843_),
    .ZN(_02307_));
 OAI21_X2 _11328_ (.A(_01523_),
    .B1(_01881_),
    .B2(net11),
    .ZN(_08890_));
 OR2_X1 _11329_ (.A1(_02307_),
    .A2(_08890_),
    .ZN(_02308_));
 NOR3_X2 _11330_ (.A1(_02103_),
    .A2(_08940_),
    .A3(_02308_),
    .ZN(_02309_));
 BUF_X1 _11331_ (.A(_09009_),
    .Z(_02310_));
 INV_X1 _11332_ (.A(_02310_),
    .ZN(_02311_));
 OAI21_X1 _11333_ (.A(_02305_),
    .B1(_02309_),
    .B2(_02311_),
    .ZN(_02312_));
 AOI21_X1 _11334_ (.A(_09005_),
    .B1(_02312_),
    .B2(_09006_),
    .ZN(_02313_));
 INV_X2 _11335_ (.A(_09024_),
    .ZN(_02314_));
 OAI21_X4 _11336_ (.A(_02304_),
    .B1(_02314_),
    .B2(_02313_),
    .ZN(_02315_));
 BUF_X1 _11337_ (.A(_09021_),
    .Z(_02316_));
 AOI21_X4 _11338_ (.A(_09020_),
    .B1(_02315_),
    .B2(_02316_),
    .ZN(_02317_));
 BUF_X1 _11339_ (.A(_09018_),
    .Z(_02318_));
 INV_X1 _11340_ (.A(_02318_),
    .ZN(_02319_));
 OAI21_X4 _11341_ (.A(_02303_),
    .B1(_02319_),
    .B2(_02317_),
    .ZN(_02320_));
 BUF_X1 _11342_ (.A(_09015_),
    .Z(_02321_));
 AOI21_X4 _11343_ (.A(_09014_),
    .B1(_02320_),
    .B2(_02321_),
    .ZN(_02322_));
 OR2_X4 _11344_ (.A1(_02302_),
    .A2(_02322_),
    .ZN(_02323_));
 NAND2_X1 _11345_ (.A1(_02301_),
    .A2(_02323_),
    .ZN(_02324_));
 XNOR2_X1 _11346_ (.A(_01122_),
    .B(_08998_),
    .ZN(_02325_));
 AOI21_X1 _11347_ (.A(_02300_),
    .B1(_02325_),
    .B2(_02324_),
    .ZN(_02326_));
 XNOR2_X2 _11348_ (.A(_09000_),
    .B(_01133_),
    .ZN(_02327_));
 NOR2_X2 _11349_ (.A1(_01117_),
    .A2(_02327_),
    .ZN(_02328_));
 NAND2_X1 _11350_ (.A1(_01089_),
    .A2(_02327_),
    .ZN(_02329_));
 XOR2_X2 _11351_ (.A(_09000_),
    .B(_01133_),
    .Z(_02330_));
 NAND2_X1 _11352_ (.A1(_01122_),
    .A2(_02330_),
    .ZN(_02331_));
 AOI22_X4 _11353_ (.A1(_02323_),
    .A2(_02301_),
    .B1(_02329_),
    .B2(_02331_),
    .ZN(_02332_));
 NOR2_X1 _11354_ (.A1(_02332_),
    .A2(_02328_),
    .ZN(_02333_));
 MUX2_X1 _11355_ (.A(_02326_),
    .B(_02333_),
    .S(_02278_),
    .Z(_02334_));
 BUF_X4 _11356_ (.A(_02334_),
    .Z(_02335_));
 AND3_X4 _11357_ (.A1(_02275_),
    .A2(_02290_),
    .A3(_02335_),
    .ZN(_02336_));
 XNOR2_X1 _11358_ (.A(_01597_),
    .B(_01310_),
    .ZN(_02337_));
 MUX2_X1 _11359_ (.A(_08890_),
    .B(_02337_),
    .S(_01721_),
    .Z(_08905_));
 AOI21_X1 _11360_ (.A(_08914_),
    .B1(_01882_),
    .B2(_08915_),
    .ZN(_02338_));
 XNOR2_X1 _11361_ (.A(_08907_),
    .B(_02338_),
    .ZN(_02339_));
 MUX2_X1 _11362_ (.A(_08905_),
    .B(_02339_),
    .S(_01819_),
    .Z(_08934_));
 XOR2_X1 _11363_ (.A(_08936_),
    .B(_01823_),
    .Z(_02340_));
 MUX2_X1 _11364_ (.A(_08934_),
    .B(_02340_),
    .S(_01916_),
    .Z(_08952_));
 OR3_X1 _11365_ (.A1(_08954_),
    .A2(_08956_),
    .A3(_01923_),
    .ZN(_02341_));
 AND2_X1 _11366_ (.A1(_01924_),
    .A2(_02341_),
    .ZN(_02342_));
 MUX2_X1 _11367_ (.A(_08952_),
    .B(_02342_),
    .S(_02017_),
    .Z(_08969_));
 XNOR2_X1 _11368_ (.A(_02105_),
    .B(_01703_),
    .ZN(_02343_));
 BUF_X8 _11369_ (.A(_02132_),
    .Z(_02344_));
 MUX2_X2 _11370_ (.A(_08969_),
    .B(_02343_),
    .S(_02344_),
    .Z(_09001_));
 AND4_X2 _11371_ (.A1(_02259_),
    .A2(_02196_),
    .A3(_02232_),
    .A4(_09001_),
    .ZN(_02345_));
 XNOR2_X2 _11372_ (.A(_09003_),
    .B(_01131_),
    .ZN(_02346_));
 BUF_X8 _11373_ (.A(_02278_),
    .Z(_02347_));
 AOI21_X4 _11374_ (.A(_02345_),
    .B1(_02346_),
    .B2(_02347_),
    .ZN(_02348_));
 INV_X1 _11375_ (.A(_02348_),
    .ZN(_09010_));
 NAND3_X1 _11376_ (.A1(_02265_),
    .A2(_02336_),
    .A3(_09010_),
    .ZN(_02349_));
 XNOR2_X2 _11377_ (.A(_02302_),
    .B(_02322_),
    .ZN(_02350_));
 NAND2_X4 _11378_ (.A1(_02256_),
    .A2(_02264_),
    .ZN(_02351_));
 NAND3_X4 _11379_ (.A1(_02275_),
    .A2(_02290_),
    .A3(_02335_),
    .ZN(_02352_));
 NOR2_X4 _11380_ (.A1(_02351_),
    .A2(_02352_),
    .ZN(_02353_));
 OAI21_X4 _11381_ (.A(_02349_),
    .B1(_02350_),
    .B2(_02353_),
    .ZN(_02354_));
 CLKBUF_X3 _11382_ (.A(_01122_),
    .Z(_02355_));
 CLKBUF_X3 _11383_ (.A(_02355_),
    .Z(_02356_));
 INV_X1 _11384_ (.A(_09037_),
    .ZN(_02357_));
 INV_X1 _11385_ (.A(_09043_),
    .ZN(_02358_));
 INV_X1 _11386_ (.A(_09031_),
    .ZN(_02359_));
 OAI21_X2 _11387_ (.A(_09032_),
    .B1(_09025_),
    .B2(_09026_),
    .ZN(_02360_));
 NAND2_X2 _11388_ (.A1(_02360_),
    .A2(_02359_),
    .ZN(_02361_));
 AND2_X4 _11389_ (.A1(_09029_),
    .A2(_02361_),
    .ZN(_02362_));
 OAI21_X4 _11390_ (.A(_09044_),
    .B1(_02362_),
    .B2(_09028_),
    .ZN(_02363_));
 NAND2_X4 _11391_ (.A1(_02358_),
    .A2(_02363_),
    .ZN(_02364_));
 AOI21_X4 _11392_ (.A(_09040_),
    .B1(_02364_),
    .B2(_09041_),
    .ZN(_02365_));
 INV_X1 _11393_ (.A(_09038_),
    .ZN(_02366_));
 OAI21_X4 _11394_ (.A(_02357_),
    .B1(_02366_),
    .B2(_02365_),
    .ZN(_02367_));
 AND2_X4 _11395_ (.A1(_09035_),
    .A2(_02367_),
    .ZN(_02368_));
 NOR2_X4 _11396_ (.A1(_02368_),
    .A2(_09034_),
    .ZN(_02369_));
 XNOR2_X2 _11397_ (.A(_02356_),
    .B(_02369_),
    .ZN(_02370_));
 OAI21_X4 _11398_ (.A(_02273_),
    .B1(_02267_),
    .B2(_02268_),
    .ZN(_02371_));
 OAI221_X2 _11399_ (.A(_02259_),
    .B1(_02266_),
    .B2(_02371_),
    .C1(_02214_),
    .C2(_02210_),
    .ZN(_02372_));
 XNOR2_X2 _11400_ (.A(_02276_),
    .B(_02372_),
    .ZN(_02373_));
 NOR3_X4 _11401_ (.A1(_02174_),
    .A2(_02266_),
    .A3(_02371_),
    .ZN(_02374_));
 NOR2_X2 _11402_ (.A1(_02279_),
    .A2(_02300_),
    .ZN(_02375_));
 INV_X1 _11403_ (.A(_08963_),
    .ZN(_02376_));
 MUX2_X2 _11404_ (.A(_02376_),
    .B(_02236_),
    .S(net7),
    .Z(_02377_));
 XNOR2_X1 _11405_ (.A(_01089_),
    .B(_02280_),
    .ZN(_02378_));
 XNOR2_X1 _11406_ (.A(_02377_),
    .B(_02378_),
    .ZN(_02379_));
 NOR2_X2 _11407_ (.A1(_02328_),
    .A2(_02379_),
    .ZN(_02380_));
 NOR3_X4 _11408_ (.A1(_02237_),
    .A2(_02238_),
    .A3(_02244_),
    .ZN(_02381_));
 AOI21_X4 _11409_ (.A(_02173_),
    .B1(_02133_),
    .B2(_02123_),
    .ZN(_02382_));
 NOR2_X2 _11410_ (.A1(_02381_),
    .A2(_02382_),
    .ZN(_02383_));
 AOI22_X4 _11411_ (.A1(_02374_),
    .A2(_02375_),
    .B1(_02380_),
    .B2(_02383_),
    .ZN(_02384_));
 INV_X1 _11412_ (.A(_02384_),
    .ZN(_02385_));
 OAI33_X1 _11413_ (.A1(_02174_),
    .A2(_02266_),
    .A3(_02371_),
    .B1(_02248_),
    .B2(_02382_),
    .B3(_02381_),
    .ZN(_02386_));
 INV_X1 _11414_ (.A(_02321_),
    .ZN(_02387_));
 INV_X1 _11415_ (.A(_09020_),
    .ZN(_02388_));
 INV_X1 _11416_ (.A(_09005_),
    .ZN(_02389_));
 OAI21_X1 _11417_ (.A(_09006_),
    .B1(_02310_),
    .B2(_09008_),
    .ZN(_02390_));
 AOI21_X1 _11418_ (.A(_02314_),
    .B1(_02389_),
    .B2(_02390_),
    .ZN(_02391_));
 NOR2_X1 _11419_ (.A1(_09023_),
    .A2(_02391_),
    .ZN(_02392_));
 INV_X1 _11420_ (.A(_02316_),
    .ZN(_02393_));
 OAI21_X1 _11421_ (.A(_02388_),
    .B1(_02392_),
    .B2(_02393_),
    .ZN(_02394_));
 AOI21_X2 _11422_ (.A(_09017_),
    .B1(_02394_),
    .B2(_02318_),
    .ZN(_02395_));
 NOR2_X1 _11423_ (.A1(_02387_),
    .A2(_02395_),
    .ZN(_02396_));
 OAI21_X1 _11424_ (.A(_09012_),
    .B1(_09014_),
    .B2(_02396_),
    .ZN(_02397_));
 AND2_X2 _11425_ (.A1(_02301_),
    .A2(_02397_),
    .ZN(_02398_));
 NOR2_X2 _11426_ (.A1(_01090_),
    .A2(_02398_),
    .ZN(_02399_));
 NAND2_X1 _11427_ (.A1(_02386_),
    .A2(_02399_),
    .ZN(_02400_));
 NOR2_X1 _11428_ (.A1(_02355_),
    .A2(_02398_),
    .ZN(_02401_));
 NAND2_X1 _11429_ (.A1(_02386_),
    .A2(_02401_),
    .ZN(_02402_));
 INV_X1 _11430_ (.A(_08998_),
    .ZN(_02403_));
 MUX2_X1 _11431_ (.A(_02403_),
    .B(_02327_),
    .S(net2),
    .Z(_02404_));
 CLKBUF_X3 _11432_ (.A(_02404_),
    .Z(_02405_));
 MUX2_X1 _11433_ (.A(_02400_),
    .B(_02402_),
    .S(_02405_),
    .Z(_02406_));
 NAND4_X2 _11434_ (.A1(_02265_),
    .A2(_02385_),
    .A3(_02352_),
    .A4(_02406_),
    .ZN(_02407_));
 XOR2_X2 _11435_ (.A(_02373_),
    .B(_02407_),
    .Z(_02408_));
 NOR3_X2 _11436_ (.A1(_02174_),
    .A2(_02215_),
    .A3(_02269_),
    .ZN(_02409_));
 NOR2_X4 _11437_ (.A1(_02196_),
    .A2(_02409_),
    .ZN(_02410_));
 OR2_X1 _11438_ (.A1(_02279_),
    .A2(_02300_),
    .ZN(_02411_));
 OR2_X1 _11439_ (.A1(_02328_),
    .A2(_02379_),
    .ZN(_02412_));
 MUX2_X1 _11440_ (.A(_02411_),
    .B(_02412_),
    .S(_02278_),
    .Z(_02413_));
 NAND2_X2 _11441_ (.A1(_02301_),
    .A2(_02397_),
    .ZN(_02414_));
 NAND3_X1 _11442_ (.A1(_01090_),
    .A2(_02327_),
    .A3(_02414_),
    .ZN(_02415_));
 NAND3_X1 _11443_ (.A1(_02355_),
    .A2(_02330_),
    .A3(_02414_),
    .ZN(_02416_));
 AOI21_X1 _11444_ (.A(_02374_),
    .B1(_02415_),
    .B2(_02416_),
    .ZN(_02417_));
 NAND2_X1 _11445_ (.A1(_08998_),
    .A2(_02399_),
    .ZN(_02418_));
 NAND2_X1 _11446_ (.A1(_02403_),
    .A2(_02401_),
    .ZN(_02419_));
 AOI21_X1 _11447_ (.A(net2),
    .B1(_02418_),
    .B2(_02419_),
    .ZN(_02420_));
 OR3_X2 _11448_ (.A1(_02413_),
    .A2(_02417_),
    .A3(_02420_),
    .ZN(_02421_));
 NAND3_X1 _11449_ (.A1(_02158_),
    .A2(_02196_),
    .A3(_02273_),
    .ZN(_02422_));
 AOI221_X2 _11450_ (.A(_02382_),
    .B1(_02422_),
    .B2(_02381_),
    .C1(_02225_),
    .C2(_02231_),
    .ZN(_02423_));
 NAND4_X2 _11451_ (.A1(_02373_),
    .A2(_02256_),
    .A3(_02264_),
    .A4(_02423_),
    .ZN(_02424_));
 OAI21_X4 _11452_ (.A(_02410_),
    .B1(_02421_),
    .B2(_02424_),
    .ZN(_02425_));
 NOR4_X2 _11453_ (.A1(_02174_),
    .A2(_02196_),
    .A3(_02215_),
    .A4(_02269_),
    .ZN(_02426_));
 AOI21_X4 _11454_ (.A(_02426_),
    .B1(_02274_),
    .B2(_02269_),
    .ZN(_02427_));
 INV_X1 _11455_ (.A(_02427_),
    .ZN(_02428_));
 NAND2_X1 _11456_ (.A1(_02290_),
    .A2(net19),
    .ZN(_02429_));
 OAI21_X2 _11457_ (.A(_02428_),
    .B1(_02429_),
    .B2(_02351_),
    .ZN(_02430_));
 NOR2_X1 _11458_ (.A1(_01097_),
    .A2(_02104_),
    .ZN(_02431_));
 AOI21_X1 _11459_ (.A(_02112_),
    .B1(net7),
    .B2(_01150_),
    .ZN(_02432_));
 INV_X1 _11460_ (.A(_02112_),
    .ZN(_02433_));
 NOR3_X4 _11461_ (.A1(_01929_),
    .A2(_02433_),
    .A3(_02122_),
    .ZN(_02434_));
 OAI21_X2 _11462_ (.A(_02431_),
    .B1(_02432_),
    .B2(_02434_),
    .ZN(_02435_));
 AND4_X1 _11463_ (.A1(_09006_),
    .A2(_02310_),
    .A3(_09012_),
    .A4(_09024_),
    .ZN(_02436_));
 NAND4_X1 _11464_ (.A1(_02321_),
    .A2(_02318_),
    .A3(_02316_),
    .A4(_02436_),
    .ZN(_02437_));
 OR4_X2 _11465_ (.A1(_08940_),
    .A2(_02308_),
    .A3(_02435_),
    .A4(_02437_),
    .ZN(_02438_));
 NOR2_X2 _11466_ (.A1(_02266_),
    .A2(_02371_),
    .ZN(_02439_));
 AOI221_X2 _11467_ (.A(_02438_),
    .B1(_02331_),
    .B2(_02329_),
    .C1(_02259_),
    .C2(_02439_),
    .ZN(_02440_));
 NAND2_X1 _11468_ (.A1(_01090_),
    .A2(_02403_),
    .ZN(_02441_));
 NAND2_X1 _11469_ (.A1(_01122_),
    .A2(_08998_),
    .ZN(_02442_));
 AOI211_X2 _11470_ (.A(net2),
    .B(_02438_),
    .C1(_02441_),
    .C2(_02442_),
    .ZN(_02443_));
 OR3_X1 _11471_ (.A1(_02410_),
    .A2(_02440_),
    .A3(_02443_),
    .ZN(_02444_));
 BUF_X4 _11472_ (.A(_02444_),
    .Z(_02445_));
 AND4_X2 _11473_ (.A1(_02256_),
    .A2(_02264_),
    .A3(_02427_),
    .A4(_02290_),
    .ZN(_02446_));
 NAND3_X2 _11474_ (.A1(_02335_),
    .A2(_02445_),
    .A3(_02446_),
    .ZN(_02447_));
 NAND3_X4 _11475_ (.A1(_02425_),
    .A2(_02430_),
    .A3(_02447_),
    .ZN(_02448_));
 NOR2_X1 _11476_ (.A1(_02174_),
    .A2(_02258_),
    .ZN(_02449_));
 NOR2_X1 _11477_ (.A1(_02262_),
    .A2(_02449_),
    .ZN(_02450_));
 NOR3_X4 _11478_ (.A1(_02410_),
    .A2(_02440_),
    .A3(_02443_),
    .ZN(_02451_));
 AND3_X1 _11479_ (.A1(_02256_),
    .A2(_02427_),
    .A3(_02290_),
    .ZN(_02452_));
 AOI21_X1 _11480_ (.A(_02450_),
    .B1(_02451_),
    .B2(_02452_),
    .ZN(_02453_));
 OAI21_X1 _11481_ (.A(_02372_),
    .B1(_02262_),
    .B2(_02449_),
    .ZN(_02454_));
 AND2_X1 _11482_ (.A1(_02301_),
    .A2(_02323_),
    .ZN(_02455_));
 XNOR2_X1 _11483_ (.A(_01090_),
    .B(_08998_),
    .ZN(_02456_));
 OAI22_X1 _11484_ (.A1(_01117_),
    .A2(_02403_),
    .B1(_02455_),
    .B2(_02456_),
    .ZN(_02457_));
 OR2_X1 _11485_ (.A1(_02328_),
    .A2(_02332_),
    .ZN(_02458_));
 MUX2_X2 _11486_ (.A(_02457_),
    .B(_02458_),
    .S(_02278_),
    .Z(_02459_));
 NOR3_X2 _11487_ (.A1(_02279_),
    .A2(_02238_),
    .A3(_02244_),
    .ZN(_02460_));
 NAND2_X1 _11488_ (.A1(_01135_),
    .A2(_02173_),
    .ZN(_02461_));
 NAND2_X1 _11489_ (.A1(_02377_),
    .A2(_02244_),
    .ZN(_02462_));
 OAI221_X2 _11490_ (.A(_02355_),
    .B1(_02377_),
    .B2(_02461_),
    .C1(_02462_),
    .C2(_01135_),
    .ZN(_02463_));
 NAND2_X1 _11491_ (.A1(_02280_),
    .A2(_02279_),
    .ZN(_02464_));
 OAI221_X2 _11492_ (.A(_01090_),
    .B1(_02279_),
    .B2(_02461_),
    .C1(_02464_),
    .C2(_02287_),
    .ZN(_02465_));
 AOI22_X4 _11493_ (.A1(_02439_),
    .A2(_02460_),
    .B1(_02463_),
    .B2(_02465_),
    .ZN(_02466_));
 NOR3_X4 _11494_ (.A1(_02254_),
    .A2(_02459_),
    .A3(_02466_),
    .ZN(_02467_));
 NOR2_X2 _11495_ (.A1(_02036_),
    .A2(_02053_),
    .ZN(_02468_));
 MUX2_X2 _11496_ (.A(_02126_),
    .B(_02257_),
    .S(_02468_),
    .Z(_02469_));
 XOR2_X2 _11497_ (.A(_02233_),
    .B(_02469_),
    .Z(_02470_));
 AOI22_X4 _11498_ (.A1(_01989_),
    .A2(_02207_),
    .B1(_02211_),
    .B2(_02203_),
    .ZN(_02471_));
 AOI21_X2 _11499_ (.A(_02471_),
    .B1(_02181_),
    .B2(_02468_),
    .ZN(_02472_));
 NAND3_X2 _11500_ (.A1(_02208_),
    .A2(net15),
    .A3(_02471_),
    .ZN(_02473_));
 AOI21_X4 _11501_ (.A(_02472_),
    .B1(_02473_),
    .B2(_02260_),
    .ZN(_02474_));
 NAND3_X1 _11502_ (.A1(_02467_),
    .A2(_02470_),
    .A3(_02474_),
    .ZN(_02475_));
 MUX2_X1 _11503_ (.A(_02453_),
    .B(_02454_),
    .S(_02475_),
    .Z(_02476_));
 BUF_X4 _11504_ (.A(_02476_),
    .Z(_02477_));
 MUX2_X2 _11505_ (.A(_08998_),
    .B(_02330_),
    .S(net2),
    .Z(_02478_));
 NOR2_X1 _11506_ (.A1(_02355_),
    .A2(_02414_),
    .ZN(_02479_));
 OAI22_X4 _11507_ (.A1(_02351_),
    .A2(_02352_),
    .B1(_02399_),
    .B2(_02479_),
    .ZN(_02480_));
 XNOR2_X2 _11508_ (.A(_02478_),
    .B(_02480_),
    .ZN(_02481_));
 NOR4_X2 _11509_ (.A1(_02408_),
    .A2(_02448_),
    .A3(_02477_),
    .A4(_02481_),
    .ZN(_02482_));
 NAND4_X4 _11510_ (.A1(_02256_),
    .A2(_02264_),
    .A3(_02427_),
    .A4(_02290_),
    .ZN(_02483_));
 OAI21_X2 _11511_ (.A(_02467_),
    .B1(_02483_),
    .B2(_02445_),
    .ZN(_02484_));
 XOR2_X2 _11512_ (.A(_02470_),
    .B(_02484_),
    .Z(_02485_));
 NOR2_X1 _11513_ (.A1(_02259_),
    .A2(_02474_),
    .ZN(_02486_));
 OAI22_X4 _11514_ (.A1(_02174_),
    .A2(_02258_),
    .B1(_02469_),
    .B2(_02474_),
    .ZN(_02487_));
 NAND2_X2 _11515_ (.A1(_02196_),
    .A2(_02232_),
    .ZN(_02488_));
 AOI21_X4 _11516_ (.A(_02486_),
    .B1(_02487_),
    .B2(_02488_),
    .ZN(_02489_));
 NOR2_X1 _11517_ (.A1(_02455_),
    .A2(_02456_),
    .ZN(_02490_));
 MUX2_X2 _11518_ (.A(_02490_),
    .B(_02332_),
    .S(net17),
    .Z(_02491_));
 NAND4_X4 _11519_ (.A1(_02234_),
    .A2(_02254_),
    .A3(_02380_),
    .A4(_02383_),
    .ZN(_02492_));
 OAI21_X1 _11520_ (.A(_02244_),
    .B1(_02238_),
    .B2(_02237_),
    .ZN(_02493_));
 NAND2_X1 _11521_ (.A1(_02381_),
    .A2(_02488_),
    .ZN(_02494_));
 NOR2_X1 _11522_ (.A1(_02254_),
    .A2(_02455_),
    .ZN(_02495_));
 NAND3_X1 _11523_ (.A1(_02493_),
    .A2(_02494_),
    .A3(_02495_),
    .ZN(_02496_));
 XNOR2_X2 _11524_ (.A(_02355_),
    .B(_02405_),
    .ZN(_02497_));
 OAI221_X2 _11525_ (.A(_02385_),
    .B1(_02491_),
    .B2(_02492_),
    .C1(_02496_),
    .C2(_02497_),
    .ZN(_02498_));
 NOR2_X4 _11526_ (.A1(_02491_),
    .A2(_02492_),
    .ZN(_02499_));
 OAI221_X2 _11527_ (.A(_02489_),
    .B1(_02498_),
    .B2(_02353_),
    .C1(_02256_),
    .C2(_02499_),
    .ZN(_02500_));
 OAI21_X2 _11528_ (.A(_02335_),
    .B1(_02445_),
    .B2(_02483_),
    .ZN(_02501_));
 NAND2_X1 _11529_ (.A1(net17),
    .A2(_02378_),
    .ZN(_02502_));
 XNOR2_X2 _11530_ (.A(_02377_),
    .B(_02502_),
    .ZN(_02503_));
 XOR2_X2 _11531_ (.A(_02501_),
    .B(_02503_),
    .Z(_02504_));
 NOR3_X1 _11532_ (.A1(_02413_),
    .A2(_02417_),
    .A3(_02420_),
    .ZN(_02505_));
 AOI21_X4 _11533_ (.A(_02382_),
    .B1(net17),
    .B2(_02381_),
    .ZN(_02506_));
 OAI21_X1 _11534_ (.A(_02506_),
    .B1(_02350_),
    .B2(_01117_),
    .ZN(_02507_));
 AOI211_X2 _11535_ (.A(_02505_),
    .B(_02507_),
    .C1(_02265_),
    .C2(_02336_),
    .ZN(_02508_));
 NAND3_X1 _11536_ (.A1(_02256_),
    .A2(_02264_),
    .A3(_02423_),
    .ZN(_02509_));
 OAI211_X2 _11537_ (.A(_02290_),
    .B(_02335_),
    .C1(_02348_),
    .C2(_01117_),
    .ZN(_02510_));
 NOR2_X2 _11538_ (.A1(_01117_),
    .A2(_02350_),
    .ZN(_02511_));
 OAI33_X1 _11539_ (.A1(_02445_),
    .A2(_02509_),
    .A3(_02510_),
    .B1(_02511_),
    .B2(_02506_),
    .B3(_02421_),
    .ZN(_02512_));
 NOR2_X4 _11540_ (.A1(_02508_),
    .A2(_02512_),
    .ZN(_02513_));
 NOR4_X2 _11541_ (.A1(_02485_),
    .A2(_02500_),
    .A3(_02504_),
    .A4(_02513_),
    .ZN(_02514_));
 AOI211_X2 _11542_ (.A(_02354_),
    .B(_02370_),
    .C1(_02482_),
    .C2(_02514_),
    .ZN(_02515_));
 XNOR2_X2 _11543_ (.A(_01091_),
    .B(_02369_),
    .ZN(_02516_));
 OR4_X4 _11544_ (.A1(_02408_),
    .A2(_02448_),
    .A3(_02477_),
    .A4(_02513_),
    .ZN(_02517_));
 XNOR2_X2 _11545_ (.A(_02470_),
    .B(_02484_),
    .ZN(_02518_));
 OAI21_X2 _11546_ (.A(_02489_),
    .B1(_02499_),
    .B2(_02256_),
    .ZN(_02519_));
 AND3_X1 _11547_ (.A1(_02493_),
    .A2(_02494_),
    .A3(_02495_),
    .ZN(_02520_));
 XNOR2_X2 _11548_ (.A(_01090_),
    .B(_02405_),
    .ZN(_02521_));
 AOI211_X2 _11549_ (.A(_02384_),
    .B(_02499_),
    .C1(_02520_),
    .C2(_02521_),
    .ZN(_02522_));
 NAND2_X4 _11550_ (.A1(_02336_),
    .A2(_02265_),
    .ZN(_02523_));
 AOI21_X4 _11551_ (.A(_02519_),
    .B1(_02522_),
    .B2(_02523_),
    .ZN(_02524_));
 OR2_X4 _11552_ (.A1(_02369_),
    .A2(_02350_),
    .ZN(_02525_));
 AND2_X1 _11553_ (.A1(_02399_),
    .A2(_02525_),
    .ZN(_02526_));
 AND3_X1 _11554_ (.A1(_02355_),
    .A2(_02398_),
    .A3(_02525_),
    .ZN(_02527_));
 MUX2_X1 _11555_ (.A(_02526_),
    .B(_02527_),
    .S(_02405_),
    .Z(_02528_));
 OR2_X4 _11556_ (.A1(_02368_),
    .A2(_09034_),
    .ZN(_02529_));
 AND2_X1 _11557_ (.A1(_02350_),
    .A2(_02529_),
    .ZN(_02530_));
 NOR3_X1 _11558_ (.A1(_02530_),
    .A2(_02398_),
    .A3(_02355_),
    .ZN(_02531_));
 NOR3_X1 _11559_ (.A1(_02530_),
    .A2(_02414_),
    .A3(_02355_),
    .ZN(_02532_));
 MUX2_X1 _11560_ (.A(_02531_),
    .B(_02532_),
    .S(_02478_),
    .Z(_02533_));
 OAI22_X4 _11561_ (.A1(_02351_),
    .A2(_02352_),
    .B1(_02533_),
    .B2(_02528_),
    .ZN(_02534_));
 NOR4_X2 _11562_ (.A1(_02174_),
    .A2(_02266_),
    .A3(_02371_),
    .A4(_09001_),
    .ZN(_02535_));
 XNOR2_X1 _11563_ (.A(_01132_),
    .B(_01131_),
    .ZN(_02536_));
 AOI211_X2 _11564_ (.A(_01090_),
    .B(_02535_),
    .C1(_02536_),
    .C2(net17),
    .ZN(_02537_));
 AOI211_X2 _11565_ (.A(_02355_),
    .B(_02345_),
    .C1(_02346_),
    .C2(net2),
    .ZN(_02538_));
 OAI21_X2 _11566_ (.A(_02529_),
    .B1(_02537_),
    .B2(_02538_),
    .ZN(_02539_));
 NAND4_X2 _11567_ (.A1(_02265_),
    .A2(_02405_),
    .A3(_02336_),
    .A4(_02539_),
    .ZN(_02540_));
 NAND2_X2 _11568_ (.A1(_02534_),
    .A2(_02540_),
    .ZN(_02541_));
 XNOR2_X2 _11569_ (.A(_02501_),
    .B(_02503_),
    .ZN(_02542_));
 NAND4_X4 _11570_ (.A1(_02518_),
    .A2(_02524_),
    .A3(_02541_),
    .A4(_02542_),
    .ZN(_02543_));
 OAI21_X1 _11571_ (.A(_02516_),
    .B1(_02517_),
    .B2(_02543_),
    .ZN(_02544_));
 AOI21_X2 _11572_ (.A(_02515_),
    .B1(_02544_),
    .B2(_02354_),
    .ZN(_02545_));
 AND2_X4 _11573_ (.A1(_02540_),
    .A2(_02534_),
    .ZN(_02546_));
 NOR4_X4 _11574_ (.A1(_02504_),
    .A2(_02500_),
    .A3(_02485_),
    .A4(_02546_),
    .ZN(_02547_));
 NOR4_X4 _11575_ (.A1(_02408_),
    .A2(_02448_),
    .A3(_02477_),
    .A4(_02513_),
    .ZN(_02548_));
 CLKBUF_X2 _11576_ (.A(_09059_),
    .Z(_02549_));
 INV_X1 _11577_ (.A(_09061_),
    .ZN(_02550_));
 INV_X1 _11578_ (.A(_09046_),
    .ZN(_02551_));
 INV_X1 _11579_ (.A(_09052_),
    .ZN(_02552_));
 OAI21_X1 _11580_ (.A(_09053_),
    .B1(_09055_),
    .B2(_09056_),
    .ZN(_02553_));
 NAND2_X1 _11581_ (.A1(_02552_),
    .A2(_02553_),
    .ZN(_02554_));
 AND2_X2 _11582_ (.A1(_02554_),
    .A2(_09050_),
    .ZN(_02555_));
 OAI21_X4 _11583_ (.A(_09047_),
    .B1(_02555_),
    .B2(_09049_),
    .ZN(_02556_));
 NAND2_X4 _11584_ (.A1(_02556_),
    .A2(_02551_),
    .ZN(_02557_));
 AND2_X4 _11585_ (.A1(_09065_),
    .A2(_02557_),
    .ZN(_02558_));
 OAI21_X4 _11586_ (.A(_09062_),
    .B1(_09064_),
    .B2(_02558_),
    .ZN(_02559_));
 NAND2_X4 _11587_ (.A1(_02559_),
    .A2(_02550_),
    .ZN(_02560_));
 AND2_X4 _11588_ (.A1(_02549_),
    .A2(_02560_),
    .ZN(_02561_));
 OR2_X4 _11589_ (.A1(_02561_),
    .A2(_09058_),
    .ZN(_02562_));
 NAND2_X1 _11590_ (.A1(_01090_),
    .A2(_02562_),
    .ZN(_02563_));
 AOI21_X2 _11591_ (.A(_01960_),
    .B1(_02356_),
    .B2(_02562_),
    .ZN(_02564_));
 NOR2_X1 _11592_ (.A1(_08915_),
    .A2(_01965_),
    .ZN(_08937_));
 OR3_X1 _11593_ (.A1(_08939_),
    .A2(_08942_),
    .A3(_08941_),
    .ZN(_02565_));
 AND2_X1 _11594_ (.A1(_01822_),
    .A2(_02565_),
    .ZN(_02566_));
 MUX2_X1 _11595_ (.A(_08937_),
    .B(_02566_),
    .S(_01916_),
    .Z(_08955_));
 XOR2_X1 _11596_ (.A(_08957_),
    .B(_01922_),
    .Z(_02567_));
 MUX2_X1 _11597_ (.A(_08955_),
    .B(_02567_),
    .S(_02017_),
    .Z(_08972_));
 XNOR2_X1 _11598_ (.A(_01140_),
    .B(_02143_),
    .ZN(_02568_));
 MUX2_X1 _11599_ (.A(_08972_),
    .B(_02568_),
    .S(_02344_),
    .Z(_08992_));
 XOR2_X1 _11600_ (.A(_08994_),
    .B(_01130_),
    .Z(_02569_));
 MUX2_X1 _11601_ (.A(_08992_),
    .B(_02569_),
    .S(_02347_),
    .Z(_09013_));
 XNOR2_X1 _11602_ (.A(_02321_),
    .B(_02395_),
    .ZN(_02570_));
 MUX2_X2 _11603_ (.A(_09013_),
    .B(_02570_),
    .S(_02523_),
    .Z(_09033_));
 MUX2_X2 _11604_ (.A(_02563_),
    .B(_02564_),
    .S(_09033_),
    .Z(_02571_));
 AND3_X2 _11605_ (.A1(_02547_),
    .A2(_02548_),
    .A3(_02571_),
    .ZN(_02572_));
 BUF_X4 _11606_ (.A(_01960_),
    .Z(_02573_));
 XOR2_X2 _11607_ (.A(_09035_),
    .B(_02367_),
    .Z(_02574_));
 NAND2_X1 _11608_ (.A1(_02573_),
    .A2(_02574_),
    .ZN(_02575_));
 OR2_X1 _11609_ (.A1(_02356_),
    .A2(_02574_),
    .ZN(_02576_));
 NAND2_X1 _11610_ (.A1(_02356_),
    .A2(_02574_),
    .ZN(_02577_));
 AND2_X1 _11611_ (.A1(_02576_),
    .A2(_02577_),
    .ZN(_02578_));
 NOR2_X4 _11612_ (.A1(_09058_),
    .A2(_02561_),
    .ZN(_02579_));
 OAI21_X2 _11613_ (.A(_02575_),
    .B1(_02578_),
    .B2(_02579_),
    .ZN(_02580_));
 AOI21_X1 _11614_ (.A(_02580_),
    .B1(_02548_),
    .B2(_02547_),
    .ZN(_02581_));
 OR2_X1 _11615_ (.A1(_02572_),
    .A2(_02581_),
    .ZN(_02582_));
 NOR2_X2 _11616_ (.A1(_02545_),
    .A2(_02582_),
    .ZN(_02583_));
 AND2_X1 _11617_ (.A1(_02545_),
    .A2(_02582_),
    .ZN(_02584_));
 BUF_X8 _11618_ (.A(_02523_),
    .Z(_02585_));
 AOI21_X2 _11619_ (.A(_02252_),
    .B1(net17),
    .B2(_02249_),
    .ZN(_02586_));
 OAI21_X2 _11620_ (.A(_02586_),
    .B1(_02491_),
    .B2(_02384_),
    .ZN(_02587_));
 OR3_X2 _11621_ (.A1(_02384_),
    .A2(_02491_),
    .A3(_02586_),
    .ZN(_02588_));
 NAND3_X4 _11622_ (.A1(net35),
    .A2(_02587_),
    .A3(_02588_),
    .ZN(_02589_));
 OAI211_X2 _11623_ (.A(_02467_),
    .B(_02470_),
    .C1(_02445_),
    .C2(_02483_),
    .ZN(_02590_));
 XNOR2_X1 _11624_ (.A(_02590_),
    .B(_02489_),
    .ZN(_02591_));
 NAND3_X1 _11625_ (.A1(_02518_),
    .A2(_02589_),
    .A3(_02591_),
    .ZN(_02592_));
 NOR4_X4 _11626_ (.A1(_01117_),
    .A2(_02351_),
    .A3(_02352_),
    .A4(_02348_),
    .ZN(_02593_));
 AOI221_X2 _11627_ (.A(_02593_),
    .B1(_02540_),
    .B2(_02534_),
    .C1(_02523_),
    .C2(_02511_),
    .ZN(_02594_));
 NAND2_X1 _11628_ (.A1(_02542_),
    .A2(_02594_),
    .ZN(_02595_));
 NOR2_X1 _11629_ (.A1(_02421_),
    .A2(_02353_),
    .ZN(_02596_));
 XNOR2_X2 _11630_ (.A(_02506_),
    .B(_02596_),
    .ZN(_02597_));
 AOI21_X2 _11631_ (.A(_02592_),
    .B1(_02595_),
    .B2(_02597_),
    .ZN(_02598_));
 AND3_X1 _11632_ (.A1(_02542_),
    .A2(_02513_),
    .A3(_02594_),
    .ZN(_02599_));
 NOR2_X2 _11633_ (.A1(_02542_),
    .A2(_02594_),
    .ZN(_02600_));
 NOR2_X4 _11634_ (.A1(_02599_),
    .A2(_02600_),
    .ZN(_02601_));
 NOR3_X4 _11635_ (.A1(_02546_),
    .A2(_02504_),
    .A3(_02513_),
    .ZN(_02602_));
 NAND2_X2 _11636_ (.A1(_02518_),
    .A2(_02524_),
    .ZN(_02603_));
 OR3_X2 _11637_ (.A1(_02408_),
    .A2(_02448_),
    .A3(_02477_),
    .ZN(_02604_));
 OAI21_X4 _11638_ (.A(_02602_),
    .B1(_02603_),
    .B2(_02604_),
    .ZN(_02605_));
 OR2_X2 _11639_ (.A1(_02508_),
    .A2(_02512_),
    .ZN(_02606_));
 NAND3_X2 _11640_ (.A1(_02541_),
    .A2(_02542_),
    .A3(_02606_),
    .ZN(_02607_));
 OAI21_X1 _11641_ (.A(_02506_),
    .B1(_02499_),
    .B2(_02256_),
    .ZN(_02608_));
 AOI211_X2 _11642_ (.A(_02413_),
    .B(_02499_),
    .C1(_02520_),
    .C2(_02521_),
    .ZN(_02609_));
 AOI21_X1 _11643_ (.A(_02608_),
    .B1(_02609_),
    .B2(net35),
    .ZN(_02610_));
 AND3_X1 _11644_ (.A1(_02542_),
    .A2(_02594_),
    .A3(_02610_),
    .ZN(_02611_));
 NOR2_X1 _11645_ (.A1(_02233_),
    .A2(_02250_),
    .ZN(_02612_));
 OAI21_X1 _11646_ (.A(_02586_),
    .B1(_02398_),
    .B2(_02497_),
    .ZN(_02613_));
 NOR3_X2 _11647_ (.A1(_02384_),
    .A2(_02353_),
    .A3(_02613_),
    .ZN(_02614_));
 XNOR2_X2 _11648_ (.A(_02612_),
    .B(_02614_),
    .ZN(_02615_));
 OAI21_X2 _11649_ (.A(_02607_),
    .B1(_02611_),
    .B2(_02615_),
    .ZN(_02616_));
 AND4_X1 _11650_ (.A1(_02598_),
    .A2(_02601_),
    .A3(_02605_),
    .A4(_02616_),
    .ZN(_02617_));
 BUF_X4 _11651_ (.A(_02617_),
    .Z(_02618_));
 NAND2_X1 _11652_ (.A1(_02405_),
    .A2(_02529_),
    .ZN(_02619_));
 NOR4_X1 _11653_ (.A1(_02459_),
    .A2(_02445_),
    .A3(_02483_),
    .A4(_02619_),
    .ZN(_02620_));
 NAND3_X1 _11654_ (.A1(_02478_),
    .A2(_02414_),
    .A3(_02529_),
    .ZN(_02621_));
 AOI21_X1 _11655_ (.A(_02621_),
    .B1(_02451_),
    .B2(net19),
    .ZN(_02622_));
 NAND2_X1 _11656_ (.A1(_02398_),
    .A2(_02529_),
    .ZN(_02623_));
 OAI221_X1 _11657_ (.A(_02356_),
    .B1(_02446_),
    .B2(_02621_),
    .C1(_02623_),
    .C2(_02478_),
    .ZN(_02624_));
 NOR3_X1 _11658_ (.A1(_02620_),
    .A2(_02622_),
    .A3(_02624_),
    .ZN(_02625_));
 NOR2_X1 _11659_ (.A1(_01960_),
    .A2(_02478_),
    .ZN(_02626_));
 NAND4_X1 _11660_ (.A1(_02265_),
    .A2(_02336_),
    .A3(_02539_),
    .A4(_02626_),
    .ZN(_02627_));
 OAI21_X1 _11661_ (.A(_01117_),
    .B1(_02528_),
    .B2(_02533_),
    .ZN(_02628_));
 OAI221_X2 _11662_ (.A(_02627_),
    .B1(_02628_),
    .B2(_02353_),
    .C1(_02356_),
    .C2(_02369_),
    .ZN(_02629_));
 AOI211_X2 _11663_ (.A(_02625_),
    .B(_02629_),
    .C1(_02481_),
    .C2(_01960_),
    .ZN(_02630_));
 NOR2_X1 _11664_ (.A1(_02356_),
    .A2(_02369_),
    .ZN(_02631_));
 AOI21_X2 _11665_ (.A(_02354_),
    .B1(_02631_),
    .B2(_02481_),
    .ZN(_02632_));
 NOR2_X2 _11666_ (.A1(_02630_),
    .A2(_02632_),
    .ZN(_02633_));
 NOR3_X4 _11667_ (.A1(_02408_),
    .A2(_02448_),
    .A3(_02477_),
    .ZN(_02634_));
 NOR4_X4 _11668_ (.A1(_02408_),
    .A2(_02448_),
    .A3(_02485_),
    .A4(_02500_),
    .ZN(_02635_));
 AOI21_X4 _11669_ (.A(_02634_),
    .B1(_02602_),
    .B2(_02635_),
    .ZN(_02636_));
 NAND3_X4 _11670_ (.A1(_02547_),
    .A2(_02548_),
    .A3(_02571_),
    .ZN(_02637_));
 NOR2_X2 _11671_ (.A1(_02354_),
    .A2(_02370_),
    .ZN(_02638_));
 OR3_X2 _11672_ (.A1(_02580_),
    .A2(_02594_),
    .A3(_02638_),
    .ZN(_02639_));
 AOI211_X2 _11673_ (.A(_02633_),
    .B(_02636_),
    .C1(_02637_),
    .C2(_02639_),
    .ZN(_02640_));
 NAND2_X4 _11674_ (.A1(_02618_),
    .A2(_02640_),
    .ZN(_02641_));
 BUF_X8 _11675_ (.A(_02641_),
    .Z(_02642_));
 AOI21_X2 _11676_ (.A(_02583_),
    .B1(_02584_),
    .B2(net18),
    .ZN(_02643_));
 CLKBUF_X3 _11677_ (.A(_02356_),
    .Z(_02644_));
 BUF_X2 _11678_ (.A(_09082_),
    .Z(_02645_));
 INV_X1 _11679_ (.A(_09084_),
    .ZN(_02646_));
 INV_X1 _11680_ (.A(_09067_),
    .ZN(_02647_));
 BUF_X2 _11681_ (.A(_09085_),
    .Z(_02648_));
 INV_X1 _11682_ (.A(_02648_),
    .ZN(_02649_));
 OAI21_X1 _11683_ (.A(_02646_),
    .B1(_02647_),
    .B2(_02649_),
    .ZN(_02650_));
 NAND2_X1 _11684_ (.A1(_02645_),
    .A2(_02650_),
    .ZN(_02651_));
 NOR2_X1 _11685_ (.A1(_02644_),
    .A2(_02651_),
    .ZN(_02652_));
 INV_X1 _11686_ (.A(_09081_),
    .ZN(_02653_));
 INV_X1 _11687_ (.A(_09070_),
    .ZN(_02654_));
 BUF_X1 _11688_ (.A(_09071_),
    .Z(_02655_));
 INV_X1 _11689_ (.A(_09076_),
    .ZN(_02656_));
 BUF_X1 rebuffer56 (.A(net415),
    .Z(net414));
 OAI21_X2 _11691_ (.A(_09077_),
    .B1(_09078_),
    .B2(_09079_),
    .ZN(_02658_));
 NAND2_X2 _11692_ (.A1(_02656_),
    .A2(_02658_),
    .ZN(_02659_));
 AND2_X4 _11693_ (.A1(_09074_),
    .A2(_02659_),
    .ZN(_02660_));
 OAI21_X2 _11694_ (.A(_02655_),
    .B1(_02660_),
    .B2(_09073_),
    .ZN(_02661_));
 NAND2_X2 _11695_ (.A1(_02654_),
    .A2(_02661_),
    .ZN(_02662_));
 NAND4_X4 _11696_ (.A1(_09068_),
    .A2(_02645_),
    .A3(_02648_),
    .A4(_02662_),
    .ZN(_02663_));
 NAND2_X4 _11697_ (.A1(_02653_),
    .A2(_02663_),
    .ZN(_02664_));
 INV_X4 _11698_ (.A(_02664_),
    .ZN(_02665_));
 NOR2_X2 _11699_ (.A1(_02644_),
    .A2(_02665_),
    .ZN(_02666_));
 NOR2_X1 _11700_ (.A1(_02666_),
    .A2(_02652_),
    .ZN(_02667_));
 OAI21_X1 _11701_ (.A(_01117_),
    .B1(_01091_),
    .B2(_02651_),
    .ZN(_02668_));
 INV_X1 _11702_ (.A(_02668_),
    .ZN(_02669_));
 NOR2_X4 _11703_ (.A1(_08940_),
    .A2(_01916_),
    .ZN(_02670_));
 AOI21_X2 _11704_ (.A(_02670_),
    .B1(_01916_),
    .B2(_08942_),
    .ZN(_08958_));
 OR3_X1 _11705_ (.A1(_08960_),
    .A2(_01920_),
    .A3(_08961_),
    .ZN(_02671_));
 AND2_X1 _11706_ (.A1(_01921_),
    .A2(_02671_),
    .ZN(_02672_));
 MUX2_X1 _11707_ (.A(_08958_),
    .B(_02672_),
    .S(_02017_),
    .Z(_08975_));
 AND2_X1 _11708_ (.A1(_01699_),
    .A2(_01698_),
    .ZN(_02673_));
 XNOR2_X1 _11709_ (.A(_08977_),
    .B(_02673_),
    .ZN(_02674_));
 MUX2_X1 _11710_ (.A(_08975_),
    .B(_02674_),
    .S(_02344_),
    .Z(_08995_));
 OR3_X1 _11711_ (.A1(_08997_),
    .A2(_08987_),
    .A3(_01128_),
    .ZN(_02675_));
 AND2_X1 _11712_ (.A1(_01129_),
    .A2(_02675_),
    .ZN(_02676_));
 MUX2_X1 _11713_ (.A(_08995_),
    .B(_02676_),
    .S(_02347_),
    .Z(_09016_));
 XNOR2_X1 _11714_ (.A(_02318_),
    .B(_02317_),
    .ZN(_02677_));
 MUX2_X2 _11715_ (.A(_09016_),
    .B(_02677_),
    .S(_02585_),
    .Z(_09036_));
 NAND3_X2 _11716_ (.A1(_02547_),
    .A2(_02548_),
    .A3(_09036_),
    .ZN(_02678_));
 XNOR2_X1 _11717_ (.A(_09038_),
    .B(_02365_),
    .ZN(_02679_));
 OAI21_X2 _11718_ (.A(_02679_),
    .B1(_02517_),
    .B2(_02543_),
    .ZN(_02680_));
 NAND2_X1 _11719_ (.A1(_02678_),
    .A2(_02680_),
    .ZN(_09057_));
 MUX2_X1 _11720_ (.A(_02667_),
    .B(_02669_),
    .S(_09057_),
    .Z(_02681_));
 XNOR2_X2 _11721_ (.A(_02549_),
    .B(_02560_),
    .ZN(_02682_));
 MUX2_X1 _11722_ (.A(_02668_),
    .B(_02652_),
    .S(_02682_),
    .Z(_02683_));
 INV_X1 _11723_ (.A(_02683_),
    .ZN(_02684_));
 MUX2_X2 _11724_ (.A(_02681_),
    .B(_02684_),
    .S(_02641_),
    .Z(_02685_));
 NAND4_X4 _11725_ (.A1(_02598_),
    .A2(_02601_),
    .A3(_02605_),
    .A4(_02616_),
    .ZN(_02686_));
 OR2_X2 _11726_ (.A1(_02630_),
    .A2(_02632_),
    .ZN(_02687_));
 AND2_X1 _11727_ (.A1(_02602_),
    .A2(_02635_),
    .ZN(_02688_));
 NOR3_X4 _11728_ (.A1(_02580_),
    .A2(_02594_),
    .A3(_02638_),
    .ZN(_02689_));
 OAI221_X2 _11729_ (.A(_02687_),
    .B1(_02688_),
    .B2(_02634_),
    .C1(_02572_),
    .C2(_02689_),
    .ZN(_02690_));
 AND2_X1 _11730_ (.A1(_02666_),
    .A2(_02682_),
    .ZN(_02691_));
 NAND2_X1 _11731_ (.A1(_02644_),
    .A2(_02664_),
    .ZN(_02692_));
 NOR2_X1 _11732_ (.A1(_02682_),
    .A2(_02692_),
    .ZN(_02693_));
 OAI22_X2 _11733_ (.A1(_02686_),
    .A2(_02690_),
    .B1(_02691_),
    .B2(_02693_),
    .ZN(_02694_));
 AOI21_X1 _11734_ (.A(_02692_),
    .B1(_02680_),
    .B2(_02678_),
    .ZN(_02695_));
 NAND3_X1 _11735_ (.A1(_02618_),
    .A2(_02640_),
    .A3(_02695_),
    .ZN(_02696_));
 AND2_X4 _11736_ (.A1(_02696_),
    .A2(_02694_),
    .ZN(_02697_));
 NAND2_X4 _11737_ (.A1(_02548_),
    .A2(_02547_),
    .ZN(_02698_));
 MUX2_X2 _11738_ (.A(_09033_),
    .B(_02574_),
    .S(_02698_),
    .Z(_02699_));
 NAND4_X1 _11739_ (.A1(_02518_),
    .A2(_02524_),
    .A3(_02542_),
    .A4(_02606_),
    .ZN(_02700_));
 OAI21_X1 _11740_ (.A(_02638_),
    .B1(_02481_),
    .B2(_02700_),
    .ZN(_02701_));
 AOI21_X2 _11741_ (.A(_02354_),
    .B1(_02516_),
    .B2(_02604_),
    .ZN(_02702_));
 NAND2_X1 _11742_ (.A1(_02354_),
    .A2(_02516_),
    .ZN(_02703_));
 AOI21_X2 _11743_ (.A(_02703_),
    .B1(_02548_),
    .B2(_02547_),
    .ZN(_02704_));
 OAI21_X1 _11744_ (.A(_02701_),
    .B1(_02702_),
    .B2(_02704_),
    .ZN(_02705_));
 NOR3_X1 _11745_ (.A1(_01547_),
    .A2(_02562_),
    .A3(_02705_),
    .ZN(_02706_));
 XNOR2_X2 _11746_ (.A(_02644_),
    .B(_02579_),
    .ZN(_02707_));
 XNOR2_X1 _11747_ (.A(_02699_),
    .B(_02707_),
    .ZN(_02708_));
 OAI33_X1 _11748_ (.A1(_02699_),
    .A2(_02641_),
    .A3(_02705_),
    .B1(_02706_),
    .B2(_02583_),
    .B3(_02708_),
    .ZN(_02709_));
 NOR2_X4 _11749_ (.A1(_02543_),
    .A2(_02517_),
    .ZN(_02710_));
 NAND4_X1 _11750_ (.A1(_02541_),
    .A2(_02542_),
    .A3(_02606_),
    .A4(_02589_),
    .ZN(_02711_));
 AOI21_X1 _11751_ (.A(_02611_),
    .B1(_02615_),
    .B2(_02711_),
    .ZN(_02712_));
 OR2_X2 _11752_ (.A1(_02710_),
    .A2(_02712_),
    .ZN(_02713_));
 OR2_X1 _11753_ (.A1(_02518_),
    .A2(_02611_),
    .ZN(_02714_));
 NAND2_X1 _11754_ (.A1(_02597_),
    .A2(_02595_),
    .ZN(_02715_));
 AND2_X1 _11755_ (.A1(_02715_),
    .A2(_02605_),
    .ZN(_02716_));
 AND3_X1 _11756_ (.A1(_02713_),
    .A2(_02714_),
    .A3(_02716_),
    .ZN(_02717_));
 NAND2_X1 _11757_ (.A1(_02601_),
    .A2(_02605_),
    .ZN(_02718_));
 AOI21_X2 _11758_ (.A(_02593_),
    .B1(_02511_),
    .B2(net35),
    .ZN(_02719_));
 NAND2_X1 _11759_ (.A1(_02541_),
    .A2(_02719_),
    .ZN(_02720_));
 XNOR2_X1 _11760_ (.A(_02405_),
    .B(_02480_),
    .ZN(_02721_));
 INV_X1 _11761_ (.A(_02719_),
    .ZN(_02722_));
 XNOR2_X1 _11762_ (.A(_02644_),
    .B(_02354_),
    .ZN(_02723_));
 AOI21_X1 _11763_ (.A(_02722_),
    .B1(_02723_),
    .B2(_02529_),
    .ZN(_02724_));
 OAI22_X2 _11764_ (.A1(_02710_),
    .A2(_02720_),
    .B1(_02721_),
    .B2(_02724_),
    .ZN(_02725_));
 OAI221_X2 _11765_ (.A(_02701_),
    .B1(_02702_),
    .B2(_02704_),
    .C1(_02581_),
    .C2(_02572_),
    .ZN(_02726_));
 AOI21_X2 _11766_ (.A(_02718_),
    .B1(_02725_),
    .B2(_02726_),
    .ZN(_02727_));
 XOR2_X2 _11767_ (.A(_02589_),
    .B(_02605_),
    .Z(_02728_));
 AOI21_X4 _11768_ (.A(_02633_),
    .B1(_02639_),
    .B2(_02637_),
    .ZN(_02729_));
 OAI22_X1 _11769_ (.A1(_02686_),
    .A2(_02690_),
    .B1(_02728_),
    .B2(_02729_),
    .ZN(_02730_));
 AND3_X2 _11770_ (.A1(_02717_),
    .A2(_02727_),
    .A3(_02730_),
    .ZN(_02731_));
 NAND4_X4 _11771_ (.A1(_02685_),
    .A2(_02697_),
    .A3(net379),
    .A4(_02731_),
    .ZN(_02732_));
 INV_X1 _11772_ (.A(_02408_),
    .ZN(_02733_));
 INV_X1 _11773_ (.A(_02477_),
    .ZN(_02734_));
 NOR2_X1 _11774_ (.A1(_02733_),
    .A2(_02734_),
    .ZN(_02735_));
 OR2_X2 _11775_ (.A1(_02408_),
    .A2(_02477_),
    .ZN(_02736_));
 NOR4_X2 _11776_ (.A1(_02736_),
    .A2(_02634_),
    .A3(_02603_),
    .A4(_02607_),
    .ZN(_02737_));
 OR2_X1 _11777_ (.A1(_02735_),
    .A2(_02737_),
    .ZN(_02738_));
 OAI21_X4 _11778_ (.A(_02687_),
    .B1(_02689_),
    .B2(_02572_),
    .ZN(_02739_));
 AOI21_X2 _11779_ (.A(_02433_),
    .B1(net29),
    .B2(_01150_),
    .ZN(_02740_));
 NAND4_X2 _11780_ (.A1(net19),
    .A2(_02451_),
    .A3(_02446_),
    .A4(_02740_),
    .ZN(_02741_));
 NOR2_X4 _11781_ (.A1(_02103_),
    .A2(_02112_),
    .ZN(_02742_));
 OAI21_X2 _11782_ (.A(_02742_),
    .B1(_02445_),
    .B2(_02459_),
    .ZN(_02743_));
 AOI21_X2 _11783_ (.A(_02109_),
    .B1(net29),
    .B2(_01150_),
    .ZN(_02744_));
 NOR3_X4 _11784_ (.A1(_01710_),
    .A2(_02434_),
    .A3(_02744_),
    .ZN(_02745_));
 AOI21_X2 _11785_ (.A(_02745_),
    .B1(_02742_),
    .B2(_02483_),
    .ZN(_02746_));
 NAND4_X1 _11786_ (.A1(_09047_),
    .A2(_09056_),
    .A3(_09050_),
    .A4(_09053_),
    .ZN(_02747_));
 NAND3_X1 _11787_ (.A1(_02549_),
    .A2(_09062_),
    .A3(_09065_),
    .ZN(_02748_));
 NOR3_X1 _11788_ (.A1(_01170_),
    .A2(_02747_),
    .A3(_02748_),
    .ZN(_02749_));
 AND4_X1 _11789_ (.A1(_02741_),
    .A2(_02743_),
    .A3(_02746_),
    .A4(_02749_),
    .ZN(_02750_));
 NOR2_X2 _11790_ (.A1(_01596_),
    .A2(net9),
    .ZN(_02751_));
 AOI21_X4 _11791_ (.A(_08940_),
    .B1(net29),
    .B2(_02751_),
    .ZN(_02752_));
 NAND2_X1 _11792_ (.A1(_02750_),
    .A2(_02752_),
    .ZN(_02753_));
 AOI221_X2 _11793_ (.A(_02753_),
    .B1(_02577_),
    .B2(_02576_),
    .C1(_02547_),
    .C2(_02548_),
    .ZN(_02754_));
 NAND4_X1 _11794_ (.A1(_02356_),
    .A2(_09033_),
    .A3(_02750_),
    .A4(_02752_),
    .ZN(_02755_));
 NOR3_X2 _11795_ (.A1(_02543_),
    .A2(_02517_),
    .A3(_02755_),
    .ZN(_02756_));
 NAND3_X4 _11796_ (.A1(_02741_),
    .A2(_02743_),
    .A3(_02746_),
    .ZN(_02757_));
 NAND2_X1 _11797_ (.A1(_02749_),
    .A2(_02752_),
    .ZN(_02758_));
 OR4_X1 _11798_ (.A1(_02356_),
    .A2(_09033_),
    .A3(_02757_),
    .A4(_02758_),
    .ZN(_02759_));
 NOR3_X2 _11799_ (.A1(_02543_),
    .A2(_02517_),
    .A3(_02759_),
    .ZN(_02760_));
 NOR4_X4 _11800_ (.A1(_02636_),
    .A2(_02754_),
    .A3(_02756_),
    .A4(_02760_),
    .ZN(_02761_));
 NOR4_X4 _11801_ (.A1(_02736_),
    .A2(_02739_),
    .A3(_02686_),
    .A4(_02761_),
    .ZN(_02762_));
 OR4_X1 _11802_ (.A1(_02636_),
    .A2(_02754_),
    .A3(_02756_),
    .A4(_02760_),
    .ZN(_02763_));
 NAND3_X1 _11803_ (.A1(_02729_),
    .A2(_02618_),
    .A3(_02763_),
    .ZN(_02764_));
 NOR2_X1 _11804_ (.A1(_02603_),
    .A2(_02607_),
    .ZN(_02765_));
 NOR2_X1 _11805_ (.A1(_02733_),
    .A2(_02765_),
    .ZN(_02766_));
 AOI211_X2 _11806_ (.A(_02738_),
    .B(_02762_),
    .C1(_02764_),
    .C2(_02766_),
    .ZN(_02767_));
 NOR3_X4 _11807_ (.A1(_02739_),
    .A2(_02686_),
    .A3(_02761_),
    .ZN(_02768_));
 AND3_X1 _11808_ (.A1(_02518_),
    .A2(_02715_),
    .A3(_02589_),
    .ZN(_02769_));
 AND2_X2 _11809_ (.A1(_02601_),
    .A2(_02605_),
    .ZN(_02770_));
 NAND4_X2 _11810_ (.A1(_02729_),
    .A2(_02769_),
    .A3(_02770_),
    .A4(_02713_),
    .ZN(_02771_));
 AOI21_X1 _11811_ (.A(_02591_),
    .B1(_02611_),
    .B2(_02518_),
    .ZN(_02772_));
 AOI21_X1 _11812_ (.A(_02772_),
    .B1(_02765_),
    .B2(_02604_),
    .ZN(_02773_));
 INV_X1 _11813_ (.A(_02773_),
    .ZN(_02774_));
 AOI21_X4 _11814_ (.A(_02768_),
    .B1(_02771_),
    .B2(_02774_),
    .ZN(_02775_));
 OR2_X1 _11815_ (.A1(_02408_),
    .A2(_02448_),
    .ZN(_02776_));
 NOR2_X1 _11816_ (.A1(_02485_),
    .A2(_02500_),
    .ZN(_02777_));
 NAND4_X1 _11817_ (.A1(_02776_),
    .A2(_02734_),
    .A3(_02777_),
    .A4(_02602_),
    .ZN(_02778_));
 OAI21_X1 _11818_ (.A(_02477_),
    .B1(_02603_),
    .B2(_02607_),
    .ZN(_02779_));
 NAND2_X1 _11819_ (.A1(_02778_),
    .A2(_02779_),
    .ZN(_02780_));
 XNOR2_X2 _11820_ (.A(_02768_),
    .B(_02780_),
    .ZN(_02781_));
 NAND3_X1 _11821_ (.A1(_02425_),
    .A2(_02777_),
    .A3(_02602_),
    .ZN(_02782_));
 OAI21_X1 _11822_ (.A(_02448_),
    .B1(_02736_),
    .B2(_02782_),
    .ZN(_02783_));
 NAND2_X1 _11823_ (.A1(_02430_),
    .A2(_02447_),
    .ZN(_02784_));
 NOR2_X2 _11824_ (.A1(_02408_),
    .A2(_02784_),
    .ZN(_02785_));
 NAND3_X1 _11825_ (.A1(_02547_),
    .A2(_02606_),
    .A3(_02785_),
    .ZN(_02786_));
 AOI21_X1 _11826_ (.A(_02425_),
    .B1(_02734_),
    .B2(_02785_),
    .ZN(_02787_));
 AOI221_X2 _11827_ (.A(_02633_),
    .B1(_02786_),
    .B2(_02787_),
    .C1(_02639_),
    .C2(_02637_),
    .ZN(_02788_));
 AOI21_X1 _11828_ (.A(_02783_),
    .B1(_02788_),
    .B2(_02618_),
    .ZN(_02789_));
 XNOR2_X2 _11829_ (.A(_02784_),
    .B(_02737_),
    .ZN(_02790_));
 AND3_X1 _11830_ (.A1(_02733_),
    .A2(_02778_),
    .A3(_02779_),
    .ZN(_02791_));
 AOI21_X1 _11831_ (.A(_02790_),
    .B1(_02791_),
    .B2(_02636_),
    .ZN(_02792_));
 AOI211_X2 _11832_ (.A(_02789_),
    .B(_02792_),
    .C1(_02790_),
    .C2(_02762_),
    .ZN(_02793_));
 NAND4_X4 _11833_ (.A1(_02767_),
    .A2(_02775_),
    .A3(_02781_),
    .A4(_02793_),
    .ZN(_02794_));
 NOR2_X4 _11834_ (.A1(_02794_),
    .A2(_02732_),
    .ZN(_02795_));
 BUF_X8 _11835_ (.A(_02795_),
    .Z(_02796_));
 BUF_X4 _11836_ (.A(_01117_),
    .Z(_02797_));
 OAI21_X1 _11837_ (.A(_02644_),
    .B1(_09081_),
    .B2(_02645_),
    .ZN(_02798_));
 NAND2_X1 _11838_ (.A1(_01150_),
    .A2(net29),
    .ZN(_02799_));
 OR3_X1 _11839_ (.A1(_02104_),
    .A2(_02112_),
    .A3(_02799_),
    .ZN(_02800_));
 OAI21_X1 _11840_ (.A(_02104_),
    .B1(_02112_),
    .B2(_02799_),
    .ZN(_02801_));
 AND2_X2 _11841_ (.A1(_02800_),
    .A2(_02801_),
    .ZN(_02802_));
 NOR2_X1 _11842_ (.A1(_01965_),
    .A2(_01882_),
    .ZN(_02803_));
 NAND2_X1 _11843_ (.A1(_02307_),
    .A2(_08890_),
    .ZN(_02804_));
 AOI21_X1 _11844_ (.A(_02803_),
    .B1(_02308_),
    .B2(_02804_),
    .ZN(_02805_));
 XNOR2_X1 _11845_ (.A(_02800_),
    .B(_02805_),
    .ZN(_02806_));
 NAND2_X1 _11846_ (.A1(_01710_),
    .A2(_02806_),
    .ZN(_02807_));
 OR3_X2 _11847_ (.A1(_02112_),
    .A2(_02802_),
    .A3(_02807_),
    .ZN(_02808_));
 AOI21_X2 _11848_ (.A(_02808_),
    .B1(_02451_),
    .B2(net19),
    .ZN(_02809_));
 NAND2_X1 _11849_ (.A1(_01710_),
    .A2(_02802_),
    .ZN(_02810_));
 NOR4_X4 _11850_ (.A1(_02459_),
    .A2(_02445_),
    .A3(_02483_),
    .A4(_02810_),
    .ZN(_02811_));
 NAND2_X1 _11851_ (.A1(_02112_),
    .A2(_02802_),
    .ZN(_02812_));
 OAI22_X4 _11852_ (.A1(_02446_),
    .A2(_02808_),
    .B1(_02812_),
    .B2(_02807_),
    .ZN(_02813_));
 NOR3_X4 _11853_ (.A1(_02809_),
    .A2(_02811_),
    .A3(_02813_),
    .ZN(_02814_));
 INV_X2 _11854_ (.A(_02752_),
    .ZN(_09007_));
 OAI211_X4 _11855_ (.A(_02742_),
    .B(_02802_),
    .C1(_02351_),
    .C2(_02352_),
    .ZN(_02815_));
 XNOR2_X2 _11856_ (.A(_09007_),
    .B(_02815_),
    .ZN(_02816_));
 AOI21_X1 _11857_ (.A(_09076_),
    .B1(_09078_),
    .B2(_09077_),
    .ZN(_02817_));
 INV_X1 _11858_ (.A(_02817_),
    .ZN(_02818_));
 NOR4_X2 _11859_ (.A1(_02757_),
    .A2(_02814_),
    .A3(_02816_),
    .A4(_02818_),
    .ZN(_02819_));
 AND2_X1 _11860_ (.A1(_09068_),
    .A2(_02655_),
    .ZN(_02820_));
 NAND2_X1 _11861_ (.A1(_02660_),
    .A2(_02820_),
    .ZN(_02821_));
 NOR2_X1 _11862_ (.A1(_02819_),
    .A2(_02821_),
    .ZN(_02822_));
 AOI21_X1 _11863_ (.A(_09070_),
    .B1(_09073_),
    .B2(_02655_),
    .ZN(_02823_));
 INV_X1 _11864_ (.A(_09068_),
    .ZN(_02824_));
 OAI21_X1 _11865_ (.A(_02647_),
    .B1(_02823_),
    .B2(_02824_),
    .ZN(_02825_));
 OAI21_X1 _11866_ (.A(_02648_),
    .B1(_02822_),
    .B2(_02825_),
    .ZN(_02826_));
 NOR3_X1 _11867_ (.A1(_02573_),
    .A2(_09081_),
    .A3(_09084_),
    .ZN(_02827_));
 AOI22_X2 _11868_ (.A1(_02797_),
    .A2(_02798_),
    .B1(_02826_),
    .B2(_02827_),
    .ZN(_02828_));
 AOI21_X2 _11869_ (.A(_02682_),
    .B1(_02640_),
    .B2(_02618_),
    .ZN(_02829_));
 AOI21_X2 _11870_ (.A(_02636_),
    .B1(_02678_),
    .B2(_02680_),
    .ZN(_02830_));
 AND3_X1 _11871_ (.A1(_02729_),
    .A2(_02618_),
    .A3(_02830_),
    .ZN(_02831_));
 OAI21_X2 _11872_ (.A(_02828_),
    .B1(_02829_),
    .B2(_02831_),
    .ZN(_02832_));
 INV_X1 _11873_ (.A(_02707_),
    .ZN(_02833_));
 OAI21_X4 _11874_ (.A(_02833_),
    .B1(_02690_),
    .B2(_02686_),
    .ZN(_02834_));
 XOR2_X2 _11875_ (.A(_02699_),
    .B(_02834_),
    .Z(_02835_));
 OAI21_X1 _11876_ (.A(_02645_),
    .B1(_02648_),
    .B2(_09084_),
    .ZN(_02836_));
 NAND2_X1 _11877_ (.A1(_02653_),
    .A2(_02836_),
    .ZN(_02837_));
 OR3_X1 _11878_ (.A1(_09081_),
    .A2(_09084_),
    .A3(_02825_),
    .ZN(_02838_));
 OAI21_X1 _11879_ (.A(_02837_),
    .B1(_02838_),
    .B2(_02822_),
    .ZN(_02839_));
 OR4_X2 _11880_ (.A1(_02644_),
    .A2(_02831_),
    .A3(_02829_),
    .A4(_02839_),
    .ZN(_02840_));
 NAND3_X1 _11881_ (.A1(_02832_),
    .A2(_02835_),
    .A3(_02840_),
    .ZN(_02841_));
 NOR2_X1 _11882_ (.A1(_02796_),
    .A2(_02841_),
    .ZN(_02842_));
 XOR2_X2 _11883_ (.A(_02643_),
    .B(_02842_),
    .Z(_02843_));
 AOI21_X2 _11884_ (.A(_02835_),
    .B1(_02697_),
    .B2(_02685_),
    .ZN(_02844_));
 NAND3_X2 _11885_ (.A1(_02729_),
    .A2(_02618_),
    .A3(_02830_),
    .ZN(_02845_));
 XOR2_X2 _11886_ (.A(_02549_),
    .B(_02560_),
    .Z(_02846_));
 OAI21_X2 _11887_ (.A(_02846_),
    .B1(_02690_),
    .B2(_02686_),
    .ZN(_02847_));
 NAND2_X2 _11888_ (.A1(_02845_),
    .A2(_02847_),
    .ZN(_02848_));
 XNOR2_X1 _11889_ (.A(_02644_),
    .B(_02839_),
    .ZN(_02849_));
 XNOR2_X2 _11890_ (.A(_02848_),
    .B(_02849_),
    .ZN(_02850_));
 AOI21_X1 _11891_ (.A(_02644_),
    .B1(_02651_),
    .B2(_02665_),
    .ZN(_02851_));
 MUX2_X1 _11892_ (.A(_02851_),
    .B(_02668_),
    .S(_09057_),
    .Z(_02852_));
 MUX2_X1 _11893_ (.A(_02852_),
    .B(_02683_),
    .S(net18),
    .Z(_02853_));
 NAND2_X1 _11894_ (.A1(_02694_),
    .A2(_02696_),
    .ZN(_02854_));
 XNOR2_X2 _11895_ (.A(_02699_),
    .B(_02834_),
    .ZN(_02855_));
 NOR3_X2 _11896_ (.A1(_02853_),
    .A2(_02854_),
    .A3(_02855_),
    .ZN(_02856_));
 NOR3_X2 _11897_ (.A1(_02844_),
    .A2(_02850_),
    .A3(_02856_),
    .ZN(_02857_));
 NOR2_X2 _11898_ (.A1(_02848_),
    .A2(_02855_),
    .ZN(_02858_));
 AOI21_X1 _11899_ (.A(_02857_),
    .B1(_02858_),
    .B2(_02796_),
    .ZN(_02859_));
 NOR2_X1 _11900_ (.A1(_01920_),
    .A2(_02064_),
    .ZN(_08978_));
 OR3_X1 _11901_ (.A1(_08980_),
    .A2(_01142_),
    .A3(_08982_),
    .ZN(_02860_));
 AND2_X1 _11902_ (.A1(_02141_),
    .A2(_02860_),
    .ZN(_02861_));
 MUX2_X1 _11903_ (.A(_08978_),
    .B(_02861_),
    .S(_02344_),
    .Z(_08986_));
 XOR2_X1 _11904_ (.A(_08988_),
    .B(_01127_),
    .Z(_02862_));
 MUX2_X1 _11905_ (.A(_08986_),
    .B(_02862_),
    .S(_02347_),
    .Z(_09019_));
 XNOR2_X1 _11906_ (.A(_02316_),
    .B(_02392_),
    .ZN(_02863_));
 MUX2_X1 _11907_ (.A(_09019_),
    .B(_02863_),
    .S(_02585_),
    .Z(_09039_));
 XOR2_X1 _11908_ (.A(_09041_),
    .B(_02364_),
    .Z(_02864_));
 MUX2_X1 _11909_ (.A(_09039_),
    .B(_02864_),
    .S(_02698_),
    .Z(_09060_));
 OR3_X1 _11910_ (.A1(_09062_),
    .A2(_09064_),
    .A3(_02558_),
    .ZN(_02865_));
 AND2_X1 _11911_ (.A1(_02559_),
    .A2(_02865_),
    .ZN(_02866_));
 MUX2_X2 _11912_ (.A(_09060_),
    .B(_02866_),
    .S(net18),
    .Z(_09080_));
 NOR3_X4 _11913_ (.A1(_02732_),
    .A2(_02794_),
    .A3(_09080_),
    .ZN(_02867_));
 CLKBUF_X3 _11914_ (.A(_02644_),
    .Z(_02868_));
 NAND2_X2 clone13 (.A1(_02886_),
    .A2(_02888_),
    .ZN(net13));
 AOI21_X2 _11916_ (.A(_09087_),
    .B1(_09088_),
    .B2(_09090_),
    .ZN(_02870_));
 INV_X2 _11917_ (.A(_02870_),
    .ZN(_02871_));
 BUF_X2 _11918_ (.A(_09106_),
    .Z(_02872_));
 AOI21_X4 _11919_ (.A(_09105_),
    .B1(_02872_),
    .B2(_02871_),
    .ZN(_02873_));
 OR2_X4 _11920_ (.A1(_02873_),
    .A2(_02868_),
    .ZN(_02874_));
 NAND2_X1 _11921_ (.A1(_09074_),
    .A2(_02659_),
    .ZN(_02875_));
 XNOR2_X1 _11922_ (.A(_02752_),
    .B(_02815_),
    .ZN(_02876_));
 AOI21_X1 _11923_ (.A(_02875_),
    .B1(_02876_),
    .B2(_02817_),
    .ZN(_02877_));
 OAI21_X1 _11924_ (.A(_02655_),
    .B1(_09073_),
    .B2(_02877_),
    .ZN(_02878_));
 AOI21_X1 _11925_ (.A(_02824_),
    .B1(_02654_),
    .B2(_02878_),
    .ZN(_02879_));
 NAND4_X2 _11926_ (.A1(_09079_),
    .A2(_09074_),
    .A3(_09077_),
    .A4(_02820_),
    .ZN(_02880_));
 NOR2_X1 _11927_ (.A1(_02880_),
    .A2(_02816_),
    .ZN(_02881_));
 NOR3_X1 _11928_ (.A1(_09067_),
    .A2(_02879_),
    .A3(_02881_),
    .ZN(_02882_));
 OAI21_X2 _11929_ (.A(_02646_),
    .B1(_02882_),
    .B2(_02649_),
    .ZN(_02883_));
 XNOR2_X2 _11930_ (.A(_02645_),
    .B(_02883_),
    .ZN(_02884_));
 AND2_X4 _11931_ (.A1(_02884_),
    .A2(_02874_),
    .ZN(_02885_));
 AND4_X4 _11932_ (.A1(_02697_),
    .A2(_02685_),
    .A3(_02709_),
    .A4(_02731_),
    .ZN(_02886_));
 BUF_X2 clone12 (.A(_03988_),
    .Z(net12));
 AND4_X4 _11934_ (.A1(_02767_),
    .A2(_02775_),
    .A3(_02781_),
    .A4(_02793_),
    .ZN(_02888_));
 NAND2_X4 _11935_ (.A1(_02888_),
    .A2(_02886_),
    .ZN(_02889_));
 AOI22_X4 _11936_ (.A1(_02867_),
    .A2(_02874_),
    .B1(_02885_),
    .B2(net13),
    .ZN(_02890_));
 XOR2_X2 _11937_ (.A(_02645_),
    .B(_02883_),
    .Z(_02891_));
 AOI21_X4 _11938_ (.A(_02891_),
    .B1(_02888_),
    .B2(_02886_),
    .ZN(_02892_));
 OAI21_X2 _11939_ (.A(_02797_),
    .B1(_01091_),
    .B2(_02873_),
    .ZN(_02893_));
 OR3_X4 _11940_ (.A1(_02892_),
    .A2(_02867_),
    .A3(_02893_),
    .ZN(_02894_));
 AOI21_X1 _11941_ (.A(_02859_),
    .B1(_02890_),
    .B2(_02894_),
    .ZN(_02895_));
 BUF_X1 _11942_ (.A(_09091_),
    .Z(_02896_));
 NAND3_X2 _11943_ (.A1(_09088_),
    .A2(_02896_),
    .A3(_02872_),
    .ZN(_02897_));
 OR2_X1 _11944_ (.A1(_02868_),
    .A2(_02897_),
    .ZN(_02898_));
 OR3_X2 _11945_ (.A1(net27),
    .A2(_02794_),
    .A3(_09080_),
    .ZN(_02899_));
 OAI21_X4 _11946_ (.A(_02884_),
    .B1(_02794_),
    .B2(_02732_),
    .ZN(_02900_));
 AOI21_X1 _11947_ (.A(_02898_),
    .B1(_02899_),
    .B2(_02900_),
    .ZN(_02901_));
 OR2_X2 _11948_ (.A1(_01091_),
    .A2(_02897_),
    .ZN(_02902_));
 NOR3_X1 _11949_ (.A1(_02892_),
    .A2(_02867_),
    .A3(_02902_),
    .ZN(_02903_));
 INV_X1 _11950_ (.A(_09096_),
    .ZN(_02904_));
 BUF_X2 _11951_ (.A(_09100_),
    .Z(_02905_));
 AOI21_X1 _11952_ (.A(_09099_),
    .B1(_09102_),
    .B2(_02905_),
    .ZN(_02906_));
 INV_X1 _11953_ (.A(_09097_),
    .ZN(_02907_));
 OAI21_X1 _11954_ (.A(_02904_),
    .B1(_02906_),
    .B2(_02907_),
    .ZN(_02908_));
 BUF_X4 _11955_ (.A(_09094_),
    .Z(_02909_));
 AOI21_X2 _11956_ (.A(_09093_),
    .B1(_02908_),
    .B2(_02909_),
    .ZN(_02910_));
 INV_X1 _11957_ (.A(_02910_),
    .ZN(_02911_));
 BUF_X4 _11958_ (.A(_09103_),
    .Z(_02912_));
 NAND4_X4 _11959_ (.A1(_09097_),
    .A2(_02909_),
    .A3(_02912_),
    .A4(_02905_),
    .ZN(_02913_));
 INV_X1 _11960_ (.A(_02757_),
    .ZN(_02914_));
 AOI211_X2 _11961_ (.A(_02914_),
    .B(_02814_),
    .C1(_02888_),
    .C2(_02886_),
    .ZN(_02915_));
 NOR2_X1 _11962_ (.A1(_02757_),
    .A2(_02814_),
    .ZN(_02916_));
 AND3_X2 _11963_ (.A1(_02886_),
    .A2(_02888_),
    .A3(_02916_),
    .ZN(_02917_));
 NOR3_X2 _11964_ (.A1(_02913_),
    .A2(_02915_),
    .A3(_02917_),
    .ZN(_02918_));
 OAI22_X2 _11965_ (.A1(_02901_),
    .A2(_02903_),
    .B1(_02911_),
    .B2(_02918_),
    .ZN(_02919_));
 BUF_X4 _11966_ (.A(_02919_),
    .Z(_02920_));
 AOI21_X2 _11967_ (.A(_02843_),
    .B1(_02895_),
    .B2(_02920_),
    .ZN(_02921_));
 OR3_X1 _11968_ (.A1(_02913_),
    .A2(_02915_),
    .A3(_02917_),
    .ZN(_02922_));
 OAI21_X1 _11969_ (.A(_01091_),
    .B1(_02892_),
    .B2(_02867_),
    .ZN(_02923_));
 NAND3_X1 _11970_ (.A1(_02868_),
    .A2(_02900_),
    .A3(_02899_),
    .ZN(_02924_));
 AOI221_X2 _11971_ (.A(_02897_),
    .B1(_02910_),
    .B2(_02922_),
    .C1(_02923_),
    .C2(_02924_),
    .ZN(_02925_));
 BUF_X4 _11972_ (.A(_02925_),
    .Z(_02926_));
 AND2_X4 _11973_ (.A1(_02890_),
    .A2(_02894_),
    .ZN(_02927_));
 BUF_X16 _11974_ (.A(_02927_),
    .Z(_02928_));
 AND2_X1 _11975_ (.A1(_02841_),
    .A2(_02643_),
    .ZN(_02929_));
 AOI22_X4 _11976_ (.A1(_02795_),
    .A2(_02858_),
    .B1(_02857_),
    .B2(_02929_),
    .ZN(_02930_));
 NOR3_X2 _11977_ (.A1(_02926_),
    .A2(_02928_),
    .A3(_02930_),
    .ZN(_02931_));
 NOR2_X2 _11978_ (.A1(_02686_),
    .A2(_02690_),
    .ZN(_02932_));
 NAND3_X2 _11979_ (.A1(_02729_),
    .A2(_02601_),
    .A3(_02716_),
    .ZN(_02933_));
 NOR3_X2 _11980_ (.A1(_02932_),
    .A2(_02728_),
    .A3(_02933_),
    .ZN(_02934_));
 NAND2_X1 _11981_ (.A1(_02518_),
    .A2(_02611_),
    .ZN(_02935_));
 OAI21_X2 _11982_ (.A(_02714_),
    .B1(_02935_),
    .B2(_02710_),
    .ZN(_02936_));
 AND2_X1 _11983_ (.A1(_02713_),
    .A2(_02936_),
    .ZN(_02937_));
 NAND2_X1 _11984_ (.A1(_02934_),
    .A2(_02937_),
    .ZN(_02938_));
 OAI21_X2 _11985_ (.A(_02938_),
    .B1(_02936_),
    .B2(_02713_),
    .ZN(_02939_));
 XNOR2_X1 _11986_ (.A(_01091_),
    .B(_02354_),
    .ZN(_02940_));
 OAI21_X2 _11987_ (.A(_02719_),
    .B1(_02940_),
    .B2(_02369_),
    .ZN(_02941_));
 AOI22_X4 _11988_ (.A1(_02698_),
    .A2(_02594_),
    .B1(_02481_),
    .B2(_02941_),
    .ZN(_02942_));
 NAND2_X1 _11989_ (.A1(_02942_),
    .A2(_02726_),
    .ZN(_02943_));
 AOI21_X2 _11990_ (.A(_02583_),
    .B1(_02943_),
    .B2(_02641_),
    .ZN(_02944_));
 NAND4_X4 _11991_ (.A1(_02832_),
    .A2(_02835_),
    .A3(_02840_),
    .A4(_02944_),
    .ZN(_02945_));
 NAND2_X2 _11992_ (.A1(_02715_),
    .A2(_02605_),
    .ZN(_02946_));
 NAND3_X1 _11993_ (.A1(_02589_),
    .A2(_02601_),
    .A3(_02605_),
    .ZN(_02947_));
 OAI21_X1 _11994_ (.A(_02589_),
    .B1(_02599_),
    .B2(_02600_),
    .ZN(_02948_));
 MUX2_X2 _11995_ (.A(_02947_),
    .B(_02948_),
    .S(_02729_),
    .Z(_02949_));
 AOI21_X2 _11996_ (.A(_02946_),
    .B1(_02949_),
    .B2(net18),
    .ZN(_02950_));
 NAND2_X1 _11997_ (.A1(_02937_),
    .A2(_02950_),
    .ZN(_02951_));
 OAI22_X2 _11998_ (.A1(net27),
    .A2(_02794_),
    .B1(_02945_),
    .B2(_02951_),
    .ZN(_02952_));
 OR2_X1 _11999_ (.A1(_02934_),
    .A2(_02936_),
    .ZN(_02953_));
 AND4_X2 _12000_ (.A1(_02832_),
    .A2(_02835_),
    .A3(_02840_),
    .A4(_02944_),
    .ZN(_02954_));
 AOI21_X2 _12001_ (.A(_02953_),
    .B1(_02950_),
    .B2(_02954_),
    .ZN(_02955_));
 NOR3_X4 _12002_ (.A1(_02939_),
    .A2(_02952_),
    .A3(_02955_),
    .ZN(_02956_));
 INV_X1 _12003_ (.A(_02781_),
    .ZN(_02957_));
 NAND3_X2 _12004_ (.A1(_02713_),
    .A2(_02714_),
    .A3(_02716_),
    .ZN(_02958_));
 AOI21_X4 _12005_ (.A(_02958_),
    .B1(_02949_),
    .B2(_02641_),
    .ZN(_02959_));
 AND2_X1 _12006_ (.A1(_02775_),
    .A2(_02959_),
    .ZN(_02960_));
 AOI21_X2 _12007_ (.A(_02957_),
    .B1(_02954_),
    .B2(_02960_),
    .ZN(_02961_));
 XNOR2_X2 _12008_ (.A(net27),
    .B(_02775_),
    .ZN(_02962_));
 AOI21_X4 _12009_ (.A(_02795_),
    .B1(_02961_),
    .B2(_02962_),
    .ZN(_02963_));
 XOR2_X2 _12010_ (.A(_02728_),
    .B(_02933_),
    .Z(_02964_));
 AOI21_X2 _12011_ (.A(_02739_),
    .B1(_02618_),
    .B2(_02761_),
    .ZN(_02965_));
 XNOR2_X2 _12012_ (.A(_02770_),
    .B(_02965_),
    .ZN(_02966_));
 OR2_X1 _12013_ (.A1(_02946_),
    .A2(_02966_),
    .ZN(_02967_));
 AOI211_X2 _12014_ (.A(_02945_),
    .B(_02967_),
    .C1(_02886_),
    .C2(_02888_),
    .ZN(_02968_));
 AND2_X1 _12015_ (.A1(_02806_),
    .A2(_02815_),
    .ZN(_02969_));
 NAND2_X1 _12016_ (.A1(_02645_),
    .A2(_02648_),
    .ZN(_02970_));
 NOR4_X1 _12017_ (.A1(_02435_),
    .A2(_09007_),
    .A3(_02970_),
    .A4(_02880_),
    .ZN(_02971_));
 AND2_X1 _12018_ (.A1(_02969_),
    .A2(_02971_),
    .ZN(_02972_));
 OAI211_X2 _12019_ (.A(_02942_),
    .B(_02972_),
    .C1(_02545_),
    .C2(_02582_),
    .ZN(_02973_));
 OAI21_X1 _12020_ (.A(_02726_),
    .B1(_02707_),
    .B2(_02699_),
    .ZN(_02974_));
 AOI221_X2 _12021_ (.A(_02973_),
    .B1(_02974_),
    .B2(_02641_),
    .C1(_02699_),
    .C2(_02834_),
    .ZN(_02975_));
 NOR3_X2 _12022_ (.A1(_02868_),
    .A2(_02831_),
    .A3(_02829_),
    .ZN(_02976_));
 AOI21_X2 _12023_ (.A(_01091_),
    .B1(_02845_),
    .B2(_02847_),
    .ZN(_02977_));
 OAI211_X4 _12024_ (.A(_02959_),
    .B(_02975_),
    .C1(_02976_),
    .C2(_02977_),
    .ZN(_02978_));
 AND3_X1 _12025_ (.A1(_02767_),
    .A2(_02775_),
    .A3(_02781_),
    .ZN(_02979_));
 AND3_X1 _12026_ (.A1(net380),
    .A2(_02731_),
    .A3(_02793_),
    .ZN(_02980_));
 AND3_X1 _12027_ (.A1(_02978_),
    .A2(_02979_),
    .A3(_02980_),
    .ZN(_02981_));
 XNOR2_X1 _12028_ (.A(_02713_),
    .B(_02934_),
    .ZN(_02982_));
 AND3_X2 _12029_ (.A1(_02685_),
    .A2(_02697_),
    .A3(_02709_),
    .ZN(_02983_));
 AND3_X1 _12030_ (.A1(_02716_),
    .A2(_02727_),
    .A3(_02730_),
    .ZN(_02984_));
 AOI21_X2 _12031_ (.A(_02982_),
    .B1(_02983_),
    .B2(_02984_),
    .ZN(_02985_));
 AND3_X1 _12032_ (.A1(_02982_),
    .A2(_02983_),
    .A3(_02984_),
    .ZN(_02986_));
 OAI33_X1 _12033_ (.A1(_02932_),
    .A2(_02964_),
    .A3(_02968_),
    .B1(_02981_),
    .B2(_02985_),
    .B3(_02986_),
    .ZN(_02987_));
 NAND2_X1 _12034_ (.A1(_02775_),
    .A2(_02781_),
    .ZN(_02988_));
 OR2_X1 _12035_ (.A1(_02732_),
    .A2(_02988_),
    .ZN(_02989_));
 AOI211_X2 _12036_ (.A(net27),
    .B(_02988_),
    .C1(_02793_),
    .C2(_02978_),
    .ZN(_02990_));
 MUX2_X2 _12037_ (.A(_02989_),
    .B(_02990_),
    .S(_02767_),
    .Z(_02991_));
 NOR4_X4 _12038_ (.A1(_02956_),
    .A2(_02963_),
    .A3(net378),
    .A4(_02991_),
    .ZN(_02992_));
 AOI21_X1 _12039_ (.A(_02765_),
    .B1(_02729_),
    .B2(_02618_),
    .ZN(_02993_));
 NOR2_X1 _12040_ (.A1(_02477_),
    .A2(_02993_),
    .ZN(_02994_));
 XOR2_X2 _12041_ (.A(_02762_),
    .B(_02790_),
    .Z(_02995_));
 AND2_X1 _12042_ (.A1(_02886_),
    .A2(_02979_),
    .ZN(_02996_));
 AOI221_X2 _12043_ (.A(_02425_),
    .B1(_02785_),
    .B2(_02994_),
    .C1(_02995_),
    .C2(_02996_),
    .ZN(_02997_));
 NAND4_X1 _12044_ (.A1(_02767_),
    .A2(_02775_),
    .A3(_02781_),
    .A4(_02959_),
    .ZN(_02998_));
 AOI211_X2 _12045_ (.A(_02945_),
    .B(_02998_),
    .C1(_02886_),
    .C2(_02888_),
    .ZN(_02999_));
 XNOR2_X2 _12046_ (.A(_02995_),
    .B(_02999_),
    .ZN(_03000_));
 INV_X1 _12047_ (.A(_02969_),
    .ZN(_03001_));
 NAND2_X1 _12048_ (.A1(net35),
    .A2(_02742_),
    .ZN(_03002_));
 XOR2_X2 _12049_ (.A(_02802_),
    .B(_03002_),
    .Z(_03003_));
 OR4_X4 _12050_ (.A1(_02913_),
    .A2(_01097_),
    .A3(_03001_),
    .A4(_03003_),
    .ZN(_03004_));
 OR2_X4 _12051_ (.A1(_02898_),
    .A2(_03004_),
    .ZN(_03005_));
 AOI21_X4 _12052_ (.A(_03005_),
    .B1(_02899_),
    .B2(_02900_),
    .ZN(_03006_));
 NOR4_X4 _12053_ (.A1(_03004_),
    .A2(_02867_),
    .A3(_02892_),
    .A4(_02902_),
    .ZN(_03007_));
 NOR4_X4 _12054_ (.A1(_03006_),
    .A2(_03000_),
    .A3(_02997_),
    .A4(_03007_),
    .ZN(_03008_));
 OAI21_X1 _12055_ (.A(_02729_),
    .B1(_02686_),
    .B2(_02763_),
    .ZN(_03009_));
 OAI21_X2 _12056_ (.A(_03009_),
    .B1(_02584_),
    .B2(_02942_),
    .ZN(_03010_));
 NAND4_X1 _12057_ (.A1(_02770_),
    .A2(_02685_),
    .A3(_02697_),
    .A4(_02709_),
    .ZN(_03011_));
 AOI21_X2 _12058_ (.A(_03010_),
    .B1(_03011_),
    .B2(_02946_),
    .ZN(_03012_));
 NAND3_X4 _12059_ (.A1(_02978_),
    .A2(_02979_),
    .A3(_02980_),
    .ZN(_03013_));
 AOI21_X4 _12060_ (.A(_03012_),
    .B1(_02983_),
    .B2(_03013_),
    .ZN(_03014_));
 OAI21_X2 _12061_ (.A(_02954_),
    .B1(_02794_),
    .B2(net27),
    .ZN(_03015_));
 XNOR2_X2 _12062_ (.A(_03015_),
    .B(_02966_),
    .ZN(_03016_));
 NOR3_X4 _12063_ (.A1(_03014_),
    .A2(_02930_),
    .A3(_03016_),
    .ZN(_03017_));
 NAND3_X4 _12064_ (.A1(_02992_),
    .A2(_03008_),
    .A3(_03017_),
    .ZN(_03018_));
 BUF_X4 _12065_ (.A(_03018_),
    .Z(_03019_));
 AOI21_X4 _12066_ (.A(_02921_),
    .B1(_02931_),
    .B2(_03019_),
    .ZN(_03020_));
 INV_X1 _12067_ (.A(_09109_),
    .ZN(_03021_));
 INV_X1 _12068_ (.A(_09114_),
    .ZN(_03022_));
 AOI21_X2 _12069_ (.A(_09120_),
    .B1(_09123_),
    .B2(_09121_),
    .ZN(_03023_));
 OAI21_X1 _12070_ (.A(_09124_),
    .B1(_09125_),
    .B2(_09126_),
    .ZN(_03024_));
 INV_X1 _12071_ (.A(_09121_),
    .ZN(_03025_));
 OAI21_X4 _12072_ (.A(_03023_),
    .B1(_03024_),
    .B2(_03025_),
    .ZN(_03026_));
 AOI21_X4 _12073_ (.A(_09117_),
    .B1(_03026_),
    .B2(_09118_),
    .ZN(_03027_));
 INV_X1 _12074_ (.A(_09115_),
    .ZN(_03028_));
 OAI21_X4 _12075_ (.A(_03022_),
    .B1(_03027_),
    .B2(_03028_),
    .ZN(_03029_));
 AOI21_X4 _12076_ (.A(_09111_),
    .B1(_03029_),
    .B2(_09112_),
    .ZN(_03030_));
 NOR2_X4 _12077_ (.A1(_03030_),
    .A2(_03021_),
    .ZN(_03031_));
 NOR2_X4 _12078_ (.A1(_09108_),
    .A2(_03031_),
    .ZN(_03032_));
 NOR2_X2 _12079_ (.A1(_02915_),
    .A2(_02917_),
    .ZN(_03033_));
 NAND2_X4 _12080_ (.A1(_02894_),
    .A2(_02890_),
    .ZN(_03034_));
 NAND2_X1 _12081_ (.A1(_02920_),
    .A2(_03034_),
    .ZN(_03035_));
 BUF_X4 _12082_ (.A(_03035_),
    .Z(_03036_));
 NOR2_X1 _12083_ (.A1(_09114_),
    .A2(_09125_),
    .ZN(_03037_));
 INV_X1 _12084_ (.A(_03023_),
    .ZN(_03038_));
 AOI21_X1 _12085_ (.A(_09117_),
    .B1(_03038_),
    .B2(_09118_),
    .ZN(_03039_));
 OAI21_X1 _12086_ (.A(_03037_),
    .B1(_03039_),
    .B2(_03028_),
    .ZN(_03040_));
 AND2_X1 _12087_ (.A1(_09109_),
    .A2(_09111_),
    .ZN(_03041_));
 OR3_X2 _12088_ (.A1(_09108_),
    .A2(_03040_),
    .A3(_03041_),
    .ZN(_03042_));
 NOR4_X4 _12089_ (.A1(_03033_),
    .A2(_03036_),
    .A3(_03019_),
    .A4(_03042_),
    .ZN(_03043_));
 NOR3_X1 _12090_ (.A1(_02914_),
    .A2(net13),
    .A3(_03003_),
    .ZN(_03044_));
 OR3_X1 _12091_ (.A1(_02809_),
    .A2(_02811_),
    .A3(_02813_),
    .ZN(_03045_));
 NOR3_X1 _12092_ (.A1(_02757_),
    .A2(_02795_),
    .A3(_03045_),
    .ZN(_03046_));
 OAI21_X1 _12093_ (.A(_01710_),
    .B1(_03044_),
    .B2(_03046_),
    .ZN(_03047_));
 NAND2_X4 _12094_ (.A1(_02889_),
    .A2(_02916_),
    .ZN(_03048_));
 NAND2_X1 _12095_ (.A1(_02969_),
    .A2(_03048_),
    .ZN(_03049_));
 OR3_X1 _12096_ (.A1(_03042_),
    .A2(_03047_),
    .A3(_03049_),
    .ZN(_03050_));
 AND3_X4 _12097_ (.A1(_02992_),
    .A2(_03017_),
    .A3(_03008_),
    .ZN(_03051_));
 BUF_X8 _12098_ (.A(_03051_),
    .Z(_03052_));
 NOR2_X4 _12099_ (.A1(_02928_),
    .A2(_02926_),
    .ZN(_03053_));
 BUF_X8 _12100_ (.A(_03053_),
    .Z(_03054_));
 AOI21_X2 _12101_ (.A(_03050_),
    .B1(net41),
    .B2(_03054_),
    .ZN(_03055_));
 NOR3_X4 _12102_ (.A1(_03032_),
    .A2(_03043_),
    .A3(_03055_),
    .ZN(_03056_));
 NAND2_X4 _12103_ (.A1(_02900_),
    .A2(_02899_),
    .ZN(_03057_));
 INV_X1 _12104_ (.A(_09105_),
    .ZN(_03058_));
 INV_X1 _12105_ (.A(_02896_),
    .ZN(_03059_));
 AOI21_X1 _12106_ (.A(_03059_),
    .B1(_02913_),
    .B2(_02910_),
    .ZN(_03060_));
 OR2_X1 _12107_ (.A1(_09090_),
    .A2(_03060_),
    .ZN(_03061_));
 AND2_X1 _12108_ (.A1(_09088_),
    .A2(_03061_),
    .ZN(_03062_));
 OAI21_X1 _12109_ (.A(_02872_),
    .B1(_09087_),
    .B2(_03062_),
    .ZN(_03063_));
 AND2_X1 _12110_ (.A1(_03058_),
    .A2(_03063_),
    .ZN(_03064_));
 INV_X1 _12111_ (.A(_03064_),
    .ZN(_03065_));
 NAND2_X1 _12112_ (.A1(_02868_),
    .A2(_03065_),
    .ZN(_03066_));
 NAND2_X1 _12113_ (.A1(_09088_),
    .A2(_03061_),
    .ZN(_03067_));
 NOR4_X2 _12114_ (.A1(_02872_),
    .A2(_02915_),
    .A3(_02917_),
    .A4(_03067_),
    .ZN(_03068_));
 NOR2_X1 _12115_ (.A1(_02872_),
    .A2(_09087_),
    .ZN(_03069_));
 AOI21_X1 _12116_ (.A(_09093_),
    .B1(_09096_),
    .B2(_02909_),
    .ZN(_03070_));
 INV_X1 _12117_ (.A(_03070_),
    .ZN(_03071_));
 AOI21_X1 _12118_ (.A(_09090_),
    .B1(_03071_),
    .B2(_02896_),
    .ZN(_03072_));
 INV_X1 _12119_ (.A(_09088_),
    .ZN(_03073_));
 OAI21_X1 _12120_ (.A(_02906_),
    .B1(_03072_),
    .B2(_03073_),
    .ZN(_03074_));
 INV_X1 _12121_ (.A(_03074_),
    .ZN(_03075_));
 OAI21_X1 _12122_ (.A(_03069_),
    .B1(_03075_),
    .B2(_03067_),
    .ZN(_03076_));
 INV_X1 _12123_ (.A(_02872_),
    .ZN(_03077_));
 NOR3_X1 _12124_ (.A1(_03077_),
    .A2(_09087_),
    .A3(_03074_),
    .ZN(_03078_));
 OR2_X1 _12125_ (.A1(_02915_),
    .A2(_02917_),
    .ZN(_03079_));
 AOI221_X1 _12126_ (.A(_03068_),
    .B1(_03076_),
    .B2(_03063_),
    .C1(_03078_),
    .C2(_03079_),
    .ZN(_03080_));
 CLKBUF_X3 _12127_ (.A(_03080_),
    .Z(_03081_));
 NOR3_X2 _12128_ (.A1(_03057_),
    .A2(_03066_),
    .A3(_03081_),
    .ZN(_03082_));
 BUF_X2 _12129_ (.A(_02868_),
    .Z(_03083_));
 NOR3_X1 _12130_ (.A1(_03083_),
    .A2(_03057_),
    .A3(_03065_),
    .ZN(_03084_));
 AOI221_X2 _12131_ (.A(_03082_),
    .B1(_03084_),
    .B2(_03081_),
    .C1(_03052_),
    .C2(net424),
    .ZN(_03085_));
 OR2_X1 _12132_ (.A1(_02803_),
    .A2(_02308_),
    .ZN(_08981_));
 XNOR2_X1 _12133_ (.A(_01142_),
    .B(_02751_),
    .ZN(_03086_));
 MUX2_X1 _12134_ (.A(_08981_),
    .B(_03086_),
    .S(_02344_),
    .Z(_08989_));
 OR3_X1 _12135_ (.A1(_08985_),
    .A2(_08991_),
    .A3(_08984_),
    .ZN(_03087_));
 AND2_X1 _12136_ (.A1(_01126_),
    .A2(_03087_),
    .ZN(_03088_));
 MUX2_X1 _12137_ (.A(_08989_),
    .B(_03088_),
    .S(_02347_),
    .Z(_09022_));
 XNOR2_X1 _12138_ (.A(_09024_),
    .B(_02313_),
    .ZN(_03089_));
 MUX2_X1 _12139_ (.A(_09022_),
    .B(_03089_),
    .S(_02585_),
    .Z(_09042_));
 OR3_X1 _12140_ (.A1(_09044_),
    .A2(_09028_),
    .A3(_02362_),
    .ZN(_03090_));
 AND2_X1 _12141_ (.A1(_02363_),
    .A2(_03090_),
    .ZN(_03091_));
 MUX2_X1 _12142_ (.A(_09042_),
    .B(_03091_),
    .S(_02698_),
    .Z(_09063_));
 XOR2_X1 _12143_ (.A(_09065_),
    .B(_02557_),
    .Z(_03092_));
 MUX2_X1 _12144_ (.A(_09063_),
    .B(_03092_),
    .S(_02642_),
    .Z(_09083_));
 OR3_X2 _12145_ (.A1(_02732_),
    .A2(_02794_),
    .A3(_09083_),
    .ZN(_03093_));
 NOR2_X1 _12146_ (.A1(_02822_),
    .A2(_02825_),
    .ZN(_03094_));
 XNOR2_X2 _12147_ (.A(_02648_),
    .B(_03094_),
    .ZN(_03095_));
 OAI21_X4 _12148_ (.A(_03093_),
    .B1(_03095_),
    .B2(_02795_),
    .ZN(_03096_));
 XNOR2_X1 _12149_ (.A(_01091_),
    .B(_03096_),
    .ZN(_03097_));
 AOI21_X1 _12150_ (.A(_03082_),
    .B1(_03097_),
    .B2(_03057_),
    .ZN(_03098_));
 NOR2_X1 _12151_ (.A1(_03035_),
    .A2(_03018_),
    .ZN(_03099_));
 BUF_X4 _12152_ (.A(_03099_),
    .Z(_03100_));
 AOI21_X2 _12153_ (.A(_03085_),
    .B1(_03098_),
    .B2(_03100_),
    .ZN(_03101_));
 CLKBUF_X3 _12154_ (.A(_03083_),
    .Z(_03102_));
 AOI21_X1 _12155_ (.A(_03068_),
    .B1(_03078_),
    .B2(_03079_),
    .ZN(_03103_));
 NAND2_X1 _12156_ (.A1(_03063_),
    .A2(_03076_),
    .ZN(_03104_));
 NAND2_X2 _12157_ (.A1(_03103_),
    .A2(_03104_),
    .ZN(_03105_));
 NAND2_X1 _12158_ (.A1(_03057_),
    .A2(_03065_),
    .ZN(_03106_));
 NAND3_X1 _12159_ (.A1(_03083_),
    .A2(_03057_),
    .A3(_03064_),
    .ZN(_03107_));
 OAI21_X1 _12160_ (.A(_03062_),
    .B1(_03074_),
    .B2(_03033_),
    .ZN(_03108_));
 AND2_X1 _12161_ (.A1(_03069_),
    .A2(_03108_),
    .ZN(_03109_));
 OAI33_X1 _12162_ (.A1(_03102_),
    .A2(_03105_),
    .A3(_03106_),
    .B1(_03107_),
    .B2(_03109_),
    .B3(_03100_),
    .ZN(_03110_));
 OAI21_X4 _12163_ (.A(_03056_),
    .B1(_03101_),
    .B2(_03110_),
    .ZN(_03111_));
 NAND2_X4 _12164_ (.A1(_03054_),
    .A2(_03052_),
    .ZN(_03112_));
 INV_X1 _12165_ (.A(_02859_),
    .ZN(_03113_));
 OAI21_X2 _12166_ (.A(_03113_),
    .B1(net425),
    .B2(_02926_),
    .ZN(_03114_));
 OAI21_X1 _12167_ (.A(_02855_),
    .B1(_02854_),
    .B2(_02853_),
    .ZN(_03115_));
 NAND2_X1 _12168_ (.A1(net13),
    .A2(_02856_),
    .ZN(_03116_));
 NAND2_X1 _12169_ (.A1(_03115_),
    .A2(_03116_),
    .ZN(_03117_));
 INV_X1 _12170_ (.A(_02850_),
    .ZN(_03118_));
 MUX2_X1 _12171_ (.A(_03118_),
    .B(_02858_),
    .S(_02795_),
    .Z(_03119_));
 OR4_X2 _12172_ (.A1(_02926_),
    .A2(_02928_),
    .A3(_03117_),
    .A4(_03119_),
    .ZN(_03120_));
 AND3_X2 _12173_ (.A1(_03112_),
    .A2(_03114_),
    .A3(_03120_),
    .ZN(_03121_));
 XNOR2_X2 _12174_ (.A(_01091_),
    .B(_03064_),
    .ZN(_03122_));
 NOR2_X1 _12175_ (.A1(_03057_),
    .A2(_03122_),
    .ZN(_03123_));
 NOR4_X1 _12176_ (.A1(_02894_),
    .A2(_03014_),
    .A3(_02930_),
    .A4(_03016_),
    .ZN(_03124_));
 AND4_X1 _12177_ (.A1(_02992_),
    .A2(_03008_),
    .A3(_02920_),
    .A4(_03124_),
    .ZN(_03125_));
 NOR2_X2 _12178_ (.A1(_03123_),
    .A2(_03125_),
    .ZN(_03126_));
 NAND2_X2 _12179_ (.A1(_03057_),
    .A2(_03122_),
    .ZN(_03127_));
 NAND2_X1 _12180_ (.A1(_02992_),
    .A2(_03008_),
    .ZN(_03128_));
 NAND4_X1 _12181_ (.A1(_02920_),
    .A2(_03034_),
    .A3(_03017_),
    .A4(_03096_),
    .ZN(_03129_));
 OAI21_X1 _12182_ (.A(_02573_),
    .B1(_03128_),
    .B2(_03129_),
    .ZN(_03130_));
 AOI21_X1 _12183_ (.A(_03105_),
    .B1(_03051_),
    .B2(_03054_),
    .ZN(_03131_));
 OAI221_X1 _12184_ (.A(_03126_),
    .B1(_03127_),
    .B2(_03099_),
    .C1(_03130_),
    .C2(_03131_),
    .ZN(_03132_));
 CLKBUF_X3 _12185_ (.A(_03132_),
    .Z(_03133_));
 NOR2_X2 _12186_ (.A1(_03121_),
    .A2(_03133_),
    .ZN(_03134_));
 OAI211_X4 _12187_ (.A(_03114_),
    .B(_03120_),
    .C1(_03036_),
    .C2(_03019_),
    .ZN(_03135_));
 OR2_X1 _12188_ (.A1(_02844_),
    .A2(_02856_),
    .ZN(_03136_));
 NAND2_X1 _12189_ (.A1(_02841_),
    .A2(_02643_),
    .ZN(_03137_));
 OAI33_X1 _12190_ (.A1(_02848_),
    .A2(net13),
    .A3(_02855_),
    .B1(_02850_),
    .B2(_03136_),
    .B3(_03137_),
    .ZN(_03138_));
 AOI21_X2 _12191_ (.A(_03010_),
    .B1(_02983_),
    .B2(_03013_),
    .ZN(_03139_));
 AND3_X1 _12192_ (.A1(_03013_),
    .A2(_02983_),
    .A3(_03010_),
    .ZN(_03140_));
 OAI21_X2 _12193_ (.A(_03138_),
    .B1(_03139_),
    .B2(_03140_),
    .ZN(_03141_));
 AND2_X1 _12194_ (.A1(_03016_),
    .A2(_03141_),
    .ZN(_03142_));
 XOR2_X1 _12195_ (.A(_03015_),
    .B(_02966_),
    .Z(_03143_));
 AOI21_X1 _12196_ (.A(_03143_),
    .B1(_03034_),
    .B2(_02920_),
    .ZN(_03144_));
 NOR4_X1 _12197_ (.A1(_02926_),
    .A2(_02928_),
    .A3(_03016_),
    .A4(_03141_),
    .ZN(_03145_));
 AOI211_X2 _12198_ (.A(_03142_),
    .B(_03144_),
    .C1(_03145_),
    .C2(_03018_),
    .ZN(_03146_));
 NAND2_X1 _12199_ (.A1(_02797_),
    .A2(_03066_),
    .ZN(_03147_));
 NOR2_X1 _12200_ (.A1(_02868_),
    .A2(_03064_),
    .ZN(_03148_));
 MUX2_X2 _12201_ (.A(_03147_),
    .B(_03148_),
    .S(_03057_),
    .Z(_03149_));
 NOR2_X1 _12202_ (.A1(_02930_),
    .A2(_03149_),
    .ZN(_03150_));
 OR3_X4 _12203_ (.A1(_03139_),
    .A2(_03140_),
    .A3(_03150_),
    .ZN(_03151_));
 NAND4_X4 _12204_ (.A1(_03135_),
    .A2(_03146_),
    .A3(_03151_),
    .A4(_03020_),
    .ZN(_03152_));
 NOR2_X1 _12205_ (.A1(_02868_),
    .A2(_03032_),
    .ZN(_03153_));
 AND2_X2 _12206_ (.A1(_03081_),
    .A2(_03153_),
    .ZN(_03154_));
 OR2_X4 _12207_ (.A1(_03031_),
    .A2(_09108_),
    .ZN(_03155_));
 NAND2_X4 _12208_ (.A1(_03155_),
    .A2(_02868_),
    .ZN(_03156_));
 INV_X4 _12209_ (.A(_03156_),
    .ZN(_03157_));
 NOR2_X4 _12210_ (.A1(_03157_),
    .A2(_02573_),
    .ZN(_03158_));
 NOR2_X2 _12211_ (.A1(_03081_),
    .A2(_03158_),
    .ZN(_03159_));
 OAI22_X4 _12212_ (.A1(_03036_),
    .A2(_03018_),
    .B1(_03159_),
    .B2(_03154_),
    .ZN(_03160_));
 NOR2_X1 _12213_ (.A1(_03158_),
    .A2(_03096_),
    .ZN(_03161_));
 AND2_X1 _12214_ (.A1(_03096_),
    .A2(_03153_),
    .ZN(_03162_));
 OAI211_X2 _12215_ (.A(_03054_),
    .B(_03052_),
    .C1(_03162_),
    .C2(_03161_),
    .ZN(_03163_));
 NAND2_X4 _12216_ (.A1(_03163_),
    .A2(_03160_),
    .ZN(_03164_));
 NOR3_X2 _12217_ (.A1(_02932_),
    .A2(_02964_),
    .A3(_02968_),
    .ZN(_03165_));
 INV_X1 _12218_ (.A(_02950_),
    .ZN(_03166_));
 NOR2_X1 _12219_ (.A1(_03015_),
    .A2(_03166_),
    .ZN(_03167_));
 NOR2_X2 _12220_ (.A1(_03165_),
    .A2(_03167_),
    .ZN(_03168_));
 NOR2_X1 _12221_ (.A1(_02920_),
    .A2(_03168_),
    .ZN(_03169_));
 AOI21_X1 _12222_ (.A(_03168_),
    .B1(_03017_),
    .B2(_03034_),
    .ZN(_03170_));
 OR2_X1 _12223_ (.A1(_03165_),
    .A2(_03167_),
    .ZN(_03171_));
 AOI21_X1 _12224_ (.A(_03171_),
    .B1(_03008_),
    .B2(_02992_),
    .ZN(_03172_));
 AND3_X1 _12225_ (.A1(_02919_),
    .A2(_03034_),
    .A3(_03017_),
    .ZN(_03173_));
 AOI211_X4 _12226_ (.A(_03169_),
    .B(_03170_),
    .C1(_03172_),
    .C2(_03173_),
    .ZN(_03174_));
 NOR3_X4 _12227_ (.A1(_02981_),
    .A2(_02985_),
    .A3(_02986_),
    .ZN(_03175_));
 AOI21_X1 _12228_ (.A(_02573_),
    .B1(_02868_),
    .B2(_03065_),
    .ZN(_03176_));
 INV_X1 _12229_ (.A(_03148_),
    .ZN(_03177_));
 MUX2_X1 _12230_ (.A(_03176_),
    .B(_03177_),
    .S(_03057_),
    .Z(_03178_));
 NAND3_X2 _12231_ (.A1(_03017_),
    .A2(_03178_),
    .A3(_03168_),
    .ZN(_03179_));
 NOR4_X4 _12232_ (.A1(_02987_),
    .A2(_03014_),
    .A3(_02930_),
    .A4(_03016_),
    .ZN(_03180_));
 NAND3_X2 _12233_ (.A1(_02920_),
    .A2(_03034_),
    .A3(_03180_),
    .ZN(_03181_));
 AOI22_X4 _12234_ (.A1(_03175_),
    .A2(_03179_),
    .B1(_03181_),
    .B2(_02956_),
    .ZN(_03182_));
 OR4_X2 _12235_ (.A1(_02987_),
    .A2(_03014_),
    .A3(_02930_),
    .A4(_03016_),
    .ZN(_03183_));
 NOR2_X2 _12236_ (.A1(_03149_),
    .A2(_03183_),
    .ZN(_03184_));
 OR3_X4 _12237_ (.A1(_02956_),
    .A2(_02963_),
    .A3(_02991_),
    .ZN(_03185_));
 OR2_X1 _12238_ (.A1(_02997_),
    .A2(_03000_),
    .ZN(_03186_));
 OR4_X2 _12239_ (.A1(_03185_),
    .A2(_03186_),
    .A3(_02926_),
    .A4(_02928_),
    .ZN(_03187_));
 AOI21_X2 _12240_ (.A(_02963_),
    .B1(_03184_),
    .B2(_03187_),
    .ZN(_03188_));
 OR2_X1 _12241_ (.A1(_02991_),
    .A2(_02997_),
    .ZN(_03189_));
 NAND4_X1 _12242_ (.A1(_02992_),
    .A2(_02920_),
    .A3(_03034_),
    .A4(_03017_),
    .ZN(_03190_));
 AOI21_X2 _12243_ (.A(_03189_),
    .B1(_03190_),
    .B2(_03000_),
    .ZN(_03191_));
 NAND4_X4 _12244_ (.A1(_03174_),
    .A2(_03182_),
    .A3(_03188_),
    .A4(_03191_),
    .ZN(_03192_));
 AOI22_X1 _12245_ (.A1(_02770_),
    .A2(_02965_),
    .B1(_02983_),
    .B2(_02727_),
    .ZN(_03193_));
 AND2_X1 _12246_ (.A1(_03013_),
    .A2(_02983_),
    .ZN(_03194_));
 OAI21_X1 _12247_ (.A(_02727_),
    .B1(_02965_),
    .B2(_03194_),
    .ZN(_03195_));
 INV_X1 _12248_ (.A(_03195_),
    .ZN(_03196_));
 MUX2_X1 _12249_ (.A(_03193_),
    .B(_03196_),
    .S(_02716_),
    .Z(_03197_));
 NOR3_X1 _12250_ (.A1(_03016_),
    .A2(_03141_),
    .A3(_03149_),
    .ZN(_03198_));
 OAI21_X1 _12251_ (.A(_03198_),
    .B1(_03018_),
    .B2(_03035_),
    .ZN(_03199_));
 XNOR2_X2 _12252_ (.A(_03197_),
    .B(_03199_),
    .ZN(_03200_));
 OAI21_X4 _12253_ (.A(_03126_),
    .B1(_03127_),
    .B2(_03100_),
    .ZN(_03201_));
 OR4_X4 _12254_ (.A1(_03164_),
    .A2(_03192_),
    .A3(_03200_),
    .A4(_03201_),
    .ZN(_03202_));
 OR4_X4 clone16 (.A1(_03192_),
    .A2(_03164_),
    .A3(_03200_),
    .A4(_03201_),
    .ZN(net16));
 OAI211_X2 _12256_ (.A(_03111_),
    .B(_03134_),
    .C1(_03152_),
    .C2(_03202_),
    .ZN(_03204_));
 XNOR2_X2 _12257_ (.A(_03020_),
    .B(_03204_),
    .ZN(_03205_));
 NAND2_X1 _12258_ (.A1(_02775_),
    .A2(_02959_),
    .ZN(_03206_));
 NOR2_X2 _12259_ (.A1(_02796_),
    .A2(_02962_),
    .ZN(_03207_));
 NAND2_X1 _12260_ (.A1(_03184_),
    .A2(_03187_),
    .ZN(_03208_));
 OAI33_X1 _12261_ (.A1(_02796_),
    .A2(_02945_),
    .A3(_03206_),
    .B1(_03207_),
    .B2(_03208_),
    .B3(_02956_),
    .ZN(_03209_));
 XNOR2_X2 _12262_ (.A(_02957_),
    .B(_03209_),
    .ZN(_03210_));
 NOR3_X4 _12263_ (.A1(_03152_),
    .A2(_03200_),
    .A3(_03133_),
    .ZN(_03211_));
 NAND2_X2 _12264_ (.A1(_03178_),
    .A2(_03180_),
    .ZN(_03212_));
 NOR4_X4 _12265_ (.A1(_03185_),
    .A2(_03186_),
    .A3(_02926_),
    .A4(net425),
    .ZN(_03213_));
 NOR3_X4 _12266_ (.A1(_02956_),
    .A2(_03212_),
    .A3(_03213_),
    .ZN(_03214_));
 XNOR2_X2 _12267_ (.A(_03207_),
    .B(_03214_),
    .ZN(_03215_));
 AND3_X1 _12268_ (.A1(_03174_),
    .A2(_03182_),
    .A3(_03215_),
    .ZN(_03216_));
 NAND4_X4 _12269_ (.A1(net16),
    .A2(_03111_),
    .A3(_03211_),
    .A4(_03216_),
    .ZN(_03217_));
 XNOR2_X2 _12270_ (.A(_03210_),
    .B(_03217_),
    .ZN(_03218_));
 NOR4_X2 _12271_ (.A1(_02956_),
    .A2(_02963_),
    .A3(_03212_),
    .A4(_03213_),
    .ZN(_03219_));
 XNOR2_X2 _12272_ (.A(_02991_),
    .B(_03219_),
    .ZN(_03220_));
 NAND3_X1 _12273_ (.A1(_03174_),
    .A2(_03182_),
    .A3(_03188_),
    .ZN(_03221_));
 NAND3_X4 _12274_ (.A1(_03146_),
    .A2(_03151_),
    .A3(_03020_),
    .ZN(_03222_));
 AND2_X1 _12275_ (.A1(_03155_),
    .A2(_03097_),
    .ZN(_03223_));
 NOR3_X1 _12276_ (.A1(_03036_),
    .A2(_03019_),
    .A3(_03223_),
    .ZN(_03224_));
 AOI221_X2 _12277_ (.A(_03154_),
    .B1(_03105_),
    .B2(_03157_),
    .C1(_03053_),
    .C2(_03051_),
    .ZN(_03225_));
 OAI21_X1 _12278_ (.A(_03135_),
    .B1(_03224_),
    .B2(_03225_),
    .ZN(_03226_));
 OR4_X2 _12279_ (.A1(_03222_),
    .A2(_03200_),
    .A3(_03133_),
    .A4(_03226_),
    .ZN(_03227_));
 NOR3_X1 _12280_ (.A1(_03191_),
    .A2(_03221_),
    .A3(_03227_),
    .ZN(_03228_));
 XOR2_X2 _12281_ (.A(_03220_),
    .B(_03228_),
    .Z(_03229_));
 XOR2_X2 _12282_ (.A(_02995_),
    .B(_02999_),
    .Z(_03230_));
 NOR4_X4 _12283_ (.A1(_03185_),
    .A2(_02926_),
    .A3(net425),
    .A4(_03183_),
    .ZN(_03231_));
 AOI21_X1 _12284_ (.A(_03000_),
    .B1(_02894_),
    .B2(_02890_),
    .ZN(_03232_));
 OAI21_X2 _12285_ (.A(_03232_),
    .B1(_03141_),
    .B2(_02920_),
    .ZN(_03233_));
 OAI211_X2 _12286_ (.A(_02992_),
    .B(_03017_),
    .C1(_02926_),
    .C2(_02997_),
    .ZN(_03234_));
 OAI22_X4 _12287_ (.A1(_03230_),
    .A2(_03231_),
    .B1(_03233_),
    .B2(_03234_),
    .ZN(_03235_));
 AND2_X1 _12288_ (.A1(_03083_),
    .A2(_03081_),
    .ZN(_03236_));
 NOR2_X1 _12289_ (.A1(_03083_),
    .A2(_03081_),
    .ZN(_03237_));
 OAI22_X2 _12290_ (.A1(_03036_),
    .A2(_03019_),
    .B1(_03236_),
    .B2(_03237_),
    .ZN(_03238_));
 NOR2_X1 _12291_ (.A1(_03083_),
    .A2(_03096_),
    .ZN(_03239_));
 INV_X1 _12292_ (.A(_03096_),
    .ZN(_09104_));
 NOR2_X1 _12293_ (.A1(_08819_),
    .A2(_09104_),
    .ZN(_03240_));
 OAI211_X2 _12294_ (.A(net424),
    .B(net41),
    .C1(_03239_),
    .C2(_03240_),
    .ZN(_03241_));
 AND2_X2 _12295_ (.A1(_03238_),
    .A2(_03241_),
    .ZN(_03242_));
 NAND2_X1 _12296_ (.A1(_03056_),
    .A2(_03242_),
    .ZN(_03243_));
 AND3_X1 _12297_ (.A1(_03174_),
    .A2(_03182_),
    .A3(_03188_),
    .ZN(_03244_));
 AND2_X1 _12298_ (.A1(_03244_),
    .A2(_03220_),
    .ZN(_03245_));
 NAND4_X2 _12299_ (.A1(_03202_),
    .A2(_03211_),
    .A3(_03243_),
    .A4(_03245_),
    .ZN(_03246_));
 XOR2_X2 _12300_ (.A(_03235_),
    .B(_03246_),
    .Z(_03247_));
 NAND4_X4 _12301_ (.A1(_03205_),
    .A2(_03218_),
    .A3(_03229_),
    .A4(_03247_),
    .ZN(_03248_));
 AOI21_X2 _12302_ (.A(_03119_),
    .B1(_03034_),
    .B2(_02920_),
    .ZN(_03249_));
 INV_X1 _12303_ (.A(_03119_),
    .ZN(_03250_));
 NOR3_X2 _12304_ (.A1(_02926_),
    .A2(net425),
    .A3(_03250_),
    .ZN(_03251_));
 AOI21_X4 _12305_ (.A(_03249_),
    .B1(_03251_),
    .B2(_03019_),
    .ZN(_03252_));
 AOI21_X1 _12306_ (.A(_03133_),
    .B1(_03242_),
    .B2(_03056_),
    .ZN(_03253_));
 OAI21_X1 _12307_ (.A(_03253_),
    .B1(net16),
    .B2(_03152_),
    .ZN(_03254_));
 XOR2_X2 _12308_ (.A(_03252_),
    .B(_03254_),
    .Z(_03255_));
 NAND2_X1 _12309_ (.A1(_02992_),
    .A2(_03017_),
    .ZN(_03256_));
 OAI21_X1 _12310_ (.A(_02997_),
    .B1(_03233_),
    .B2(_03256_),
    .ZN(_03257_));
 INV_X1 _12311_ (.A(_03257_),
    .ZN(_03258_));
 NAND3_X1 _12312_ (.A1(net424),
    .A2(net41),
    .A3(_03096_),
    .ZN(_03259_));
 OAI21_X1 _12313_ (.A(_03081_),
    .B1(_03019_),
    .B2(_03036_),
    .ZN(_03260_));
 AND4_X1 _12314_ (.A1(_09108_),
    .A2(_03083_),
    .A3(_03259_),
    .A4(_03260_),
    .ZN(_03261_));
 OR4_X2 _12315_ (.A1(_03152_),
    .A2(_03200_),
    .A3(_03133_),
    .A4(_03261_),
    .ZN(_03262_));
 AND2_X1 _12316_ (.A1(_09108_),
    .A2(_08819_),
    .ZN(_03263_));
 NAND2_X1 _12317_ (.A1(_03081_),
    .A2(_03263_),
    .ZN(_03264_));
 AOI21_X2 _12318_ (.A(_03264_),
    .B1(net41),
    .B2(net424),
    .ZN(_03265_));
 AND4_X1 _12319_ (.A1(net424),
    .A2(_03052_),
    .A3(_03096_),
    .A4(_03263_),
    .ZN(_03266_));
 NOR4_X2 _12320_ (.A1(_02991_),
    .A2(_03235_),
    .A3(_03265_),
    .A4(_03266_),
    .ZN(_03267_));
 NAND3_X1 _12321_ (.A1(_03031_),
    .A2(_03238_),
    .A3(_03241_),
    .ZN(_03268_));
 BUF_X4 _12322_ (.A(_03201_),
    .Z(_03269_));
 OAI211_X2 _12323_ (.A(_03244_),
    .B(_03267_),
    .C1(_03268_),
    .C2(_03269_),
    .ZN(_03270_));
 OAI21_X4 _12324_ (.A(_03258_),
    .B1(_03262_),
    .B2(_03270_),
    .ZN(_03271_));
 NOR2_X1 _12325_ (.A1(_03164_),
    .A2(_03269_),
    .ZN(_03272_));
 OR3_X2 _12326_ (.A1(_03032_),
    .A2(_03043_),
    .A3(_03055_),
    .ZN(_03273_));
 XNOR2_X2 _12327_ (.A(_03273_),
    .B(_03242_),
    .ZN(_03274_));
 AND2_X1 _12328_ (.A1(_03164_),
    .A2(_03269_),
    .ZN(_03275_));
 OR2_X1 _12329_ (.A1(_03192_),
    .A2(_03269_),
    .ZN(_03276_));
 AND2_X2 _12330_ (.A1(_03259_),
    .A2(_03260_),
    .ZN(_03277_));
 OAI33_X1 _12331_ (.A1(_03272_),
    .A2(_03274_),
    .A3(_03275_),
    .B1(_03227_),
    .B2(_03276_),
    .B3(_03277_),
    .ZN(_03278_));
 NOR2_X1 _12332_ (.A1(_03250_),
    .A2(_03149_),
    .ZN(_03279_));
 OAI21_X1 _12333_ (.A(_03279_),
    .B1(_03019_),
    .B2(_03036_),
    .ZN(_03280_));
 XNOR2_X2 _12334_ (.A(_03117_),
    .B(_03280_),
    .ZN(_03281_));
 OR3_X1 _12335_ (.A1(net41),
    .A2(_03141_),
    .A3(_03149_),
    .ZN(_03282_));
 NAND2_X1 _12336_ (.A1(_03151_),
    .A2(_03282_),
    .ZN(_03283_));
 NOR2_X1 _12337_ (.A1(_03281_),
    .A2(_03283_),
    .ZN(_03284_));
 NAND3_X2 _12338_ (.A1(_03271_),
    .A2(_03278_),
    .A3(_03284_),
    .ZN(_03285_));
 INV_X1 _12339_ (.A(_09131_),
    .ZN(_03286_));
 INV_X1 _12340_ (.A(_09137_),
    .ZN(_03287_));
 INV_X1 _12341_ (.A(_09143_),
    .ZN(_03288_));
 OAI21_X2 _12342_ (.A(_09144_),
    .B1(_09147_),
    .B2(_09146_),
    .ZN(_03289_));
 NAND2_X2 _12343_ (.A1(_03289_),
    .A2(_03288_),
    .ZN(_03290_));
 AND2_X4 _12344_ (.A1(_09141_),
    .A2(_03290_),
    .ZN(_03291_));
 OAI21_X4 _12345_ (.A(_09138_),
    .B1(_03291_),
    .B2(_09140_),
    .ZN(_03292_));
 NAND2_X4 _12346_ (.A1(_03287_),
    .A2(_03292_),
    .ZN(_03293_));
 AOI21_X4 _12347_ (.A(_09134_),
    .B1(_03293_),
    .B2(_09135_),
    .ZN(_03294_));
 INV_X1 _12348_ (.A(_09132_),
    .ZN(_03295_));
 OAI21_X4 _12349_ (.A(_03286_),
    .B1(_03295_),
    .B2(_03294_),
    .ZN(_03296_));
 AND2_X4 _12350_ (.A1(_09129_),
    .A2(_03296_),
    .ZN(_03297_));
 NOR2_X1 _12351_ (.A1(_09128_),
    .A2(_03297_),
    .ZN(_03298_));
 NOR2_X1 _12352_ (.A1(_03102_),
    .A2(_03298_),
    .ZN(_03299_));
 OR2_X4 _12353_ (.A1(_03297_),
    .A2(_09128_),
    .ZN(_03300_));
 NAND2_X2 _12354_ (.A1(_03300_),
    .A2(_03102_),
    .ZN(_03301_));
 NAND2_X1 _12355_ (.A1(_02797_),
    .A2(_03301_),
    .ZN(_03302_));
 XNOR2_X2 _12356_ (.A(_09109_),
    .B(_03030_),
    .ZN(_03303_));
 MUX2_X1 _12357_ (.A(_03299_),
    .B(_03302_),
    .S(_03303_),
    .Z(_03304_));
 NOR2_X1 _12358_ (.A1(_08985_),
    .A2(_02374_),
    .ZN(_09004_));
 OR3_X1 _12359_ (.A1(_09006_),
    .A2(_02310_),
    .A3(_09008_),
    .ZN(_03305_));
 AND2_X1 _12360_ (.A1(_02390_),
    .A2(_03305_),
    .ZN(_03306_));
 MUX2_X1 _12361_ (.A(_09004_),
    .B(_03306_),
    .S(_02585_),
    .Z(_09027_));
 XOR2_X1 _12362_ (.A(_09029_),
    .B(_02361_),
    .Z(_03307_));
 MUX2_X1 _12363_ (.A(_09027_),
    .B(_03307_),
    .S(_02698_),
    .Z(_09045_));
 OR3_X1 _12364_ (.A1(_09047_),
    .A2(_09049_),
    .A3(_02555_),
    .ZN(_03308_));
 AND2_X1 _12365_ (.A1(_02556_),
    .A2(_03308_),
    .ZN(_03309_));
 MUX2_X1 _12366_ (.A(_09045_),
    .B(_03309_),
    .S(net18),
    .Z(_09066_));
 NOR2_X1 _12367_ (.A1(_09068_),
    .A2(_02662_),
    .ZN(_03310_));
 NOR3_X1 _12368_ (.A1(_02879_),
    .A2(_02881_),
    .A3(_03310_),
    .ZN(_03311_));
 MUX2_X1 _12369_ (.A(_09066_),
    .B(_03311_),
    .S(_02889_),
    .Z(_09086_));
 XNOR2_X1 _12370_ (.A(_03073_),
    .B(_03061_),
    .ZN(_03312_));
 BUF_X8 _12371_ (.A(_03112_),
    .Z(_03313_));
 MUX2_X2 _12372_ (.A(_09086_),
    .B(_03312_),
    .S(net39),
    .Z(_09107_));
 MUX2_X1 _12373_ (.A(_03299_),
    .B(_03302_),
    .S(_09107_),
    .Z(_03314_));
 NOR2_X4 _12374_ (.A1(_03152_),
    .A2(_03202_),
    .ZN(_03315_));
 MUX2_X2 _12375_ (.A(_03304_),
    .B(_03314_),
    .S(_03315_),
    .Z(_03316_));
 OR3_X4 _12376_ (.A1(_03255_),
    .A2(_03316_),
    .A3(_03285_),
    .ZN(_03317_));
 OAI21_X1 _12377_ (.A(_03174_),
    .B1(_03192_),
    .B2(_03269_),
    .ZN(_03318_));
 OR2_X2 _12378_ (.A1(_03227_),
    .A2(_03318_),
    .ZN(_03319_));
 AND2_X1 _12379_ (.A1(_03175_),
    .A2(_03179_),
    .ZN(_03320_));
 INV_X1 _12380_ (.A(_03320_),
    .ZN(_03321_));
 NOR2_X1 _12381_ (.A1(_03036_),
    .A2(_03183_),
    .ZN(_03322_));
 INV_X1 _12382_ (.A(_02956_),
    .ZN(_03323_));
 OAI21_X1 _12383_ (.A(_03212_),
    .B1(_03322_),
    .B2(_03323_),
    .ZN(_03324_));
 AOI21_X1 _12384_ (.A(_03321_),
    .B1(_03324_),
    .B2(net39),
    .ZN(_03325_));
 NOR2_X1 _12385_ (.A1(_03323_),
    .A2(_03181_),
    .ZN(_03326_));
 NOR2_X1 _12386_ (.A1(_03100_),
    .A2(_03149_),
    .ZN(_03327_));
 AOI21_X2 _12387_ (.A(_03325_),
    .B1(_03326_),
    .B2(_03327_),
    .ZN(_03328_));
 AND4_X1 _12388_ (.A1(_03174_),
    .A2(_03202_),
    .A3(_03211_),
    .A4(_03243_),
    .ZN(_03329_));
 AOI221_X2 _12389_ (.A(_03320_),
    .B1(_03184_),
    .B2(_03187_),
    .C1(_03181_),
    .C2(_02956_),
    .ZN(_03330_));
 OAI21_X2 _12390_ (.A(_03330_),
    .B1(_03318_),
    .B2(_03227_),
    .ZN(_03331_));
 OAI22_X4 _12391_ (.A1(_03319_),
    .A2(_03328_),
    .B1(_03329_),
    .B2(_03331_),
    .ZN(_03332_));
 NAND3_X1 _12392_ (.A1(_03202_),
    .A2(_03111_),
    .A3(_03211_),
    .ZN(_03333_));
 XNOR2_X2 _12393_ (.A(_03174_),
    .B(_03333_),
    .ZN(_03334_));
 AOI21_X1 _12394_ (.A(_03197_),
    .B1(_03198_),
    .B2(net39),
    .ZN(_03335_));
 AND3_X1 _12395_ (.A1(net39),
    .A2(_03197_),
    .A3(_03198_),
    .ZN(_03336_));
 NOR3_X1 _12396_ (.A1(_03222_),
    .A2(_03133_),
    .A3(_03226_),
    .ZN(_03337_));
 OR2_X1 _12397_ (.A1(_03222_),
    .A2(_03200_),
    .ZN(_03338_));
 NOR4_X1 _12398_ (.A1(_03121_),
    .A2(_03164_),
    .A3(_03192_),
    .A4(_03269_),
    .ZN(_03339_));
 OR2_X1 _12399_ (.A1(_03133_),
    .A2(_03226_),
    .ZN(_03340_));
 OAI33_X1 _12400_ (.A1(_03335_),
    .A2(_03336_),
    .A3(_03337_),
    .B1(_03338_),
    .B2(_03339_),
    .B3(_03340_),
    .ZN(_03341_));
 NAND2_X1 _12401_ (.A1(_03151_),
    .A2(_03020_),
    .ZN(_03342_));
 AOI21_X2 _12402_ (.A(_03342_),
    .B1(_03056_),
    .B2(_03242_),
    .ZN(_03343_));
 AOI21_X2 _12403_ (.A(_03146_),
    .B1(_03134_),
    .B2(_03343_),
    .ZN(_03344_));
 AND3_X1 _12404_ (.A1(_03146_),
    .A2(_03134_),
    .A3(_03343_),
    .ZN(_03345_));
 NOR2_X4 _12405_ (.A1(_03121_),
    .A2(_03222_),
    .ZN(_03346_));
 NOR4_X4 _12406_ (.A1(_03164_),
    .A2(_03192_),
    .A3(_03200_),
    .A4(_03269_),
    .ZN(_03347_));
 NAND2_X4 _12407_ (.A1(_03346_),
    .A2(_03347_),
    .ZN(_03348_));
 AOI211_X2 _12408_ (.A(_03341_),
    .B(_03344_),
    .C1(_03345_),
    .C2(_03348_),
    .ZN(_03349_));
 NAND4_X4 _12409_ (.A1(_03215_),
    .A2(_03332_),
    .A3(_03334_),
    .A4(_03349_),
    .ZN(_03350_));
 OR3_X4 _12410_ (.A1(_03317_),
    .A2(_03248_),
    .A3(_03350_),
    .ZN(_03351_));
 OR3_X4 clone30 (.A1(_03317_),
    .A2(_03248_),
    .A3(_03350_),
    .ZN(net30));
 BUF_X8 _12412_ (.A(_03351_),
    .Z(_03353_));
 BUF_X8 _12413_ (.A(_03353_),
    .Z(_03354_));
 XNOR2_X1 _12414_ (.A(_03295_),
    .B(_03294_),
    .ZN(_03355_));
 NAND2_X1 _12415_ (.A1(_03354_),
    .A2(_03355_),
    .ZN(_03356_));
 NOR2_X1 _12416_ (.A1(_09026_),
    .A2(_02710_),
    .ZN(_09051_));
 OR3_X1 _12417_ (.A1(_09056_),
    .A2(_09053_),
    .A3(_09055_),
    .ZN(_03357_));
 AND2_X1 _12418_ (.A1(_02553_),
    .A2(_03357_),
    .ZN(_03358_));
 MUX2_X1 _12419_ (.A(_09051_),
    .B(_03358_),
    .S(_02642_),
    .Z(_09072_));
 XOR2_X1 _12420_ (.A(_09074_),
    .B(_02659_),
    .Z(_03359_));
 MUX2_X1 _12421_ (.A(_09072_),
    .B(_03359_),
    .S(_02889_),
    .Z(_09092_));
 INV_X1 _12422_ (.A(_09099_),
    .ZN(_03360_));
 OAI21_X1 _12423_ (.A(_02905_),
    .B1(_09102_),
    .B2(_02912_),
    .ZN(_03361_));
 AOI21_X1 _12424_ (.A(_02907_),
    .B1(_03360_),
    .B2(_03361_),
    .ZN(_03362_));
 NOR2_X1 _12425_ (.A1(_09096_),
    .A2(_03362_),
    .ZN(_03363_));
 XNOR2_X1 _12426_ (.A(_02909_),
    .B(_03363_),
    .ZN(_03364_));
 MUX2_X1 _12427_ (.A(_09092_),
    .B(_03364_),
    .S(_03313_),
    .Z(_09113_));
 XNOR2_X1 _12428_ (.A(_09115_),
    .B(_03027_),
    .ZN(_03365_));
 MUX2_X1 _12429_ (.A(_09113_),
    .B(_03365_),
    .S(_03348_),
    .Z(_09130_));
 OAI21_X1 _12430_ (.A(_03356_),
    .B1(_03354_),
    .B2(_09130_),
    .ZN(_03366_));
 INV_X1 _12431_ (.A(_09154_),
    .ZN(_03367_));
 INV_X1 _12432_ (.A(_09160_),
    .ZN(_03368_));
 OAI21_X2 _12433_ (.A(_09161_),
    .B1(_09163_),
    .B2(_09164_),
    .ZN(_03369_));
 NOR3_X4 _12434_ (.A1(_09163_),
    .A2(_09160_),
    .A3(_09166_),
    .ZN(_03370_));
 OAI21_X2 _12435_ (.A(_09167_),
    .B1(_09148_),
    .B2(_09149_),
    .ZN(_03371_));
 AOI22_X2 _12436_ (.A1(_03368_),
    .A2(_03369_),
    .B1(_03370_),
    .B2(_03371_),
    .ZN(_03372_));
 NAND2_X2 _12437_ (.A1(_03372_),
    .A2(_09158_),
    .ZN(_03373_));
 INV_X4 _12438_ (.A(_03373_),
    .ZN(_03374_));
 OAI21_X4 _12439_ (.A(_09155_),
    .B1(_03374_),
    .B2(_09157_),
    .ZN(_03375_));
 NAND2_X4 _12440_ (.A1(_03367_),
    .A2(_03375_),
    .ZN(_03376_));
 XNOR2_X1 _12441_ (.A(_09152_),
    .B(_03376_),
    .ZN(_03377_));
 INV_X1 _12442_ (.A(_03301_),
    .ZN(_03378_));
 AND3_X1 _12443_ (.A1(_03346_),
    .A2(_03347_),
    .A3(_09107_),
    .ZN(_03379_));
 INV_X1 _12444_ (.A(_03303_),
    .ZN(_03380_));
 AOI21_X4 _12445_ (.A(_03380_),
    .B1(_03347_),
    .B2(_03346_),
    .ZN(_03381_));
 OAI22_X2 _12446_ (.A1(_02573_),
    .A2(_03378_),
    .B1(_03379_),
    .B2(_03381_),
    .ZN(_03382_));
 NAND3_X2 _12447_ (.A1(_03346_),
    .A2(_03347_),
    .A3(_09107_),
    .ZN(_03383_));
 OAI21_X2 _12448_ (.A(_03303_),
    .B1(net16),
    .B2(_03152_),
    .ZN(_03384_));
 NAND3_X1 _12449_ (.A1(_03299_),
    .A2(_03383_),
    .A3(_03384_),
    .ZN(_03385_));
 NAND3_X2 _12450_ (.A1(_03278_),
    .A2(_03382_),
    .A3(_03385_),
    .ZN(_03386_));
 AND2_X2 _12451_ (.A1(_03255_),
    .A2(_03386_),
    .ZN(_03387_));
 AND4_X1 _12452_ (.A1(_03160_),
    .A2(_03163_),
    .A3(_03269_),
    .A4(_03252_),
    .ZN(_03388_));
 OAI21_X1 _12453_ (.A(_03122_),
    .B1(_03019_),
    .B2(_03036_),
    .ZN(_03389_));
 XNOR2_X1 _12454_ (.A(_03057_),
    .B(_03389_),
    .ZN(_03390_));
 AND2_X1 _12455_ (.A1(_03390_),
    .A2(_03252_),
    .ZN(_03391_));
 NAND2_X1 _12456_ (.A1(_03259_),
    .A2(_03260_),
    .ZN(_03392_));
 NAND2_X1 _12457_ (.A1(_03238_),
    .A2(_03241_),
    .ZN(_03393_));
 OAI22_X2 _12458_ (.A1(_02797_),
    .A2(_03392_),
    .B1(_03273_),
    .B2(_03393_),
    .ZN(_03394_));
 OR2_X1 _12459_ (.A1(_03032_),
    .A2(_03252_),
    .ZN(_03395_));
 NOR2_X1 _12460_ (.A1(_03083_),
    .A2(_09104_),
    .ZN(_03396_));
 NAND2_X1 _12461_ (.A1(_02797_),
    .A2(_03083_),
    .ZN(_03397_));
 NOR2_X1 _12462_ (.A1(_03096_),
    .A2(_03397_),
    .ZN(_03398_));
 OAI21_X1 _12463_ (.A(_03100_),
    .B1(_03396_),
    .B2(_03398_),
    .ZN(_03399_));
 NOR2_X1 _12464_ (.A1(_03083_),
    .A2(_03105_),
    .ZN(_03400_));
 NOR2_X1 _12465_ (.A1(_03081_),
    .A2(_03397_),
    .ZN(_03401_));
 OAI21_X1 _12466_ (.A(net39),
    .B1(_03400_),
    .B2(_03401_),
    .ZN(_03402_));
 AOI221_X2 _12467_ (.A(_03395_),
    .B1(_03399_),
    .B2(_03402_),
    .C1(_03056_),
    .C2(_03242_),
    .ZN(_03403_));
 AOI221_X2 _12468_ (.A(_03388_),
    .B1(_03391_),
    .B2(_03394_),
    .C1(_03390_),
    .C2(_03403_),
    .ZN(_03404_));
 INV_X1 _12469_ (.A(_03304_),
    .ZN(_03405_));
 OAI21_X1 _12470_ (.A(_03405_),
    .B1(net16),
    .B2(_03152_),
    .ZN(_03406_));
 OAI33_X1 _12471_ (.A1(_03277_),
    .A2(_03348_),
    .A3(_03314_),
    .B1(_03404_),
    .B2(_03274_),
    .B3(_03406_),
    .ZN(_03407_));
 BUF_X4 _12472_ (.A(_03407_),
    .Z(_03408_));
 OR2_X1 _12473_ (.A1(_03255_),
    .A2(_03285_),
    .ZN(_03409_));
 OR3_X1 _12474_ (.A1(_03409_),
    .A2(_03248_),
    .A3(_03350_),
    .ZN(_03410_));
 BUF_X4 _12475_ (.A(_03410_),
    .Z(_03411_));
 AOI21_X4 _12476_ (.A(_03387_),
    .B1(_03408_),
    .B2(_03411_),
    .ZN(_03412_));
 AOI21_X4 _12477_ (.A(_09151_),
    .B1(_03376_),
    .B2(_09152_),
    .ZN(_03413_));
 NOR2_X1 _12478_ (.A1(_03102_),
    .A2(_03413_),
    .ZN(_03414_));
 OAI21_X4 _12479_ (.A(_02797_),
    .B1(_03413_),
    .B2(_08819_),
    .ZN(_03415_));
 XNOR2_X1 _12480_ (.A(_02310_),
    .B(_02309_),
    .ZN(_03416_));
 MUX2_X1 _12481_ (.A(_09007_),
    .B(_03416_),
    .S(_02585_),
    .Z(_09030_));
 OR3_X1 _12482_ (.A1(_09026_),
    .A2(_09032_),
    .A3(_09025_),
    .ZN(_03417_));
 AND2_X1 _12483_ (.A1(_02360_),
    .A2(_03417_),
    .ZN(_03418_));
 MUX2_X1 _12484_ (.A(_09030_),
    .B(_03418_),
    .S(_02698_),
    .Z(_09048_));
 XOR2_X1 _12485_ (.A(_09050_),
    .B(_02554_),
    .Z(_03419_));
 MUX2_X1 _12486_ (.A(_09048_),
    .B(_03419_),
    .S(_02642_),
    .Z(_09069_));
 INV_X1 _12487_ (.A(_09073_),
    .ZN(_03420_));
 OAI21_X1 _12488_ (.A(_03420_),
    .B1(_02875_),
    .B2(_02819_),
    .ZN(_03421_));
 XOR2_X1 _12489_ (.A(_02655_),
    .B(_03421_),
    .Z(_03422_));
 MUX2_X1 _12490_ (.A(_09069_),
    .B(_03422_),
    .S(_02889_),
    .Z(_09089_));
 NOR2_X1 _12491_ (.A1(_02911_),
    .A2(_02918_),
    .ZN(_03423_));
 XNOR2_X1 _12492_ (.A(_02896_),
    .B(_03423_),
    .ZN(_03424_));
 MUX2_X1 _12493_ (.A(_09089_),
    .B(_03424_),
    .S(_03313_),
    .Z(_09110_));
 NOR3_X1 _12494_ (.A1(_03100_),
    .A2(_03047_),
    .A3(_03049_),
    .ZN(_03425_));
 AOI21_X1 _12495_ (.A(_03425_),
    .B1(_03100_),
    .B2(_03079_),
    .ZN(_03426_));
 OAI21_X1 _12496_ (.A(_03029_),
    .B1(_03040_),
    .B2(_03426_),
    .ZN(_03427_));
 XNOR2_X1 _12497_ (.A(_09112_),
    .B(_03427_),
    .ZN(_03428_));
 MUX2_X1 _12498_ (.A(_09110_),
    .B(_03428_),
    .S(_03348_),
    .Z(_03429_));
 CLKBUF_X3 _12499_ (.A(_03429_),
    .Z(_09127_));
 MUX2_X1 _12500_ (.A(_03414_),
    .B(_03415_),
    .S(_09127_),
    .Z(_03430_));
 XOR2_X2 _12501_ (.A(_09129_),
    .B(_03296_),
    .Z(_03431_));
 MUX2_X1 _12502_ (.A(_03414_),
    .B(_03415_),
    .S(_03431_),
    .Z(_03432_));
 OAI21_X1 _12503_ (.A(_03300_),
    .B1(_03379_),
    .B2(_03381_),
    .ZN(_03433_));
 NAND3_X1 _12504_ (.A1(_03298_),
    .A2(_03383_),
    .A3(_03384_),
    .ZN(_03434_));
 XNOR2_X1 _12505_ (.A(_03102_),
    .B(_03056_),
    .ZN(_03435_));
 OAI21_X2 _12506_ (.A(_03435_),
    .B1(net16),
    .B2(_03152_),
    .ZN(_03436_));
 XNOR2_X2 _12507_ (.A(_03277_),
    .B(_03436_),
    .ZN(_03437_));
 MUX2_X1 _12508_ (.A(_03433_),
    .B(_03434_),
    .S(_03437_),
    .Z(_03438_));
 XNOR2_X1 _12509_ (.A(_02797_),
    .B(_03277_),
    .ZN(_03439_));
 XNOR2_X1 _12510_ (.A(_03436_),
    .B(_03439_),
    .ZN(_03440_));
 AOI21_X1 _12511_ (.A(_03300_),
    .B1(_03383_),
    .B2(_03384_),
    .ZN(_03441_));
 NOR3_X1 _12512_ (.A1(_03298_),
    .A2(_03379_),
    .A3(_03381_),
    .ZN(_03442_));
 XNOR2_X1 _12513_ (.A(_03392_),
    .B(_03436_),
    .ZN(_03443_));
 AOI22_X1 _12514_ (.A1(_03440_),
    .A2(_03441_),
    .B1(_03442_),
    .B2(_03443_),
    .ZN(_03444_));
 MUX2_X1 _12515_ (.A(_03438_),
    .B(_03444_),
    .S(_08819_),
    .Z(_03445_));
 OAI22_X4 _12516_ (.A1(_03351_),
    .A2(_03430_),
    .B1(_03432_),
    .B2(_03445_),
    .ZN(_03446_));
 AND2_X1 _12517_ (.A1(_03348_),
    .A2(_03345_),
    .ZN(_03447_));
 OR2_X1 _12518_ (.A1(_03447_),
    .A2(_03344_),
    .ZN(_03448_));
 AND3_X1 _12519_ (.A1(_03151_),
    .A2(_03281_),
    .A3(_03282_),
    .ZN(_03449_));
 OAI21_X1 _12520_ (.A(_03252_),
    .B1(_03225_),
    .B2(_03224_),
    .ZN(_03450_));
 OR2_X1 _12521_ (.A1(_03133_),
    .A2(_03450_),
    .ZN(_03451_));
 MUX2_X1 _12522_ (.A(_03449_),
    .B(_03284_),
    .S(_03451_),
    .Z(_03452_));
 OR2_X2 _12523_ (.A1(_03315_),
    .A2(_03452_),
    .ZN(_03453_));
 AND2_X1 _12524_ (.A1(_03205_),
    .A2(_03453_),
    .ZN(_03454_));
 NAND2_X1 _12525_ (.A1(_03164_),
    .A2(_03269_),
    .ZN(_03455_));
 OR2_X1 _12526_ (.A1(_03164_),
    .A2(_03269_),
    .ZN(_03456_));
 OAI21_X1 _12527_ (.A(_03455_),
    .B1(_03315_),
    .B2(_03456_),
    .ZN(_03457_));
 INV_X1 _12528_ (.A(_03457_),
    .ZN(_03458_));
 NOR3_X1 _12529_ (.A1(_03277_),
    .A2(_03348_),
    .A3(_03314_),
    .ZN(_03459_));
 NOR2_X1 _12530_ (.A1(_03274_),
    .A2(_03406_),
    .ZN(_03460_));
 OR2_X2 _12531_ (.A1(_03459_),
    .A2(_03460_),
    .ZN(_03461_));
 OAI211_X2 _12532_ (.A(_03454_),
    .B(_03386_),
    .C1(_03458_),
    .C2(_03461_),
    .ZN(_03462_));
 NOR2_X1 _12533_ (.A1(_03102_),
    .A2(_03300_),
    .ZN(_03463_));
 NOR2_X2 _12534_ (.A1(_03379_),
    .A2(_03381_),
    .ZN(_03464_));
 NOR3_X1 _12535_ (.A1(_02573_),
    .A2(_03443_),
    .A3(_03464_),
    .ZN(_03465_));
 NOR2_X1 _12536_ (.A1(_02797_),
    .A2(_03437_),
    .ZN(_03466_));
 OAI21_X2 _12537_ (.A(_03463_),
    .B1(_03465_),
    .B2(_03466_),
    .ZN(_03467_));
 NAND2_X1 _12538_ (.A1(_03383_),
    .A2(_03384_),
    .ZN(_03468_));
 NOR2_X2 _12539_ (.A1(_03437_),
    .A2(_03468_),
    .ZN(_03469_));
 NAND2_X1 _12540_ (.A1(_03300_),
    .A2(_03437_),
    .ZN(_03470_));
 NOR2_X1 _12541_ (.A1(_08819_),
    .A2(_03441_),
    .ZN(_03471_));
 AOI21_X2 _12542_ (.A(_03469_),
    .B1(_03470_),
    .B2(_03471_),
    .ZN(_03472_));
 AOI221_X2 _12543_ (.A(_03448_),
    .B1(_03351_),
    .B2(_03462_),
    .C1(_03467_),
    .C2(_03472_),
    .ZN(_03473_));
 AND3_X4 _12544_ (.A1(_03446_),
    .A2(_03412_),
    .A3(_03473_),
    .ZN(_03474_));
 BUF_X2 clone11 (.A(_01407_),
    .Z(net11));
 XOR2_X2 _12546_ (.A(_03207_),
    .B(_03214_),
    .Z(_03476_));
 MUX2_X1 _12547_ (.A(_03171_),
    .B(_03172_),
    .S(_03173_),
    .Z(_03477_));
 NOR2_X1 _12548_ (.A1(_03323_),
    .A2(_03322_),
    .ZN(_03478_));
 OR2_X1 _12549_ (.A1(_03227_),
    .A2(_03339_),
    .ZN(_03479_));
 NOR4_X2 _12550_ (.A1(_03477_),
    .A2(_03320_),
    .A3(_03478_),
    .A4(_03479_),
    .ZN(_03480_));
 XNOR2_X2 _12551_ (.A(_03476_),
    .B(_03480_),
    .ZN(_03481_));
 AND3_X1 _12552_ (.A1(_03332_),
    .A2(_03334_),
    .A3(_03349_),
    .ZN(_03482_));
 AND3_X2 _12553_ (.A1(_03205_),
    .A2(_03453_),
    .A3(_03408_),
    .ZN(_03483_));
 AOI21_X4 _12554_ (.A(_03481_),
    .B1(_03482_),
    .B2(_03483_),
    .ZN(_03484_));
 AND3_X1 _12555_ (.A1(_03218_),
    .A2(_03229_),
    .A3(_03247_),
    .ZN(_03485_));
 NAND2_X1 _12556_ (.A1(_03271_),
    .A2(_03485_),
    .ZN(_03486_));
 NOR2_X4 _12557_ (.A1(_03484_),
    .A2(_03486_),
    .ZN(_03487_));
 OAI21_X1 _12558_ (.A(_03200_),
    .B1(_03340_),
    .B2(_03222_),
    .ZN(_03488_));
 AND2_X1 _12559_ (.A1(_03479_),
    .A2(_03488_),
    .ZN(_03489_));
 NOR2_X2 _12560_ (.A1(_03447_),
    .A2(_03344_),
    .ZN(_03490_));
 AOI21_X2 _12561_ (.A(_03489_),
    .B1(_03490_),
    .B2(_03483_),
    .ZN(_03491_));
 AND2_X1 _12562_ (.A1(_03349_),
    .A2(_03483_),
    .ZN(_03492_));
 AOI21_X4 _12563_ (.A(_03491_),
    .B1(_03492_),
    .B2(_03351_),
    .ZN(_03493_));
 INV_X1 _12564_ (.A(_03332_),
    .ZN(_03494_));
 NAND2_X1 _12565_ (.A1(_03334_),
    .A2(_03349_),
    .ZN(_03495_));
 NAND3_X4 _12566_ (.A1(_03205_),
    .A2(_03453_),
    .A3(_03408_),
    .ZN(_03496_));
 NOR2_X1 _12567_ (.A1(_03495_),
    .A2(_03496_),
    .ZN(_03497_));
 NAND2_X1 _12568_ (.A1(_03349_),
    .A2(_03483_),
    .ZN(_03498_));
 INV_X1 _12569_ (.A(_03334_),
    .ZN(_03499_));
 AOI221_X4 _12570_ (.A(_03494_),
    .B1(_03351_),
    .B2(_03497_),
    .C1(_03498_),
    .C2(_03499_),
    .ZN(_03500_));
 AND3_X4 _12571_ (.A1(_03487_),
    .A2(_03493_),
    .A3(_03500_),
    .ZN(_03501_));
 NAND2_X4 _12572_ (.A1(_03474_),
    .A2(_03501_),
    .ZN(_03502_));
 MUX2_X2 _12573_ (.A(_03366_),
    .B(_03377_),
    .S(_03502_),
    .Z(_03503_));
 INV_X1 _12574_ (.A(_03503_),
    .ZN(_09186_));
 NAND3_X4 _12575_ (.A1(_03446_),
    .A2(_03412_),
    .A3(_03473_),
    .ZN(_03504_));
 NAND3_X4 _12576_ (.A1(_03487_),
    .A2(_03493_),
    .A3(_03500_),
    .ZN(_03505_));
 NOR2_X4 _12577_ (.A1(_03504_),
    .A2(_03505_),
    .ZN(_03506_));
 NAND2_X1 _12578_ (.A1(_02751_),
    .A2(net29),
    .ZN(_03507_));
 INV_X1 _12579_ (.A(_08981_),
    .ZN(_03508_));
 NAND2_X1 _12580_ (.A1(_02309_),
    .A2(net35),
    .ZN(_03509_));
 NAND3_X2 _12581_ (.A1(_03507_),
    .A2(_03508_),
    .A3(_03509_),
    .ZN(_09054_));
 NOR2_X4 _12582_ (.A1(_09054_),
    .A2(_02642_),
    .ZN(_03510_));
 AOI21_X4 _12583_ (.A(_03510_),
    .B1(_02642_),
    .B2(_09056_),
    .ZN(_09075_));
 NAND2_X1 _12584_ (.A1(_03045_),
    .A2(_02876_),
    .ZN(_03511_));
 AOI21_X1 _12585_ (.A(_09078_),
    .B1(_03511_),
    .B2(_09079_),
    .ZN(_03512_));
 XNOR2_X1 _12586_ (.A(_09077_),
    .B(_03512_),
    .ZN(_03513_));
 MUX2_X1 _12587_ (.A(_09075_),
    .B(_03513_),
    .S(_02889_),
    .Z(_09095_));
 AOI21_X1 _12588_ (.A(_09102_),
    .B1(_03033_),
    .B2(_02912_),
    .ZN(_03514_));
 INV_X1 _12589_ (.A(_02905_),
    .ZN(_03515_));
 OAI21_X1 _12590_ (.A(_03360_),
    .B1(_03514_),
    .B2(_03515_),
    .ZN(_03516_));
 XNOR2_X1 _12591_ (.A(_02907_),
    .B(_03516_),
    .ZN(_03517_));
 MUX2_X1 _12592_ (.A(_09095_),
    .B(_03517_),
    .S(_03313_),
    .Z(_09116_));
 AOI21_X1 _12593_ (.A(_09125_),
    .B1(_03426_),
    .B2(_09126_),
    .ZN(_03518_));
 NAND2_X1 _12594_ (.A1(_09121_),
    .A2(_09124_),
    .ZN(_03519_));
 OAI21_X1 _12595_ (.A(_03023_),
    .B1(_03518_),
    .B2(_03519_),
    .ZN(_03520_));
 XOR2_X1 _12596_ (.A(_09118_),
    .B(_03520_),
    .Z(_03521_));
 MUX2_X1 _12597_ (.A(_09116_),
    .B(_03521_),
    .S(_03348_),
    .Z(_09133_));
 XOR2_X1 _12598_ (.A(_09135_),
    .B(_03293_),
    .Z(_03522_));
 MUX2_X1 _12599_ (.A(_09133_),
    .B(_03522_),
    .S(_03354_),
    .Z(_09153_));
 NAND2_X1 _12600_ (.A1(_03506_),
    .A2(_09153_),
    .ZN(_03523_));
 BUF_X8 _12601_ (.A(_03502_),
    .Z(_03524_));
 NOR2_X1 _12602_ (.A1(_09148_),
    .A2(_03003_),
    .ZN(_03525_));
 NAND2_X1 _12603_ (.A1(_03048_),
    .A2(_03525_),
    .ZN(_03526_));
 NOR2_X1 _12604_ (.A1(_02103_),
    .A2(_02796_),
    .ZN(_03527_));
 XNOR2_X1 _12605_ (.A(_02757_),
    .B(_03527_),
    .ZN(_03528_));
 NAND3_X2 _12606_ (.A1(_03054_),
    .A2(_03052_),
    .A3(_03528_),
    .ZN(_03529_));
 NAND2_X1 _12607_ (.A1(_02799_),
    .A2(_02353_),
    .ZN(_03530_));
 XNOR2_X1 _12608_ (.A(_02112_),
    .B(_02796_),
    .ZN(_03531_));
 XNOR2_X1 _12609_ (.A(_03530_),
    .B(_03531_),
    .ZN(_03532_));
 AOI21_X2 _12610_ (.A(_02745_),
    .B1(_03532_),
    .B2(_01710_),
    .ZN(_03533_));
 OAI21_X4 _12611_ (.A(_03533_),
    .B1(_03019_),
    .B2(_03036_),
    .ZN(_03534_));
 AOI211_X2 _12612_ (.A(_01929_),
    .B(_03526_),
    .C1(_03529_),
    .C2(_03534_),
    .ZN(_03535_));
 AOI21_X2 _12613_ (.A(_03373_),
    .B1(_03535_),
    .B2(_03370_),
    .ZN(_03536_));
 NOR2_X1 _12614_ (.A1(_09157_),
    .A2(_03536_),
    .ZN(_03537_));
 XNOR2_X1 _12615_ (.A(_09155_),
    .B(_03537_),
    .ZN(_03538_));
 NAND2_X1 _12616_ (.A1(_03524_),
    .A2(_03538_),
    .ZN(_03539_));
 AND2_X1 _12617_ (.A1(_03523_),
    .A2(_03539_),
    .ZN(_03540_));
 CLKBUF_X2 _12618_ (.A(_09191_),
    .Z(_03541_));
 INV_X1 _12619_ (.A(_03541_),
    .ZN(_03542_));
 AOI21_X2 _12620_ (.A(_09169_),
    .B1(_09172_),
    .B2(_09170_),
    .ZN(_03543_));
 INV_X1 _12621_ (.A(_09178_),
    .ZN(_03544_));
 BUF_X1 _12622_ (.A(_09182_),
    .Z(_03545_));
 AOI21_X1 _12623_ (.A(_09181_),
    .B1(_09184_),
    .B2(_03545_),
    .ZN(_03546_));
 INV_X1 _12624_ (.A(_09179_),
    .ZN(_03547_));
 OAI21_X1 _12625_ (.A(_03544_),
    .B1(_03546_),
    .B2(_03547_),
    .ZN(_03548_));
 BUF_X2 _12626_ (.A(_09176_),
    .Z(_03549_));
 AOI21_X1 _12627_ (.A(_09175_),
    .B1(_03548_),
    .B2(_03549_),
    .ZN(_03550_));
 AND2_X1 _12628_ (.A1(_09170_),
    .A2(_09173_),
    .ZN(_03551_));
 NAND2_X4 _12629_ (.A1(_03534_),
    .A2(_03529_),
    .ZN(_03552_));
 XNOR2_X2 _12630_ (.A(net38),
    .B(_03552_),
    .ZN(_03553_));
 OAI21_X2 _12631_ (.A(_03551_),
    .B1(_03553_),
    .B2(_01929_),
    .ZN(_03554_));
 NAND4_X1 _12632_ (.A1(_03542_),
    .A2(_03543_),
    .A3(_03550_),
    .A4(_03554_),
    .ZN(_03555_));
 NAND2_X1 _12633_ (.A1(_03545_),
    .A2(_09185_),
    .ZN(_03556_));
 NAND2_X1 _12634_ (.A1(_03549_),
    .A2(_09179_),
    .ZN(_03557_));
 OR4_X1 _12635_ (.A1(_03542_),
    .A2(_03556_),
    .A3(_03557_),
    .A4(_03554_),
    .ZN(_03558_));
 NOR4_X1 _12636_ (.A1(_03542_),
    .A2(_03543_),
    .A3(_03556_),
    .A4(_03557_),
    .ZN(_03559_));
 NOR2_X2 _12637_ (.A1(_03556_),
    .A2(_03557_),
    .ZN(_03560_));
 NOR2_X1 _12638_ (.A1(_03541_),
    .A2(_03560_),
    .ZN(_03561_));
 MUX2_X1 _12639_ (.A(_03541_),
    .B(_03561_),
    .S(_03550_),
    .Z(_03562_));
 NOR2_X1 _12640_ (.A1(_03559_),
    .A2(_03562_),
    .ZN(_03563_));
 NAND3_X1 _12641_ (.A1(_03555_),
    .A2(_03558_),
    .A3(_03563_),
    .ZN(_03564_));
 BUF_X2 _12642_ (.A(_09188_),
    .Z(_03565_));
 INV_X1 _12643_ (.A(_09190_),
    .ZN(_03566_));
 INV_X1 _12644_ (.A(_09184_),
    .ZN(_03567_));
 INV_X1 _12645_ (.A(_09185_),
    .ZN(_03568_));
 OAI21_X2 _12646_ (.A(_03567_),
    .B1(_03568_),
    .B2(_03543_),
    .ZN(_03569_));
 AOI21_X2 _12647_ (.A(_09181_),
    .B1(_03569_),
    .B2(_03545_),
    .ZN(_03570_));
 OAI21_X2 _12648_ (.A(_03544_),
    .B1(_03570_),
    .B2(_03547_),
    .ZN(_03571_));
 AOI21_X2 _12649_ (.A(_09175_),
    .B1(_03549_),
    .B2(_03571_),
    .ZN(_03572_));
 OAI21_X2 _12650_ (.A(_03566_),
    .B1(_03572_),
    .B2(_03542_),
    .ZN(_03573_));
 AOI21_X2 _12651_ (.A(_09187_),
    .B1(_03565_),
    .B2(_03573_),
    .ZN(_03574_));
 NAND4_X2 _12652_ (.A1(_03565_),
    .A2(_03541_),
    .A3(_03560_),
    .A4(_03551_),
    .ZN(_03575_));
 AOI21_X1 _12653_ (.A(_01929_),
    .B1(_03534_),
    .B2(_03529_),
    .ZN(_03576_));
 OAI21_X1 _12654_ (.A(_03574_),
    .B1(_03575_),
    .B2(_03576_),
    .ZN(_03577_));
 AND2_X1 _12655_ (.A1(_03468_),
    .A2(_09127_),
    .ZN(_03578_));
 INV_X1 _12656_ (.A(_03431_),
    .ZN(_03579_));
 NOR2_X1 _12657_ (.A1(_03378_),
    .A2(_03463_),
    .ZN(_03580_));
 XNOR2_X1 _12658_ (.A(_03464_),
    .B(_03580_),
    .ZN(_03581_));
 NOR2_X1 _12659_ (.A1(_03579_),
    .A2(_03581_),
    .ZN(_03582_));
 MUX2_X1 _12660_ (.A(_03578_),
    .B(_03582_),
    .S(net32),
    .Z(_03583_));
 AND2_X1 _12661_ (.A1(_09152_),
    .A2(_09155_),
    .ZN(_03584_));
 NAND2_X1 _12662_ (.A1(_09155_),
    .A2(_09157_),
    .ZN(_03585_));
 NAND2_X1 _12663_ (.A1(_03367_),
    .A2(_03585_),
    .ZN(_03586_));
 AOI221_X2 _12664_ (.A(_09151_),
    .B1(_03536_),
    .B2(_03584_),
    .C1(_03586_),
    .C2(_09152_),
    .ZN(_03587_));
 XNOR2_X2 _12665_ (.A(_03102_),
    .B(_03587_),
    .ZN(_03588_));
 NOR2_X1 _12666_ (.A1(_03415_),
    .A2(_03588_),
    .ZN(_03589_));
 INV_X1 _12667_ (.A(_03415_),
    .ZN(_03590_));
 NOR2_X1 _12668_ (.A1(_03590_),
    .A2(_03588_),
    .ZN(_03591_));
 NAND2_X1 _12669_ (.A1(_03464_),
    .A2(_03580_),
    .ZN(_03592_));
 OR2_X1 _12670_ (.A1(_03464_),
    .A2(_03580_),
    .ZN(_03593_));
 NOR3_X4 _12671_ (.A1(_03248_),
    .A2(_03317_),
    .A3(_03350_),
    .ZN(_03594_));
 OR2_X1 _12672_ (.A1(_03350_),
    .A2(_03468_),
    .ZN(_03595_));
 OR2_X2 _12673_ (.A1(_03248_),
    .A2(_03317_),
    .ZN(_03596_));
 OAI221_X2 _12674_ (.A(_03592_),
    .B1(_03593_),
    .B2(_03594_),
    .C1(_03595_),
    .C2(_03596_),
    .ZN(_03597_));
 BUF_X4 _12675_ (.A(_03597_),
    .Z(_03598_));
 AOI22_X2 _12676_ (.A1(_03583_),
    .A2(_03589_),
    .B1(_03591_),
    .B2(_03598_),
    .ZN(_03599_));
 OR2_X1 _12677_ (.A1(_03102_),
    .A2(_03413_),
    .ZN(_03600_));
 NAND2_X1 _12678_ (.A1(_03600_),
    .A2(_03588_),
    .ZN(_03601_));
 NOR2_X1 _12679_ (.A1(_09127_),
    .A2(_03601_),
    .ZN(_03602_));
 NOR2_X1 _12680_ (.A1(_03431_),
    .A2(_03601_),
    .ZN(_03603_));
 MUX2_X1 _12681_ (.A(_03602_),
    .B(_03603_),
    .S(_03353_),
    .Z(_03604_));
 INV_X1 _12682_ (.A(_09127_),
    .ZN(_03605_));
 MUX2_X2 _12683_ (.A(_03605_),
    .B(_03579_),
    .S(_03353_),
    .Z(_03606_));
 AOI21_X2 _12684_ (.A(_03604_),
    .B1(_03598_),
    .B2(_03606_),
    .ZN(_03607_));
 AND2_X1 _12685_ (.A1(_03599_),
    .A2(_03607_),
    .ZN(_03608_));
 OR2_X1 _12686_ (.A1(_03102_),
    .A2(_03587_),
    .ZN(_03609_));
 NOR2_X1 _12687_ (.A1(_09127_),
    .A2(_03609_),
    .ZN(_03610_));
 NOR2_X1 _12688_ (.A1(_03431_),
    .A2(_03609_),
    .ZN(_03611_));
 MUX2_X2 _12689_ (.A(_03610_),
    .B(_03611_),
    .S(net30),
    .Z(_03612_));
 MUX2_X1 _12690_ (.A(_03604_),
    .B(_03612_),
    .S(_03597_),
    .Z(_03613_));
 NOR2_X1 _12691_ (.A1(_03606_),
    .A2(_03588_),
    .ZN(_03614_));
 XNOR2_X1 _12692_ (.A(_03415_),
    .B(_03598_),
    .ZN(_03615_));
 AOI21_X1 _12693_ (.A(_03613_),
    .B1(_03614_),
    .B2(_03615_),
    .ZN(_03616_));
 OR2_X1 _12694_ (.A1(_02745_),
    .A2(_03575_),
    .ZN(_03617_));
 NAND2_X1 _12695_ (.A1(_03574_),
    .A2(_03617_),
    .ZN(_03618_));
 OAI21_X1 _12696_ (.A(_03408_),
    .B1(_03248_),
    .B2(_03409_),
    .ZN(_03619_));
 AOI22_X2 _12697_ (.A1(_03255_),
    .A2(_03386_),
    .B1(_03408_),
    .B2(_03350_),
    .ZN(_03620_));
 NAND2_X2 _12698_ (.A1(_03619_),
    .A2(_03620_),
    .ZN(_03621_));
 AND2_X1 _12699_ (.A1(_03316_),
    .A2(_03437_),
    .ZN(_03622_));
 INV_X1 _12700_ (.A(_03622_),
    .ZN(_03623_));
 NOR2_X1 _12701_ (.A1(_03459_),
    .A2(_03460_),
    .ZN(_03624_));
 OAI21_X2 _12702_ (.A(_03623_),
    .B1(_03594_),
    .B2(_03624_),
    .ZN(_03625_));
 OR2_X1 _12703_ (.A1(_03621_),
    .A2(_03625_),
    .ZN(_03626_));
 NAND2_X1 _12704_ (.A1(_03412_),
    .A2(_03625_),
    .ZN(_03627_));
 OR2_X1 _12705_ (.A1(_09127_),
    .A2(_03609_),
    .ZN(_03628_));
 OR2_X1 _12706_ (.A1(_03431_),
    .A2(_03609_),
    .ZN(_03629_));
 MUX2_X2 _12707_ (.A(_03628_),
    .B(_03629_),
    .S(net30),
    .Z(_03630_));
 OAI21_X2 _12708_ (.A(_02797_),
    .B1(_08819_),
    .B2(_03587_),
    .ZN(_03631_));
 NAND2_X1 _12709_ (.A1(_09127_),
    .A2(_03631_),
    .ZN(_03632_));
 NAND2_X1 _12710_ (.A1(_03431_),
    .A2(_03631_),
    .ZN(_03633_));
 MUX2_X1 _12711_ (.A(_03632_),
    .B(_03633_),
    .S(net30),
    .Z(_03634_));
 AND3_X2 _12712_ (.A1(_03630_),
    .A2(_03634_),
    .A3(_03597_),
    .ZN(_03635_));
 MUX2_X2 _12713_ (.A(_03626_),
    .B(_03627_),
    .S(_03635_),
    .Z(_03636_));
 OAI33_X1 _12714_ (.A1(_03577_),
    .A2(_03502_),
    .A3(_03608_),
    .B1(_03618_),
    .B2(_03616_),
    .B3(_03636_),
    .ZN(_03637_));
 INV_X1 _12715_ (.A(_03625_),
    .ZN(_03638_));
 NAND2_X2 _12716_ (.A1(_03467_),
    .A2(_03472_),
    .ZN(_03639_));
 NAND2_X2 _12717_ (.A1(net403),
    .A2(_03639_),
    .ZN(_03640_));
 AOI21_X4 _12718_ (.A(_03638_),
    .B1(_03635_),
    .B2(_03640_),
    .ZN(_03641_));
 OAI21_X2 _12719_ (.A(_03386_),
    .B1(_03458_),
    .B2(_03461_),
    .ZN(_03642_));
 NAND2_X1 _12720_ (.A1(_03354_),
    .A2(_03642_),
    .ZN(_03643_));
 NAND2_X1 _12721_ (.A1(_03281_),
    .A2(_03451_),
    .ZN(_03644_));
 OAI21_X2 _12722_ (.A(_03644_),
    .B1(_03340_),
    .B2(_03315_),
    .ZN(_03645_));
 NAND2_X1 _12723_ (.A1(_03645_),
    .A2(_03408_),
    .ZN(_03646_));
 OR2_X1 _12724_ (.A1(_03645_),
    .A2(_03408_),
    .ZN(_03647_));
 NAND3_X4 _12725_ (.A1(_03411_),
    .A2(_03646_),
    .A3(_03647_),
    .ZN(_03648_));
 NAND2_X1 _12726_ (.A1(_03643_),
    .A2(_03648_),
    .ZN(_03649_));
 NOR2_X2 _12727_ (.A1(_03641_),
    .A2(_03649_),
    .ZN(_03650_));
 INV_X1 _12728_ (.A(_03645_),
    .ZN(_03651_));
 AOI21_X2 _12729_ (.A(_03205_),
    .B1(_03651_),
    .B2(_03408_),
    .ZN(_03652_));
 XOR2_X1 _12730_ (.A(_03020_),
    .B(_03204_),
    .Z(_03653_));
 NOR2_X1 _12731_ (.A1(_03653_),
    .A2(_03645_),
    .ZN(_03654_));
 AND2_X1 _12732_ (.A1(_03408_),
    .A2(_03654_),
    .ZN(_03655_));
 AOI21_X4 _12733_ (.A(_03652_),
    .B1(_03655_),
    .B2(_03411_),
    .ZN(_03656_));
 INV_X1 _12734_ (.A(_03656_),
    .ZN(_03657_));
 OR3_X1 _12735_ (.A1(_03645_),
    .A2(_03622_),
    .A3(_03457_),
    .ZN(_03658_));
 AOI211_X2 _12736_ (.A(_03658_),
    .B(_03387_),
    .C1(_03411_),
    .C2(_03461_),
    .ZN(_03659_));
 NAND4_X2 _12737_ (.A1(_03630_),
    .A2(_03634_),
    .A3(_03598_),
    .A4(_03659_),
    .ZN(_03660_));
 AOI211_X2 _12738_ (.A(_03657_),
    .B(_03660_),
    .C1(_03474_),
    .C2(_03501_),
    .ZN(_03661_));
 AND4_X1 _12739_ (.A1(_03630_),
    .A2(_03634_),
    .A3(_03598_),
    .A4(_03659_),
    .ZN(_03662_));
 NOR2_X2 _12740_ (.A1(_03656_),
    .A2(_03662_),
    .ZN(_03663_));
 NAND2_X2 _12741_ (.A1(_03353_),
    .A2(_03462_),
    .ZN(_03664_));
 NAND4_X4 _12742_ (.A1(_03412_),
    .A2(_03664_),
    .A3(_03446_),
    .A4(_03639_),
    .ZN(_03665_));
 NAND2_X2 _12743_ (.A1(_03448_),
    .A2(_03483_),
    .ZN(_03666_));
 NAND2_X2 _12744_ (.A1(_03490_),
    .A2(_03496_),
    .ZN(_03667_));
 NAND3_X4 _12745_ (.A1(net30),
    .A2(_03666_),
    .A3(_03667_),
    .ZN(_03668_));
 AND4_X2 _12746_ (.A1(_03487_),
    .A2(_03493_),
    .A3(_03500_),
    .A4(_03668_),
    .ZN(_03669_));
 AOI221_X2 _12747_ (.A(_03387_),
    .B1(_03408_),
    .B2(_03411_),
    .C1(_03642_),
    .C2(_03353_),
    .ZN(_03670_));
 AND4_X1 _12748_ (.A1(_03446_),
    .A2(_03639_),
    .A3(_03654_),
    .A4(_03670_),
    .ZN(_03671_));
 NOR2_X1 _12749_ (.A1(_03594_),
    .A2(_03496_),
    .ZN(_03672_));
 NAND3_X1 _12750_ (.A1(_03135_),
    .A2(_03020_),
    .A3(_03272_),
    .ZN(_03673_));
 NOR3_X1 _12751_ (.A1(_03315_),
    .A2(_03283_),
    .A3(_03673_),
    .ZN(_03674_));
 AOI21_X1 _12752_ (.A(_03674_),
    .B1(_03673_),
    .B2(_03283_),
    .ZN(_03675_));
 AOI21_X1 _12753_ (.A(_03675_),
    .B1(_03655_),
    .B2(_03411_),
    .ZN(_03676_));
 NOR2_X1 _12754_ (.A1(_03672_),
    .A2(_03676_),
    .ZN(_03677_));
 OAI22_X4 _12755_ (.A1(_03665_),
    .A2(_03669_),
    .B1(_03671_),
    .B2(_03677_),
    .ZN(_03678_));
 NOR3_X4 _12756_ (.A1(_03661_),
    .A2(_03663_),
    .A3(_03678_),
    .ZN(_03679_));
 NAND3_X4 _12757_ (.A1(_03679_),
    .A2(_03650_),
    .A3(net376),
    .ZN(_03680_));
 XOR2_X2 _12758_ (.A(_03210_),
    .B(_03217_),
    .Z(_03681_));
 AND4_X1 _12759_ (.A1(_03271_),
    .A2(_03218_),
    .A3(_03229_),
    .A4(_03247_),
    .ZN(_03682_));
 NOR3_X4 _12760_ (.A1(_03350_),
    .A2(_03496_),
    .A3(_03682_),
    .ZN(_03683_));
 XNOR2_X2 _12761_ (.A(_03681_),
    .B(_03683_),
    .ZN(_03684_));
 INV_X1 _12762_ (.A(_03684_),
    .ZN(_03685_));
 XNOR2_X1 _12763_ (.A(_03490_),
    .B(_03483_),
    .ZN(_03686_));
 NAND2_X1 _12764_ (.A1(_03489_),
    .A2(_03334_),
    .ZN(_03687_));
 OAI21_X1 _12765_ (.A(net32),
    .B1(_03686_),
    .B2(_03687_),
    .ZN(_03688_));
 NOR2_X1 _12766_ (.A1(_03478_),
    .A2(_03214_),
    .ZN(_03689_));
 AND3_X1 _12767_ (.A1(_03321_),
    .A2(_03208_),
    .A3(_03329_),
    .ZN(_03690_));
 XNOR2_X2 _12768_ (.A(_03689_),
    .B(_03690_),
    .ZN(_03691_));
 OR2_X1 _12769_ (.A1(_03495_),
    .A2(_03496_),
    .ZN(_03692_));
 OAI21_X1 _12770_ (.A(_03691_),
    .B1(_03692_),
    .B2(_03594_),
    .ZN(_03693_));
 NAND3_X1 _12771_ (.A1(_03332_),
    .A2(_03334_),
    .A3(_03349_),
    .ZN(_03694_));
 NOR4_X2 _12772_ (.A1(_03255_),
    .A2(_03285_),
    .A3(_03476_),
    .A4(_03316_),
    .ZN(_03695_));
 AND4_X1 _12773_ (.A1(_03205_),
    .A2(_03218_),
    .A3(_03229_),
    .A4(_03247_),
    .ZN(_03696_));
 AOI211_X2 _12774_ (.A(_03496_),
    .B(_03694_),
    .C1(_03695_),
    .C2(_03696_),
    .ZN(_03697_));
 NAND2_X1 _12775_ (.A1(_03321_),
    .A2(_03208_),
    .ZN(_03698_));
 XNOR2_X2 _12776_ (.A(_03319_),
    .B(_03698_),
    .ZN(_03699_));
 NOR4_X2 _12777_ (.A1(_03484_),
    .A2(_03697_),
    .A3(_03699_),
    .A4(_03683_),
    .ZN(_03700_));
 AND3_X2 _12778_ (.A1(_03688_),
    .A2(_03693_),
    .A3(_03700_),
    .ZN(_03701_));
 INV_X1 _12779_ (.A(_03701_),
    .ZN(_03702_));
 AND2_X2 _12780_ (.A1(_03412_),
    .A2(_03664_),
    .ZN(_03703_));
 AND2_X1 _12781_ (.A1(_09127_),
    .A2(_03631_),
    .ZN(_03704_));
 AND2_X1 _12782_ (.A1(_03431_),
    .A2(_03631_),
    .ZN(_03705_));
 MUX2_X2 _12783_ (.A(_03704_),
    .B(_03705_),
    .S(net30),
    .Z(_03706_));
 NAND2_X1 _12784_ (.A1(_03102_),
    .A2(_03438_),
    .ZN(_03707_));
 NAND2_X1 _12785_ (.A1(_08819_),
    .A2(_03444_),
    .ZN(_03708_));
 AOI22_X4 _12786_ (.A1(_03594_),
    .A2(_03469_),
    .B1(_03707_),
    .B2(_03708_),
    .ZN(_03709_));
 NOR3_X4 _12787_ (.A1(_03612_),
    .A2(_03706_),
    .A3(_03709_),
    .ZN(_03710_));
 OAI211_X4 _12788_ (.A(_03703_),
    .B(_03710_),
    .C1(_03505_),
    .C2(net402),
    .ZN(_03711_));
 OAI21_X4 _12789_ (.A(_03685_),
    .B1(_03702_),
    .B2(_03711_),
    .ZN(_03712_));
 NAND2_X1 _12790_ (.A1(_03412_),
    .A2(_03664_),
    .ZN(_03713_));
 OR3_X2 _12791_ (.A1(_03612_),
    .A2(_03706_),
    .A3(_03709_),
    .ZN(_03714_));
 AOI211_X4 _12792_ (.A(_03713_),
    .B(_03714_),
    .C1(_03501_),
    .C2(_03474_),
    .ZN(_03715_));
 NAND3_X4 _12793_ (.A1(_03684_),
    .A2(_03701_),
    .A3(_03715_),
    .ZN(_03716_));
 NOR2_X1 _12794_ (.A1(_03484_),
    .A2(_03683_),
    .ZN(_03717_));
 OR2_X1 _12795_ (.A1(_03484_),
    .A2(_03486_),
    .ZN(_03718_));
 NAND2_X1 _12796_ (.A1(_03718_),
    .A2(_03717_),
    .ZN(_03719_));
 NAND2_X1 _12797_ (.A1(_03493_),
    .A2(_03500_),
    .ZN(_03720_));
 NOR2_X1 _12798_ (.A1(_03504_),
    .A2(_03720_),
    .ZN(_03721_));
 MUX2_X2 _12799_ (.A(_03717_),
    .B(_03719_),
    .S(_03721_),
    .Z(_03722_));
 NAND3_X4 _12800_ (.A1(_03712_),
    .A2(_03716_),
    .A3(_03722_),
    .ZN(_03723_));
 OR2_X1 _12801_ (.A1(_03350_),
    .A2(_03496_),
    .ZN(_03724_));
 NAND2_X1 _12802_ (.A1(_03681_),
    .A2(_03724_),
    .ZN(_03725_));
 NAND4_X1 _12803_ (.A1(_03688_),
    .A2(_03693_),
    .A3(_03700_),
    .A4(_03725_),
    .ZN(_03726_));
 OAI33_X1 _12804_ (.A1(_03681_),
    .A2(_03682_),
    .A3(_03724_),
    .B1(_03726_),
    .B2(_03665_),
    .B3(_03669_),
    .ZN(_03727_));
 XOR2_X2 _12805_ (.A(_03229_),
    .B(_03727_),
    .Z(_03728_));
 NOR2_X2 _12806_ (.A1(_03350_),
    .A2(_03496_),
    .ZN(_03729_));
 NAND4_X2 _12807_ (.A1(_03218_),
    .A2(_03229_),
    .A3(_03596_),
    .A4(_03729_),
    .ZN(_03730_));
 XOR2_X2 _12808_ (.A(_03247_),
    .B(_03730_),
    .Z(_03731_));
 AND2_X1 _12809_ (.A1(_03229_),
    .A2(_03684_),
    .ZN(_03732_));
 AND2_X1 _12810_ (.A1(_03701_),
    .A2(_03732_),
    .ZN(_03733_));
 AOI21_X4 _12811_ (.A(_03731_),
    .B1(_03733_),
    .B2(_03715_),
    .ZN(_03734_));
 AND4_X2 _12812_ (.A1(_03701_),
    .A2(_03715_),
    .A3(_03731_),
    .A4(_03732_),
    .ZN(_03735_));
 OAI21_X4 _12813_ (.A(_03728_),
    .B1(_03734_),
    .B2(_03735_),
    .ZN(_03736_));
 NAND2_X2 _12814_ (.A1(net32),
    .A2(_03497_),
    .ZN(_03737_));
 NAND2_X1 _12815_ (.A1(_03499_),
    .A2(_03498_),
    .ZN(_03738_));
 AND2_X2 _12816_ (.A1(_03737_),
    .A2(_03738_),
    .ZN(_03739_));
 AND3_X2 _12817_ (.A1(net32),
    .A2(_03666_),
    .A3(_03667_),
    .ZN(_03740_));
 NOR2_X4 _12818_ (.A1(net377),
    .A2(_03740_),
    .ZN(_03741_));
 OAI211_X4 _12819_ (.A(net402),
    .B(_03741_),
    .C1(_03714_),
    .C2(_03713_),
    .ZN(_03742_));
 NAND4_X4 _12820_ (.A1(_03703_),
    .A2(_03493_),
    .A3(_03740_),
    .A4(_03710_),
    .ZN(_03743_));
 NAND3_X4 _12821_ (.A1(_03502_),
    .A2(_03742_),
    .A3(_03743_),
    .ZN(_03744_));
 XNOR2_X2 _12822_ (.A(_03737_),
    .B(_03699_),
    .ZN(_03745_));
 OR3_X1 _12823_ (.A1(_03697_),
    .A2(_03691_),
    .A3(_03745_),
    .ZN(_03746_));
 INV_X2 _12824_ (.A(_03746_),
    .ZN(_03747_));
 NAND3_X4 _12825_ (.A1(_03739_),
    .A2(_03744_),
    .A3(_03747_),
    .ZN(_03748_));
 NOR4_X4 _12826_ (.A1(_03680_),
    .A2(_03723_),
    .A3(_03736_),
    .A4(_03748_),
    .ZN(_03749_));
 OR2_X1 _12827_ (.A1(_03504_),
    .A2(_03720_),
    .ZN(_03750_));
 OAI21_X2 _12828_ (.A(_03724_),
    .B1(_03750_),
    .B2(_03484_),
    .ZN(_03751_));
 AOI21_X4 _12829_ (.A(_03271_),
    .B1(_03485_),
    .B2(_03751_),
    .ZN(_03752_));
 AOI211_X2 _12830_ (.A(_03504_),
    .B(_03505_),
    .C1(_03599_),
    .C2(_03607_),
    .ZN(_03753_));
 OR2_X1 _12831_ (.A1(_09127_),
    .A2(_03601_),
    .ZN(_03754_));
 NAND3_X1 _12832_ (.A1(_03600_),
    .A2(_03579_),
    .A3(_03588_),
    .ZN(_03755_));
 MUX2_X1 _12833_ (.A(_03754_),
    .B(_03755_),
    .S(_03354_),
    .Z(_03756_));
 MUX2_X1 _12834_ (.A(_03756_),
    .B(_03630_),
    .S(_03598_),
    .Z(_03757_));
 OR2_X1 _12835_ (.A1(_03606_),
    .A2(_03588_),
    .ZN(_03758_));
 XNOR2_X1 _12836_ (.A(_03590_),
    .B(_03598_),
    .ZN(_03759_));
 OAI21_X2 _12837_ (.A(_03757_),
    .B1(_03758_),
    .B2(_03759_),
    .ZN(_03760_));
 AND2_X2 _12838_ (.A1(net32),
    .A2(_03642_),
    .ZN(_03761_));
 NOR2_X1 _12839_ (.A1(_03761_),
    .A2(_03625_),
    .ZN(_03762_));
 AND2_X1 _12840_ (.A1(_03643_),
    .A2(_03625_),
    .ZN(_03763_));
 MUX2_X1 _12841_ (.A(_03762_),
    .B(_03763_),
    .S(_03635_),
    .Z(_03764_));
 AOI21_X1 _12842_ (.A(_03753_),
    .B1(_03760_),
    .B2(_03764_),
    .ZN(_03765_));
 OAI211_X2 _12843_ (.A(_03656_),
    .B(_03662_),
    .C1(_03504_),
    .C2(_03505_),
    .ZN(_03766_));
 NAND2_X1 _12844_ (.A1(_03657_),
    .A2(_03660_),
    .ZN(_03767_));
 AND4_X1 _12845_ (.A1(_03412_),
    .A2(_03664_),
    .A3(net403),
    .A4(_03639_),
    .ZN(_03768_));
 NAND4_X2 _12846_ (.A1(_03487_),
    .A2(_03493_),
    .A3(_03500_),
    .A4(_03668_),
    .ZN(_03769_));
 NAND4_X2 _12847_ (.A1(_03446_),
    .A2(_03639_),
    .A3(_03654_),
    .A4(_03670_),
    .ZN(_03770_));
 OR2_X1 _12848_ (.A1(_03672_),
    .A2(_03676_),
    .ZN(_03771_));
 AOI22_X4 _12849_ (.A1(_03768_),
    .A2(_03769_),
    .B1(_03770_),
    .B2(_03771_),
    .ZN(_03772_));
 NOR2_X4 _12850_ (.A1(_03315_),
    .A2(_02103_),
    .ZN(_03773_));
 XNOR2_X1 _12851_ (.A(_03552_),
    .B(_03773_),
    .ZN(_03774_));
 NOR3_X1 _12852_ (.A1(_01170_),
    .A2(_03575_),
    .A3(_03774_),
    .ZN(_03775_));
 NAND4_X1 _12853_ (.A1(_03766_),
    .A2(_03767_),
    .A3(_03772_),
    .A4(_03775_),
    .ZN(_03776_));
 NAND2_X1 _12854_ (.A1(_01150_),
    .A2(_03552_),
    .ZN(_03777_));
 AND2_X1 _12855_ (.A1(_03412_),
    .A2(_03648_),
    .ZN(_03778_));
 AND2_X1 _12856_ (.A1(_03621_),
    .A2(_03648_),
    .ZN(_03779_));
 NOR4_X4 _12857_ (.A1(_03761_),
    .A2(_03612_),
    .A3(_03706_),
    .A4(_03709_),
    .ZN(_03780_));
 MUX2_X1 _12858_ (.A(_03778_),
    .B(_03779_),
    .S(_03780_),
    .Z(_03781_));
 AND4_X1 _12859_ (.A1(_03703_),
    .A2(_03493_),
    .A3(_03740_),
    .A4(_03710_),
    .ZN(_03782_));
 NAND2_X2 _12860_ (.A1(_03489_),
    .A2(_03668_),
    .ZN(_03783_));
 AOI211_X2 _12861_ (.A(_03474_),
    .B(_03783_),
    .C1(_03710_),
    .C2(_03703_),
    .ZN(_03784_));
 OAI211_X2 _12862_ (.A(_03777_),
    .B(_03781_),
    .C1(_03782_),
    .C2(_03784_),
    .ZN(_03785_));
 AOI211_X2 _12863_ (.A(_03765_),
    .B(_03776_),
    .C1(_03502_),
    .C2(_03785_),
    .ZN(_03786_));
 NOR2_X4 _12864_ (.A1(_03752_),
    .A2(_03786_),
    .ZN(_03787_));
 BUF_X8 _12865_ (.A(_03787_),
    .Z(_03788_));
 NAND2_X4 _12866_ (.A1(_03749_),
    .A2(_03788_),
    .ZN(_03789_));
 MUX2_X2 _12867_ (.A(_03540_),
    .B(_03564_),
    .S(_03789_),
    .Z(_03790_));
 INV_X1 _12868_ (.A(_03790_),
    .ZN(_09200_));
 BUF_X8 _12869_ (.A(_03789_),
    .Z(_03791_));
 INV_X1 _12870_ (.A(_09181_),
    .ZN(_03792_));
 NAND2_X1 _12871_ (.A1(_09170_),
    .A2(_09173_),
    .ZN(_03793_));
 NAND2_X1 _12872_ (.A1(_03543_),
    .A2(_03793_),
    .ZN(_03794_));
 AOI21_X1 _12873_ (.A(_09184_),
    .B1(_03794_),
    .B2(_09185_),
    .ZN(_03795_));
 INV_X1 _12874_ (.A(_03545_),
    .ZN(_03796_));
 OAI21_X1 _12875_ (.A(_03792_),
    .B1(_03795_),
    .B2(_03796_),
    .ZN(_03797_));
 AOI21_X2 _12876_ (.A(_09178_),
    .B1(_03797_),
    .B2(_09179_),
    .ZN(_03798_));
 XOR2_X1 _12877_ (.A(_03549_),
    .B(_03798_),
    .Z(_03799_));
 NAND2_X1 _12878_ (.A1(net23),
    .A2(_03799_),
    .ZN(_03800_));
 NOR2_X2 _12879_ (.A1(_09079_),
    .A2(_02796_),
    .ZN(_09098_));
 OR3_X1 _12880_ (.A1(_02912_),
    .A2(_02905_),
    .A3(_09102_),
    .ZN(_03801_));
 AND2_X1 _12881_ (.A1(_03361_),
    .A2(_03801_),
    .ZN(_03802_));
 MUX2_X1 _12882_ (.A(_09098_),
    .B(_03802_),
    .S(_03313_),
    .Z(_09119_));
 INV_X1 _12883_ (.A(_09123_),
    .ZN(_03803_));
 NAND2_X1 _12884_ (.A1(_03803_),
    .A2(_03024_),
    .ZN(_03804_));
 XNOR2_X1 _12885_ (.A(_03025_),
    .B(_03804_),
    .ZN(_03805_));
 MUX2_X1 _12886_ (.A(_09119_),
    .B(_03805_),
    .S(_03348_),
    .Z(_09136_));
 OR3_X1 _12887_ (.A1(_09138_),
    .A2(_09140_),
    .A3(_03291_),
    .ZN(_03806_));
 AND2_X1 _12888_ (.A1(_03292_),
    .A2(_03806_),
    .ZN(_03807_));
 MUX2_X1 _12889_ (.A(_09136_),
    .B(_03807_),
    .S(_03354_),
    .Z(_09156_));
 XOR2_X1 _12890_ (.A(_09158_),
    .B(_03372_),
    .Z(_03808_));
 MUX2_X1 _12891_ (.A(_09156_),
    .B(_03808_),
    .S(_03524_),
    .Z(_09174_));
 OAI21_X1 _12892_ (.A(_03800_),
    .B1(_09174_),
    .B2(net23),
    .ZN(_03809_));
 INV_X1 _12893_ (.A(_03809_),
    .ZN(_09203_));
 INV_X1 _12894_ (.A(_09207_),
    .ZN(_03810_));
 INV_X1 _12895_ (.A(_09213_),
    .ZN(_03811_));
 INV_X1 _12896_ (.A(_09196_),
    .ZN(_03812_));
 OAI21_X2 _12897_ (.A(_09197_),
    .B1(_09198_),
    .B2(_09199_),
    .ZN(_03813_));
 NAND2_X2 _12898_ (.A1(_03813_),
    .A2(_03812_),
    .ZN(_03814_));
 AND2_X4 _12899_ (.A1(_09194_),
    .A2(_03814_),
    .ZN(_03815_));
 OAI21_X4 _12900_ (.A(_09214_),
    .B1(_09193_),
    .B2(_03815_),
    .ZN(_03816_));
 NAND2_X4 _12901_ (.A1(_03816_),
    .A2(_03811_),
    .ZN(_03817_));
 AND2_X4 _12902_ (.A1(_09211_),
    .A2(_03817_),
    .ZN(_03818_));
 OAI21_X4 _12903_ (.A(_09208_),
    .B1(_03818_),
    .B2(_09210_),
    .ZN(_03819_));
 NAND2_X4 _12904_ (.A1(_03810_),
    .A2(_03819_),
    .ZN(_03820_));
 XNOR2_X1 _12905_ (.A(_09205_),
    .B(_03820_),
    .ZN(_03821_));
 INV_X1 _12906_ (.A(_03821_),
    .ZN(_03822_));
 INV_X1 _12907_ (.A(_03739_),
    .ZN(_03823_));
 AOI21_X4 _12908_ (.A(_03823_),
    .B1(_03741_),
    .B2(_03715_),
    .ZN(_03824_));
 NOR3_X4 _12909_ (.A1(_03739_),
    .A2(_03783_),
    .A3(_03711_),
    .ZN(_03825_));
 OAI21_X2 _12910_ (.A(_03747_),
    .B1(_03824_),
    .B2(_03825_),
    .ZN(_03826_));
 AOI21_X2 _12911_ (.A(_03668_),
    .B1(_03710_),
    .B2(_03703_),
    .ZN(_03827_));
 AOI211_X2 _12912_ (.A(_03678_),
    .B(_03827_),
    .C1(_03715_),
    .C2(_03668_),
    .ZN(_03828_));
 NAND3_X1 _12913_ (.A1(_03332_),
    .A2(_03737_),
    .A3(_03738_),
    .ZN(_03829_));
 OAI21_X1 _12914_ (.A(_03493_),
    .B1(_03829_),
    .B2(_03718_),
    .ZN(_03830_));
 MUX2_X2 _12915_ (.A(_03493_),
    .B(_03830_),
    .S(net21),
    .Z(_03831_));
 NAND2_X1 _12916_ (.A1(_03828_),
    .A2(_03831_),
    .ZN(_03832_));
 OR2_X2 _12917_ (.A1(_03826_),
    .A2(_03832_),
    .ZN(_03833_));
 NAND2_X2 _12918_ (.A1(_03712_),
    .A2(_03716_),
    .ZN(_03834_));
 NAND2_X1 _12919_ (.A1(_03598_),
    .A2(_03656_),
    .ZN(_03835_));
 NAND3_X1 _12920_ (.A1(_03630_),
    .A2(_03634_),
    .A3(_03659_),
    .ZN(_03836_));
 MUX2_X2 _12921_ (.A(_03415_),
    .B(_03414_),
    .S(_03606_),
    .Z(_03837_));
 AOI221_X2 _12922_ (.A(_03835_),
    .B1(_03836_),
    .B2(_03837_),
    .C1(_03474_),
    .C2(_03501_),
    .ZN(_03838_));
 AND2_X1 _12923_ (.A1(_03411_),
    .A2(_03655_),
    .ZN(_03839_));
 NOR3_X1 _12924_ (.A1(_03598_),
    .A2(_03652_),
    .A3(_03839_),
    .ZN(_03840_));
 MUX2_X1 _12925_ (.A(_03657_),
    .B(_03840_),
    .S(_03837_),
    .Z(_03841_));
 NOR3_X2 _12926_ (.A1(_03663_),
    .A2(_03838_),
    .A3(_03841_),
    .ZN(_03842_));
 NAND3_X1 _12927_ (.A1(_03549_),
    .A2(_03565_),
    .A3(_03541_),
    .ZN(_03843_));
 NOR2_X1 _12928_ (.A1(_03798_),
    .A2(_03843_),
    .ZN(_03844_));
 INV_X1 _12929_ (.A(_03565_),
    .ZN(_03845_));
 AOI21_X1 _12930_ (.A(_09190_),
    .B1(_09175_),
    .B2(_03541_),
    .ZN(_03846_));
 NOR2_X1 _12931_ (.A1(_03845_),
    .A2(_03846_),
    .ZN(_03847_));
 NOR3_X2 _12932_ (.A1(_09187_),
    .A2(_03844_),
    .A3(_03847_),
    .ZN(_03848_));
 XNOR2_X2 _12933_ (.A(_03606_),
    .B(_03588_),
    .ZN(_03849_));
 AND2_X1 _12934_ (.A1(_03643_),
    .A2(_03648_),
    .ZN(_03850_));
 OAI211_X2 _12935_ (.A(_03849_),
    .B(_03850_),
    .C1(net402),
    .C2(_03505_),
    .ZN(_03851_));
 OAI33_X1 _12936_ (.A1(_03718_),
    .A2(_03750_),
    .A3(_03608_),
    .B1(_03636_),
    .B2(_03641_),
    .B3(_03851_),
    .ZN(_03852_));
 NAND3_X2 _12937_ (.A1(_03842_),
    .A2(_03848_),
    .A3(_03852_),
    .ZN(_03853_));
 NOR3_X1 _12938_ (.A1(_03834_),
    .A2(_03722_),
    .A3(_03853_),
    .ZN(_03854_));
 NOR4_X2 _12939_ (.A1(_03641_),
    .A2(_03649_),
    .A3(_03661_),
    .A4(_03663_),
    .ZN(_03855_));
 AND2_X1 _12940_ (.A1(net376),
    .A2(_03855_),
    .ZN(_03856_));
 AND3_X1 _12941_ (.A1(_03834_),
    .A2(_03722_),
    .A3(_03856_),
    .ZN(_03857_));
 AOI21_X1 _12942_ (.A(_03854_),
    .B1(_03857_),
    .B2(_03853_),
    .ZN(_03858_));
 NAND2_X1 _12943_ (.A1(net376),
    .A2(_03855_),
    .ZN(_03859_));
 NOR2_X1 _12944_ (.A1(_03859_),
    .A2(_03833_),
    .ZN(_03860_));
 OAI221_X2 _12945_ (.A(_03789_),
    .B1(_03833_),
    .B2(_03858_),
    .C1(_03860_),
    .C2(_03723_),
    .ZN(_03861_));
 NOR2_X1 _12946_ (.A1(_03826_),
    .A2(_03832_),
    .ZN(_03862_));
 NOR2_X2 _12947_ (.A1(_03723_),
    .A2(_03853_),
    .ZN(_03863_));
 AOI21_X2 _12948_ (.A(_03728_),
    .B1(_03862_),
    .B2(_03863_),
    .ZN(_03864_));
 AND3_X1 _12949_ (.A1(_03728_),
    .A2(_03862_),
    .A3(_03863_),
    .ZN(_03865_));
 AOI21_X4 _12950_ (.A(_03864_),
    .B1(_03865_),
    .B2(_03789_),
    .ZN(_03866_));
 BUF_X4 _12951_ (.A(_03866_),
    .Z(_03867_));
 INV_X1 _12952_ (.A(_03271_),
    .ZN(_03868_));
 NAND3_X2 _12953_ (.A1(_03218_),
    .A2(_03229_),
    .A3(_03247_),
    .ZN(_03869_));
 AOI21_X2 _12954_ (.A(_03729_),
    .B1(_03717_),
    .B2(_03721_),
    .ZN(_03870_));
 OAI21_X4 _12955_ (.A(_03868_),
    .B1(_03869_),
    .B2(_03870_),
    .ZN(_03871_));
 NOR3_X2 _12956_ (.A1(_03736_),
    .A2(_03826_),
    .A3(_03832_),
    .ZN(_03872_));
 AOI21_X4 _12957_ (.A(_03871_),
    .B1(_03863_),
    .B2(_03872_),
    .ZN(_03873_));
 OR4_X1 _12958_ (.A1(_03680_),
    .A2(_03723_),
    .A3(_03736_),
    .A4(_03748_),
    .ZN(_03874_));
 BUF_X4 _12959_ (.A(_03874_),
    .Z(_03875_));
 OAI211_X4 _12960_ (.A(_03747_),
    .B(_03728_),
    .C1(_03824_),
    .C2(_03825_),
    .ZN(_03876_));
 NAND4_X4 _12961_ (.A1(_03744_),
    .A2(_03712_),
    .A3(_03716_),
    .A4(_03722_),
    .ZN(_03877_));
 NOR3_X4 _12962_ (.A1(_03680_),
    .A2(_03876_),
    .A3(_03877_),
    .ZN(_03878_));
 OR2_X2 _12963_ (.A1(_03734_),
    .A2(_03735_),
    .ZN(_03879_));
 OAI22_X4 _12964_ (.A1(_03875_),
    .A2(_03787_),
    .B1(_03878_),
    .B2(_03879_),
    .ZN(_03880_));
 NOR2_X4 _12965_ (.A1(_03873_),
    .A2(_03880_),
    .ZN(_03881_));
 OR2_X1 _12966_ (.A1(_03737_),
    .A2(_03699_),
    .ZN(_03882_));
 AOI21_X2 _12967_ (.A(_03697_),
    .B1(_03882_),
    .B2(_03691_),
    .ZN(_03883_));
 NOR2_X1 _12968_ (.A1(_03687_),
    .A2(_03686_),
    .ZN(_03884_));
 NOR2_X2 _12969_ (.A1(_03594_),
    .A2(_03884_),
    .ZN(_03885_));
 NOR3_X2 _12970_ (.A1(_03699_),
    .A2(_03885_),
    .A3(_03711_),
    .ZN(_03886_));
 XOR2_X2 _12971_ (.A(_03883_),
    .B(_03886_),
    .Z(_03887_));
 INV_X2 _12972_ (.A(_03577_),
    .ZN(_03888_));
 NAND2_X2 _12973_ (.A1(_03888_),
    .A2(_03753_),
    .ZN(_03889_));
 AND2_X2 _12974_ (.A1(_03574_),
    .A2(_03617_),
    .ZN(_03890_));
 NAND3_X1 _12975_ (.A1(_03760_),
    .A2(_03890_),
    .A3(_03764_),
    .ZN(_03891_));
 NAND2_X1 _12976_ (.A1(_03889_),
    .A2(_03891_),
    .ZN(_03892_));
 OAI21_X1 _12977_ (.A(_03781_),
    .B1(_03782_),
    .B2(_03784_),
    .ZN(_03893_));
 NAND2_X1 _12978_ (.A1(net38),
    .A2(_03893_),
    .ZN(_03894_));
 AND3_X2 _12979_ (.A1(_03679_),
    .A2(_03892_),
    .A3(_03894_),
    .ZN(_03895_));
 NOR2_X2 _12980_ (.A1(_03824_),
    .A2(_03825_),
    .ZN(_03896_));
 NOR3_X4 _12981_ (.A1(_03665_),
    .A2(_03669_),
    .A3(_03885_),
    .ZN(_03897_));
 XOR2_X2 _12982_ (.A(_03745_),
    .B(_03897_),
    .Z(_03898_));
 NOR2_X1 _12983_ (.A1(_03896_),
    .A2(_03898_),
    .ZN(_03899_));
 AOI21_X4 _12984_ (.A(_03887_),
    .B1(_03895_),
    .B2(_03899_),
    .ZN(_03900_));
 NOR3_X4 _12985_ (.A1(_03723_),
    .A2(_03736_),
    .A3(_03748_),
    .ZN(_03901_));
 AOI211_X2 _12986_ (.A(_03859_),
    .B(_03833_),
    .C1(_03901_),
    .C2(_03787_),
    .ZN(_03902_));
 AOI21_X2 _12987_ (.A(_03827_),
    .B1(_03715_),
    .B2(_03668_),
    .ZN(_03903_));
 AND2_X1 _12988_ (.A1(_03678_),
    .A2(_03903_),
    .ZN(_03904_));
 AND3_X2 _12989_ (.A1(_03842_),
    .A2(_03848_),
    .A3(_03852_),
    .ZN(_03905_));
 MUX2_X1 _12990_ (.A(_03772_),
    .B(_03904_),
    .S(_03905_),
    .Z(_03906_));
 MUX2_X1 _12991_ (.A(_03856_),
    .B(_03680_),
    .S(_03903_),
    .Z(_03907_));
 AOI22_X4 _12992_ (.A1(_03749_),
    .A2(_03788_),
    .B1(_03906_),
    .B2(_03907_),
    .ZN(_03908_));
 NOR3_X4 _12993_ (.A1(_03900_),
    .A2(_03902_),
    .A3(_03908_),
    .ZN(_03909_));
 AND4_X4 _12994_ (.A1(_03861_),
    .A2(_03867_),
    .A3(_03881_),
    .A4(_03909_),
    .ZN(_03910_));
 XNOR2_X2 _12995_ (.A(_03745_),
    .B(_03897_),
    .ZN(_03911_));
 NAND2_X1 _12996_ (.A1(_03896_),
    .A2(_03911_),
    .ZN(_03912_));
 AND4_X1 _12997_ (.A1(_03766_),
    .A2(_03767_),
    .A3(_03772_),
    .A4(_03775_),
    .ZN(_03913_));
 AND2_X1 _12998_ (.A1(_03760_),
    .A2(_03764_),
    .ZN(_03914_));
 NAND2_X1 _12999_ (.A1(_03412_),
    .A2(_03648_),
    .ZN(_03915_));
 NAND2_X1 _13000_ (.A1(_03621_),
    .A2(_03648_),
    .ZN(_03916_));
 MUX2_X1 _13001_ (.A(_03915_),
    .B(_03916_),
    .S(_03780_),
    .Z(_03917_));
 AOI221_X2 _13002_ (.A(_03917_),
    .B1(_03743_),
    .B2(_03742_),
    .C1(_01150_),
    .C2(_03552_),
    .ZN(_03918_));
 OAI221_X2 _13003_ (.A(_03913_),
    .B1(_03914_),
    .B2(_03753_),
    .C1(net428),
    .C2(_03918_),
    .ZN(_03919_));
 NAND2_X4 _13004_ (.A1(_03871_),
    .A2(_03919_),
    .ZN(_03920_));
 OAI21_X2 _13005_ (.A(_03895_),
    .B1(_03920_),
    .B2(_03875_),
    .ZN(_03921_));
 MUX2_X1 _13006_ (.A(_03912_),
    .B(_03896_),
    .S(_03921_),
    .Z(_03922_));
 NAND2_X1 _13007_ (.A1(_03828_),
    .A2(_03905_),
    .ZN(_03923_));
 AOI21_X4 _13008_ (.A(_03923_),
    .B1(_03787_),
    .B2(_03749_),
    .ZN(_03924_));
 XNOR2_X2 _13009_ (.A(_03831_),
    .B(_03924_),
    .ZN(_03925_));
 NOR3_X4 _13010_ (.A1(_03898_),
    .A2(_03922_),
    .A3(_03925_),
    .ZN(_03926_));
 OAI21_X1 _13011_ (.A(net38),
    .B1(_03636_),
    .B2(_03761_),
    .ZN(_03927_));
 XNOR2_X2 _13012_ (.A(_03598_),
    .B(_03837_),
    .ZN(_03928_));
 OR2_X2 _13013_ (.A1(_03506_),
    .A2(_03928_),
    .ZN(_03929_));
 OAI21_X1 _13014_ (.A(_03849_),
    .B1(_03505_),
    .B2(net402),
    .ZN(_03930_));
 OAI21_X2 _13015_ (.A(_03930_),
    .B1(_03608_),
    .B2(net20),
    .ZN(_03931_));
 AND2_X1 _13016_ (.A1(_03848_),
    .A2(_03931_),
    .ZN(_03932_));
 NAND3_X1 _13017_ (.A1(_03927_),
    .A2(_03929_),
    .A3(_03932_),
    .ZN(_03933_));
 AOI21_X2 _13018_ (.A(_03933_),
    .B1(_03787_),
    .B2(_03749_),
    .ZN(_03934_));
 NAND2_X1 _13019_ (.A1(net38),
    .A2(_03648_),
    .ZN(_03935_));
 NOR3_X1 _13020_ (.A1(_03621_),
    .A2(_03761_),
    .A3(_03640_),
    .ZN(_03936_));
 MUX2_X2 _13021_ (.A(_03648_),
    .B(_03935_),
    .S(_03936_),
    .Z(_03937_));
 XOR2_X2 _13022_ (.A(_03934_),
    .B(_03937_),
    .Z(_03938_));
 NOR2_X1 _13023_ (.A1(_03412_),
    .A2(_03780_),
    .ZN(_03939_));
 AOI21_X1 _13024_ (.A(_03621_),
    .B1(net21),
    .B2(_03501_),
    .ZN(_03940_));
 AOI21_X2 _13025_ (.A(_03939_),
    .B1(_03940_),
    .B2(_03780_),
    .ZN(_03941_));
 OAI22_X1 _13026_ (.A1(net38),
    .A2(_03608_),
    .B1(_03616_),
    .B2(_03636_),
    .ZN(_03942_));
 NAND3_X1 _13027_ (.A1(_03650_),
    .A2(_03679_),
    .A3(_03942_),
    .ZN(_03943_));
 NAND3_X2 _13028_ (.A1(_03892_),
    .A2(_03941_),
    .A3(_03943_),
    .ZN(_03944_));
 MUX2_X1 _13029_ (.A(_03621_),
    .B(_03940_),
    .S(_03780_),
    .Z(_03945_));
 AOI21_X2 _13030_ (.A(_03945_),
    .B1(_03891_),
    .B2(_03889_),
    .ZN(_03946_));
 OAI21_X2 _13031_ (.A(_03946_),
    .B1(_03877_),
    .B2(_03876_),
    .ZN(_03947_));
 OAI21_X2 _13032_ (.A(_03946_),
    .B1(_03786_),
    .B2(_03752_),
    .ZN(_03948_));
 OR3_X1 _13033_ (.A1(_03734_),
    .A2(_03735_),
    .A3(_03945_),
    .ZN(_03949_));
 MUX2_X1 _13034_ (.A(_03941_),
    .B(_03949_),
    .S(_03892_),
    .Z(_03950_));
 NAND4_X4 _13035_ (.A1(_03944_),
    .A2(_03947_),
    .A3(_03948_),
    .A4(_03950_),
    .ZN(_03951_));
 NAND3_X4 _13036_ (.A1(_03679_),
    .A2(_03901_),
    .A3(_03788_),
    .ZN(_03952_));
 AOI22_X1 _13037_ (.A1(_03637_),
    .A2(_03650_),
    .B1(_03766_),
    .B2(_03767_),
    .ZN(_03953_));
 OR2_X2 _13038_ (.A1(_03856_),
    .A2(_03953_),
    .ZN(_03954_));
 AOI21_X4 _13039_ (.A(_03951_),
    .B1(_03952_),
    .B2(_03954_),
    .ZN(_03955_));
 AOI21_X1 _13040_ (.A(_03714_),
    .B1(_03501_),
    .B2(net21),
    .ZN(_03956_));
 NOR2_X2 _13041_ (.A1(_03641_),
    .A2(_03956_),
    .ZN(_03957_));
 NOR2_X1 _13042_ (.A1(_03761_),
    .A2(net428),
    .ZN(_03958_));
 MUX2_X2 _13043_ (.A(_03958_),
    .B(_03761_),
    .S(_03640_),
    .Z(_03959_));
 AOI22_X4 _13044_ (.A1(_03888_),
    .A2(_03753_),
    .B1(_03760_),
    .B2(_03890_),
    .ZN(_03960_));
 NOR3_X1 _13045_ (.A1(_03957_),
    .A2(_03959_),
    .A3(_03960_),
    .ZN(_03961_));
 OR2_X1 _13046_ (.A1(net428),
    .A2(_03764_),
    .ZN(_03962_));
 AND2_X1 _13047_ (.A1(_03962_),
    .A2(_03960_),
    .ZN(_03963_));
 AOI211_X2 _13048_ (.A(_03961_),
    .B(_03963_),
    .C1(_03749_),
    .C2(_03788_),
    .ZN(_03964_));
 AOI21_X4 _13049_ (.A(_09204_),
    .B1(_03820_),
    .B2(_09205_),
    .ZN(_03965_));
 INV_X4 _13050_ (.A(_03965_),
    .ZN(_03966_));
 AOI21_X4 _13051_ (.A(_09201_),
    .B1(_03966_),
    .B2(_09202_),
    .ZN(_03967_));
 AOI221_X2 _13052_ (.A(_09175_),
    .B1(_03560_),
    .B2(_03794_),
    .C1(_03548_),
    .C2(_03549_),
    .ZN(_03968_));
 OAI21_X2 _13053_ (.A(_03566_),
    .B1(_03968_),
    .B2(_03542_),
    .ZN(_03969_));
 XNOR2_X2 _13054_ (.A(_03565_),
    .B(_03969_),
    .ZN(_03970_));
 NAND2_X1 _13055_ (.A1(_03967_),
    .A2(_03970_),
    .ZN(_03971_));
 MUX2_X1 _13056_ (.A(_03888_),
    .B(_03890_),
    .S(net20),
    .Z(_03972_));
 XNOR2_X2 _13057_ (.A(_03931_),
    .B(_03972_),
    .ZN(_03973_));
 NOR2_X2 _13058_ (.A1(_03971_),
    .A2(_03973_),
    .ZN(_03974_));
 AND4_X4 _13059_ (.A1(_03967_),
    .A2(_03849_),
    .A3(_03928_),
    .A4(net20),
    .ZN(_03975_));
 INV_X1 _13060_ (.A(_09201_),
    .ZN(_03976_));
 INV_X1 _13061_ (.A(_09202_),
    .ZN(_03977_));
 OAI21_X4 _13062_ (.A(_03976_),
    .B1(_03977_),
    .B2(_03965_),
    .ZN(_03978_));
 NOR3_X2 _13063_ (.A1(net20),
    .A2(_03608_),
    .A3(_03978_),
    .ZN(_03979_));
 XNOR2_X2 _13064_ (.A(_03845_),
    .B(_03969_),
    .ZN(_03980_));
 NOR2_X1 _13065_ (.A1(_03890_),
    .A2(_03980_),
    .ZN(_03981_));
 NOR2_X1 _13066_ (.A1(_03888_),
    .A2(_03980_),
    .ZN(_03982_));
 MUX2_X1 _13067_ (.A(_03981_),
    .B(_03982_),
    .S(_03506_),
    .Z(_03983_));
 OAI222_X2 _13068_ (.A1(_03734_),
    .A2(_03735_),
    .B1(_03975_),
    .B2(_03979_),
    .C1(_03983_),
    .C2(_03503_),
    .ZN(_03984_));
 NOR4_X4 _13069_ (.A1(_03877_),
    .A2(_03876_),
    .A3(_03984_),
    .A4(_03680_),
    .ZN(_03985_));
 AOI22_X4 _13070_ (.A1(_03929_),
    .A2(_03974_),
    .B1(_03985_),
    .B2(_03787_),
    .ZN(_03986_));
 NOR2_X4 _13071_ (.A1(_03964_),
    .A2(_03986_),
    .ZN(_03987_));
 AND3_X4 _13072_ (.A1(_03938_),
    .A2(_03955_),
    .A3(_03987_),
    .ZN(_03988_));
 BUF_X8 _13073_ (.A(_03988_),
    .Z(_03989_));
 NAND3_X4 _13074_ (.A1(_03989_),
    .A2(_03926_),
    .A3(_03910_),
    .ZN(_03990_));
 BUF_X8 _13075_ (.A(_03990_),
    .Z(_03991_));
 MUX2_X2 _13076_ (.A(_09203_),
    .B(_03822_),
    .S(net14),
    .Z(_09227_));
 XNOR2_X2 _13077_ (.A(_03048_),
    .B(_02816_),
    .ZN(_09101_));
 XNOR2_X1 _13078_ (.A(_02912_),
    .B(_03079_),
    .ZN(_03992_));
 MUX2_X1 _13079_ (.A(_09101_),
    .B(_03992_),
    .S(_03313_),
    .Z(_09122_));
 XNOR2_X1 _13080_ (.A(_09124_),
    .B(_03518_),
    .ZN(_03993_));
 MUX2_X1 _13081_ (.A(_09122_),
    .B(_03993_),
    .S(_03348_),
    .Z(_09139_));
 XOR2_X1 _13082_ (.A(_09141_),
    .B(_03290_),
    .Z(_03994_));
 MUX2_X1 _13083_ (.A(_09139_),
    .B(_03994_),
    .S(_03354_),
    .Z(_09159_));
 NOR2_X1 _13084_ (.A1(_09149_),
    .A2(_09148_),
    .ZN(_03995_));
 NOR2_X1 _13085_ (.A1(_03995_),
    .A2(_03535_),
    .ZN(_03996_));
 AOI21_X1 _13086_ (.A(_09166_),
    .B1(_03996_),
    .B2(_09167_),
    .ZN(_03997_));
 INV_X1 _13087_ (.A(_03997_),
    .ZN(_03998_));
 AOI21_X1 _13088_ (.A(_09163_),
    .B1(_03998_),
    .B2(_09164_),
    .ZN(_03999_));
 XNOR2_X1 _13089_ (.A(_09161_),
    .B(_03999_),
    .ZN(_04000_));
 MUX2_X1 _13090_ (.A(_09159_),
    .B(_04000_),
    .S(_03524_),
    .Z(_09177_));
 OAI21_X1 _13091_ (.A(_03570_),
    .B1(_03556_),
    .B2(_03554_),
    .ZN(_04001_));
 XNOR2_X1 _13092_ (.A(_03547_),
    .B(_04001_),
    .ZN(_04002_));
 MUX2_X1 _13093_ (.A(_09177_),
    .B(_04002_),
    .S(_03791_),
    .Z(_09206_));
 OR3_X1 _13094_ (.A1(_09208_),
    .A2(_09210_),
    .A3(_03818_),
    .ZN(_04003_));
 AND2_X1 _13095_ (.A1(_03819_),
    .A2(_04003_),
    .ZN(_04004_));
 MUX2_X1 _13096_ (.A(_09206_),
    .B(_04004_),
    .S(_03991_),
    .Z(_09230_));
 BUF_X2 _13097_ (.A(_09232_),
    .Z(_04005_));
 INV_X1 _13098_ (.A(_09237_),
    .ZN(_04006_));
 INV_X1 _13099_ (.A(_09219_),
    .ZN(_04007_));
 BUF_X1 _13100_ (.A(_09226_),
    .Z(_04008_));
 AOI21_X1 _13101_ (.A(_09225_),
    .B1(_02103_),
    .B2(_04008_),
    .ZN(_04009_));
 INV_X1 _13102_ (.A(_04009_),
    .ZN(_04010_));
 AOI21_X2 _13103_ (.A(_09222_),
    .B1(_04010_),
    .B2(_09223_),
    .ZN(_04011_));
 INV_X1 _13104_ (.A(_09220_),
    .ZN(_04012_));
 OAI21_X2 _13105_ (.A(_04007_),
    .B1(_04011_),
    .B2(_04012_),
    .ZN(_04013_));
 BUF_X1 _13106_ (.A(_09217_),
    .Z(_04014_));
 AOI21_X2 _13107_ (.A(_09216_),
    .B1(_04013_),
    .B2(_04014_),
    .ZN(_04015_));
 INV_X1 _13108_ (.A(_09238_),
    .ZN(_04016_));
 OAI21_X2 _13109_ (.A(_04006_),
    .B1(_04015_),
    .B2(_04016_),
    .ZN(_04017_));
 BUF_X1 _13110_ (.A(_09235_),
    .Z(_04018_));
 AOI21_X2 _13111_ (.A(_09234_),
    .B1(_04018_),
    .B2(_04017_),
    .ZN(_04019_));
 XNOR2_X1 _13112_ (.A(_04005_),
    .B(_04019_),
    .ZN(_04020_));
 INV_X1 _13113_ (.A(_03896_),
    .ZN(_04021_));
 NOR2_X1 _13114_ (.A1(_04021_),
    .A2(_03898_),
    .ZN(_04022_));
 MUX2_X2 _13115_ (.A(_04022_),
    .B(_04021_),
    .S(_03921_),
    .Z(_04023_));
 XOR2_X2 _13116_ (.A(_03831_),
    .B(_03924_),
    .Z(_04024_));
 NAND3_X4 _13117_ (.A1(_03911_),
    .A2(_04023_),
    .A3(_04024_),
    .ZN(_04025_));
 NAND4_X4 _13118_ (.A1(_03861_),
    .A2(_03866_),
    .A3(_03881_),
    .A4(_03909_),
    .ZN(_04026_));
 OAI21_X4 _13119_ (.A(_03989_),
    .B1(_04025_),
    .B2(_04026_),
    .ZN(_04027_));
 NAND3_X4 _13120_ (.A1(_03938_),
    .A2(_03955_),
    .A3(_03987_),
    .ZN(_04028_));
 NAND3_X1 _13121_ (.A1(_03772_),
    .A2(net5),
    .A3(_03905_),
    .ZN(_04029_));
 OAI21_X2 _13122_ (.A(_04029_),
    .B1(_03905_),
    .B2(_03772_),
    .ZN(_04030_));
 NAND2_X2 _13123_ (.A1(_04028_),
    .A2(_04030_),
    .ZN(_04031_));
 XNOR2_X2 _13124_ (.A(_03934_),
    .B(_03937_),
    .ZN(_04032_));
 OR3_X2 _13125_ (.A1(_03951_),
    .A2(_03964_),
    .A3(_03986_),
    .ZN(_04033_));
 NOR2_X4 _13126_ (.A1(_04032_),
    .A2(_04033_),
    .ZN(_04034_));
 NAND2_X4 _13127_ (.A1(_03952_),
    .A2(_03954_),
    .ZN(_04035_));
 OAI211_X4 _13128_ (.A(_04027_),
    .B(_04031_),
    .C1(_04034_),
    .C2(_04035_),
    .ZN(_04036_));
 NAND4_X2 _13129_ (.A1(_03911_),
    .A2(_04023_),
    .A3(_04024_),
    .A4(_04035_),
    .ZN(_04037_));
 OAI21_X4 _13130_ (.A(_04034_),
    .B1(_04037_),
    .B2(_04026_),
    .ZN(_04038_));
 AND2_X1 _13131_ (.A1(_03944_),
    .A2(_03947_),
    .ZN(_04039_));
 AND2_X1 _13132_ (.A1(_03948_),
    .A2(_03950_),
    .ZN(_04040_));
 OR3_X1 _13133_ (.A1(_03957_),
    .A2(_03959_),
    .A3(_03960_),
    .ZN(_04041_));
 NAND2_X1 _13134_ (.A1(_03962_),
    .A2(_03960_),
    .ZN(_04042_));
 OAI211_X2 _13135_ (.A(_04041_),
    .B(_04042_),
    .C1(_03875_),
    .C2(_03920_),
    .ZN(_04043_));
 NOR2_X1 _13136_ (.A1(net428),
    .A2(_03928_),
    .ZN(_04044_));
 NAND2_X1 _13137_ (.A1(_03503_),
    .A2(_03967_),
    .ZN(_04045_));
 OAI33_X1 _13138_ (.A1(_04044_),
    .A2(_03971_),
    .A3(_03973_),
    .B1(_04045_),
    .B2(_03875_),
    .B3(_03920_),
    .ZN(_04046_));
 AOI22_X4 _13139_ (.A1(_04039_),
    .A2(_04040_),
    .B1(_04043_),
    .B2(net375),
    .ZN(_04047_));
 OR2_X1 _13140_ (.A1(_03641_),
    .A2(_03956_),
    .ZN(_04048_));
 OR2_X2 _13141_ (.A1(_04048_),
    .A2(_03960_),
    .ZN(_04049_));
 AOI21_X2 _13142_ (.A(_04049_),
    .B1(_03919_),
    .B2(_03871_),
    .ZN(_04050_));
 AND4_X1 _13143_ (.A1(_03744_),
    .A2(_03712_),
    .A3(_03716_),
    .A4(_03722_),
    .ZN(_04051_));
 XNOR2_X1 _13144_ (.A(_03229_),
    .B(_03727_),
    .ZN(_04052_));
 OAI21_X1 _13145_ (.A(_03500_),
    .B1(_03783_),
    .B2(_03711_),
    .ZN(_04053_));
 NOR2_X1 _13146_ (.A1(_03739_),
    .A2(_03745_),
    .ZN(_04054_));
 NAND4_X1 _13147_ (.A1(_03883_),
    .A2(_03741_),
    .A3(_03715_),
    .A4(_04054_),
    .ZN(_04055_));
 AOI21_X1 _13148_ (.A(_04052_),
    .B1(_04053_),
    .B2(_04055_),
    .ZN(_04056_));
 AOI21_X2 _13149_ (.A(_04049_),
    .B1(_04051_),
    .B2(_04056_),
    .ZN(_04057_));
 OR4_X1 _13150_ (.A1(_03734_),
    .A2(_03735_),
    .A3(_04048_),
    .A4(_03960_),
    .ZN(_04058_));
 NAND2_X1 _13151_ (.A1(_04048_),
    .A2(_03960_),
    .ZN(_04059_));
 AND3_X1 _13152_ (.A1(net376),
    .A2(_03650_),
    .A3(_03679_),
    .ZN(_04060_));
 OAI211_X2 _13153_ (.A(_04058_),
    .B(_04059_),
    .C1(_04060_),
    .C2(_04049_),
    .ZN(_04061_));
 NOR3_X2 _13154_ (.A1(_04050_),
    .A2(_04057_),
    .A3(_04061_),
    .ZN(_04062_));
 NAND2_X2 _13155_ (.A1(net375),
    .A2(_04062_),
    .ZN(_04063_));
 NAND3_X2 _13156_ (.A1(_03957_),
    .A2(_03929_),
    .A3(_03932_),
    .ZN(_04064_));
 AOI21_X4 _13157_ (.A(_04064_),
    .B1(_03788_),
    .B2(net1),
    .ZN(_04065_));
 XOR2_X2 _13158_ (.A(_03959_),
    .B(_04065_),
    .Z(_04066_));
 AOI21_X4 _13159_ (.A(_04047_),
    .B1(_04063_),
    .B2(_04066_),
    .ZN(_04067_));
 NAND2_X2 _13160_ (.A1(_04032_),
    .A2(_04033_),
    .ZN(_04068_));
 NAND3_X4 _13161_ (.A1(_04038_),
    .A2(_04067_),
    .A3(_04068_),
    .ZN(_04069_));
 NOR3_X4 _13162_ (.A1(_04025_),
    .A2(_04028_),
    .A3(_04026_),
    .ZN(_04070_));
 NOR2_X1 _13163_ (.A1(_03503_),
    .A2(_03967_),
    .ZN(_04071_));
 NOR2_X1 _13164_ (.A1(net5),
    .A2(_04071_),
    .ZN(_04072_));
 XNOR2_X2 _13165_ (.A(_04044_),
    .B(_03932_),
    .ZN(_04073_));
 AOI21_X2 _13166_ (.A(_04073_),
    .B1(_03970_),
    .B2(_03967_),
    .ZN(_04074_));
 NOR2_X1 _13167_ (.A1(_03973_),
    .A2(_04074_),
    .ZN(_04075_));
 NAND2_X1 _13168_ (.A1(_03978_),
    .A2(_03980_),
    .ZN(_04076_));
 AOI21_X2 _13169_ (.A(_04072_),
    .B1(_04075_),
    .B2(_04076_),
    .ZN(_04077_));
 OAI21_X1 _13170_ (.A(net5),
    .B1(_03973_),
    .B2(_04074_),
    .ZN(_04078_));
 NAND3_X2 _13171_ (.A1(_03986_),
    .A2(_04062_),
    .A3(_04078_),
    .ZN(_04079_));
 NOR3_X4 _13172_ (.A1(_03503_),
    .A2(_03875_),
    .A3(_03920_),
    .ZN(_04080_));
 AOI21_X4 _13173_ (.A(_03970_),
    .B1(_03788_),
    .B2(net1),
    .ZN(_04081_));
 NOR3_X4 _13174_ (.A1(_03978_),
    .A2(_04080_),
    .A3(_04081_),
    .ZN(_04082_));
 NOR3_X2 _13175_ (.A1(_04077_),
    .A2(_04079_),
    .A3(_04082_),
    .ZN(_04083_));
 NOR2_X4 _13176_ (.A1(_04070_),
    .A2(_04083_),
    .ZN(_04084_));
 INV_X1 _13177_ (.A(_09228_),
    .ZN(_04085_));
 CLKBUF_X2 _13178_ (.A(_09229_),
    .Z(_04086_));
 INV_X1 _13179_ (.A(_04086_),
    .ZN(_04087_));
 INV_X2 _13180_ (.A(_04019_),
    .ZN(_04088_));
 AOI21_X4 _13181_ (.A(_09231_),
    .B1(_04088_),
    .B2(_04005_),
    .ZN(_04089_));
 OAI21_X4 _13182_ (.A(_04085_),
    .B1(_04087_),
    .B2(_04089_),
    .ZN(_04090_));
 INV_X4 _13183_ (.A(_04090_),
    .ZN(_04091_));
 XNOR2_X2 _13184_ (.A(_03977_),
    .B(_03965_),
    .ZN(_04092_));
 NAND2_X1 _13185_ (.A1(_04091_),
    .A2(_04092_),
    .ZN(_04093_));
 NAND2_X1 _13186_ (.A1(_03790_),
    .A2(_04091_),
    .ZN(_04094_));
 MUX2_X2 _13187_ (.A(_04093_),
    .B(_04094_),
    .S(_04070_),
    .Z(_04095_));
 OR4_X4 _13188_ (.A1(_04095_),
    .A2(_04036_),
    .A3(_04084_),
    .A4(_04069_),
    .ZN(_04096_));
 AND3_X1 _13189_ (.A1(_03789_),
    .A2(_03862_),
    .A3(_03905_),
    .ZN(_04097_));
 XNOR2_X2 _13190_ (.A(_03722_),
    .B(_04097_),
    .ZN(_04098_));
 AND4_X2 _13191_ (.A1(_03911_),
    .A2(_03909_),
    .A3(_04023_),
    .A4(_04024_),
    .ZN(_04099_));
 NAND3_X2 _13192_ (.A1(_03989_),
    .A2(_04098_),
    .A3(_04099_),
    .ZN(_04100_));
 XOR2_X2 _13193_ (.A(_03722_),
    .B(_04097_),
    .Z(_04101_));
 AND3_X1 _13194_ (.A1(_03989_),
    .A2(_04101_),
    .A3(_04099_),
    .ZN(_04102_));
 BUF_X4 _13195_ (.A(_04102_),
    .Z(_04103_));
 OAI211_X4 _13196_ (.A(_03990_),
    .B(_04100_),
    .C1(_04103_),
    .C2(_04098_),
    .ZN(_04104_));
 NAND3_X1 _13197_ (.A1(_03861_),
    .A2(_03867_),
    .A3(_03881_),
    .ZN(_04105_));
 NOR2_X1 _13198_ (.A1(_03900_),
    .A2(_03902_),
    .ZN(_04106_));
 XNOR2_X2 _13199_ (.A(_03959_),
    .B(_04065_),
    .ZN(_04107_));
 OR3_X2 _13200_ (.A1(_04050_),
    .A2(_04057_),
    .A3(_04061_),
    .ZN(_04108_));
 NOR3_X2 _13201_ (.A1(_03908_),
    .A2(_03986_),
    .A3(_04108_),
    .ZN(_04109_));
 AND4_X2 _13202_ (.A1(_03938_),
    .A2(_03955_),
    .A3(_04107_),
    .A4(_04109_),
    .ZN(_04110_));
 NAND4_X2 _13203_ (.A1(_04105_),
    .A2(_04106_),
    .A3(_03926_),
    .A4(_04110_),
    .ZN(_04111_));
 NAND4_X4 _13204_ (.A1(_03938_),
    .A2(_03955_),
    .A3(_04107_),
    .A4(_04109_),
    .ZN(_04112_));
 OAI22_X4 _13205_ (.A1(_03900_),
    .A2(_03902_),
    .B1(_04025_),
    .B2(_04112_),
    .ZN(_04113_));
 OAI211_X2 _13206_ (.A(_04024_),
    .B(_04110_),
    .C1(_04025_),
    .C2(_04026_),
    .ZN(_04114_));
 AOI21_X1 _13207_ (.A(_03911_),
    .B1(_03924_),
    .B2(_03831_),
    .ZN(_04115_));
 OR2_X1 _13208_ (.A1(_03922_),
    .A2(_04115_),
    .ZN(_04116_));
 AOI21_X1 _13209_ (.A(_04116_),
    .B1(_04112_),
    .B2(_03925_),
    .ZN(_04117_));
 AND4_X4 _13210_ (.A1(_04111_),
    .A2(_04113_),
    .A3(_04114_),
    .A4(_04117_),
    .ZN(_04118_));
 NAND2_X1 _13211_ (.A1(_03722_),
    .A2(_03856_),
    .ZN(_04119_));
 AOI211_X2 _13212_ (.A(_03833_),
    .B(_04119_),
    .C1(net1),
    .C2(_03788_),
    .ZN(_04120_));
 XOR2_X2 _13213_ (.A(_03834_),
    .B(_04120_),
    .Z(_04121_));
 AND3_X1 _13214_ (.A1(_03867_),
    .A2(_03881_),
    .A3(_04121_),
    .ZN(_04122_));
 NAND4_X2 _13215_ (.A1(_03989_),
    .A2(_04101_),
    .A3(_04099_),
    .A4(_04122_),
    .ZN(_04123_));
 XNOR2_X2 _13216_ (.A(_03834_),
    .B(_04120_),
    .ZN(_04124_));
 NAND3_X1 _13217_ (.A1(_03867_),
    .A2(_03881_),
    .A3(_04124_),
    .ZN(_04125_));
 OAI211_X4 _13218_ (.A(_03990_),
    .B(_04123_),
    .C1(_04125_),
    .C2(_04103_),
    .ZN(_04126_));
 OAI21_X1 _13219_ (.A(_04110_),
    .B1(_04025_),
    .B2(_04026_),
    .ZN(_04127_));
 XNOR2_X1 _13220_ (.A(_03680_),
    .B(_03903_),
    .ZN(_04128_));
 AOI21_X2 _13221_ (.A(_04128_),
    .B1(_03788_),
    .B2(_03901_),
    .ZN(_04129_));
 OAI21_X1 _13222_ (.A(_04129_),
    .B1(_04030_),
    .B2(_04028_),
    .ZN(_04130_));
 AND2_X1 _13223_ (.A1(_04127_),
    .A2(_04130_),
    .ZN(_04131_));
 BUF_X4 _13224_ (.A(_04131_),
    .Z(_04132_));
 NAND4_X4 _13225_ (.A1(_04104_),
    .A2(_04118_),
    .A3(_04126_),
    .A4(_04132_),
    .ZN(_04133_));
 OR2_X4 _13226_ (.A1(_04096_),
    .A2(_04133_),
    .ZN(_04134_));
 BUF_X8 _13227_ (.A(_04134_),
    .Z(_04135_));
 MUX2_X1 _13228_ (.A(_09230_),
    .B(_04020_),
    .S(net40),
    .Z(_09259_));
 INV_X1 _13229_ (.A(_09255_),
    .ZN(_04136_));
 INV_X1 _13230_ (.A(_09257_),
    .ZN(_04137_));
 INV_X1 _13231_ (.A(_09251_),
    .ZN(_04138_));
 INV_X1 _13232_ (.A(_09245_),
    .ZN(_04139_));
 OAI21_X2 _13233_ (.A(_09246_),
    .B1(_09240_),
    .B2(_09239_),
    .ZN(_04140_));
 NAND2_X2 _13234_ (.A1(_04140_),
    .A2(_04139_),
    .ZN(_04141_));
 AOI21_X4 _13235_ (.A(_09242_),
    .B1(_09243_),
    .B2(_04141_),
    .ZN(_04142_));
 INV_X1 _13236_ (.A(_09252_),
    .ZN(_04143_));
 OAI21_X4 _13237_ (.A(_04138_),
    .B1(_04142_),
    .B2(_04143_),
    .ZN(_04144_));
 AOI21_X4 _13238_ (.A(_09248_),
    .B1(_09249_),
    .B2(_04144_),
    .ZN(_04145_));
 INV_X1 _13239_ (.A(_09258_),
    .ZN(_04146_));
 OAI21_X4 _13240_ (.A(_04137_),
    .B1(_04145_),
    .B2(_04146_),
    .ZN(_04147_));
 XNOR2_X1 _13241_ (.A(_04136_),
    .B(_04147_),
    .ZN(_04148_));
 NOR2_X1 _13242_ (.A1(_09126_),
    .A2(_03315_),
    .ZN(_09142_));
 OR3_X1 _13243_ (.A1(_09147_),
    .A2(_09144_),
    .A3(_09146_),
    .ZN(_04149_));
 AND2_X1 _13244_ (.A1(_03289_),
    .A2(_04149_),
    .ZN(_04150_));
 MUX2_X1 _13245_ (.A(_09142_),
    .B(_04150_),
    .S(_03354_),
    .Z(_09162_));
 INV_X1 _13246_ (.A(_09166_),
    .ZN(_04151_));
 NAND2_X1 _13247_ (.A1(_04151_),
    .A2(_03371_),
    .ZN(_04152_));
 XOR2_X1 _13248_ (.A(_09164_),
    .B(_04152_),
    .Z(_04153_));
 MUX2_X1 _13249_ (.A(_09162_),
    .B(_04153_),
    .S(_03524_),
    .Z(_09180_));
 XNOR2_X1 _13250_ (.A(_03545_),
    .B(_03795_),
    .ZN(_04154_));
 MUX2_X1 _13251_ (.A(_09180_),
    .B(_04154_),
    .S(_03791_),
    .Z(_09209_));
 XOR2_X1 _13252_ (.A(_09211_),
    .B(_03817_),
    .Z(_04155_));
 MUX2_X1 _13253_ (.A(_09209_),
    .B(_04155_),
    .S(_03991_),
    .Z(_09233_));
 INV_X1 _13254_ (.A(_09216_),
    .ZN(_04156_));
 INV_X1 _13255_ (.A(_09222_),
    .ZN(_04157_));
 OAI21_X1 _13256_ (.A(_09223_),
    .B1(_09225_),
    .B2(_04008_),
    .ZN(_04158_));
 AOI21_X1 _13257_ (.A(_04012_),
    .B1(_04157_),
    .B2(_04158_),
    .ZN(_04159_));
 NOR2_X1 _13258_ (.A1(_09219_),
    .A2(_04159_),
    .ZN(_04160_));
 INV_X1 _13259_ (.A(_04014_),
    .ZN(_04161_));
 OAI21_X1 _13260_ (.A(_04156_),
    .B1(_04160_),
    .B2(_04161_),
    .ZN(_04162_));
 AOI21_X2 _13261_ (.A(_09237_),
    .B1(_04162_),
    .B2(_09238_),
    .ZN(_04163_));
 XNOR2_X1 _13262_ (.A(_04018_),
    .B(_04163_),
    .ZN(_04164_));
 MUX2_X1 _13263_ (.A(_09233_),
    .B(_04164_),
    .S(net40),
    .Z(_09253_));
 BUF_X8 _13264_ (.A(_04070_),
    .Z(_04165_));
 NOR2_X1 _13265_ (.A1(_04063_),
    .A2(_04165_),
    .ZN(_04166_));
 NAND2_X1 _13266_ (.A1(_03986_),
    .A2(_04108_),
    .ZN(_04167_));
 NAND3_X1 _13267_ (.A1(_09186_),
    .A2(net1),
    .A3(_03788_),
    .ZN(_04168_));
 OAI21_X1 _13268_ (.A(_03980_),
    .B1(_03920_),
    .B2(_03875_),
    .ZN(_04169_));
 AOI21_X2 _13269_ (.A(_03978_),
    .B1(_04168_),
    .B2(_04169_),
    .ZN(_04170_));
 NOR3_X2 _13270_ (.A1(net6),
    .A2(_04080_),
    .A3(_04081_),
    .ZN(_04171_));
 OAI211_X2 _13271_ (.A(_04091_),
    .B(_04092_),
    .C1(_04170_),
    .C2(_04171_),
    .ZN(_04172_));
 NOR2_X2 _13272_ (.A1(_04080_),
    .A2(_04081_),
    .ZN(_04173_));
 INV_X1 _13273_ (.A(_03540_),
    .ZN(_09189_));
 XNOR2_X1 _13274_ (.A(_09202_),
    .B(_03965_),
    .ZN(_04174_));
 NOR2_X1 _13275_ (.A1(net6),
    .A2(_04174_),
    .ZN(_04175_));
 INV_X1 _13276_ (.A(_04175_),
    .ZN(_04176_));
 NAND2_X1 _13277_ (.A1(_09189_),
    .A2(_04176_),
    .ZN(_04177_));
 NAND4_X1 _13278_ (.A1(_03555_),
    .A2(_03558_),
    .A3(_03563_),
    .A4(_04176_),
    .ZN(_04178_));
 MUX2_X1 _13279_ (.A(_04177_),
    .B(_04178_),
    .S(net5),
    .Z(_04179_));
 NAND3_X1 _13280_ (.A1(_04091_),
    .A2(_04173_),
    .A3(_04179_),
    .ZN(_04180_));
 OAI21_X2 _13281_ (.A(_04172_),
    .B1(_04180_),
    .B2(_03990_),
    .ZN(_04181_));
 AOI21_X1 _13282_ (.A(_04167_),
    .B1(_04181_),
    .B2(_04078_),
    .ZN(_04182_));
 OR2_X1 _13283_ (.A1(_04166_),
    .A2(_04182_),
    .ZN(_04183_));
 NOR4_X4 _13284_ (.A1(_04036_),
    .A2(_04069_),
    .A3(_04084_),
    .A4(_04095_),
    .ZN(_04184_));
 BUF_X4 _13285_ (.A(_04184_),
    .Z(_04185_));
 AND2_X2 _13286_ (.A1(_04104_),
    .A2(_04118_),
    .ZN(_04186_));
 AND2_X2 _13287_ (.A1(_04126_),
    .A2(_04132_),
    .ZN(_04187_));
 NAND3_X2 _13288_ (.A1(_04185_),
    .A2(_04186_),
    .A3(_04187_),
    .ZN(_04188_));
 OAI21_X1 _13289_ (.A(_04092_),
    .B1(_04170_),
    .B2(_04171_),
    .ZN(_04189_));
 NOR2_X1 _13290_ (.A1(_04090_),
    .A2(_04189_),
    .ZN(_04190_));
 INV_X1 _13291_ (.A(_04180_),
    .ZN(_04191_));
 AOI21_X2 _13292_ (.A(_04190_),
    .B1(_04191_),
    .B2(net408),
    .ZN(_04192_));
 NOR2_X1 _13293_ (.A1(net14),
    .A2(_04192_),
    .ZN(_04193_));
 AND2_X1 _13294_ (.A1(_04172_),
    .A2(_04180_),
    .ZN(_04194_));
 OR2_X1 _13295_ (.A1(_04079_),
    .A2(_04172_),
    .ZN(_04195_));
 AOI21_X2 _13296_ (.A(_04194_),
    .B1(_04195_),
    .B2(_03990_),
    .ZN(_04196_));
 AOI221_X2 _13297_ (.A(_04183_),
    .B1(_04188_),
    .B2(_04193_),
    .C1(_04134_),
    .C2(_04196_),
    .ZN(_04197_));
 NOR2_X2 _13298_ (.A1(_03974_),
    .A2(_04073_),
    .ZN(_04198_));
 AOI22_X4 _13299_ (.A1(net426),
    .A2(net14),
    .B1(_04198_),
    .B2(net23),
    .ZN(_04199_));
 AND3_X2 _13300_ (.A1(_04185_),
    .A2(_04186_),
    .A3(_04187_),
    .ZN(_04200_));
 NAND2_X1 _13301_ (.A1(net5),
    .A2(_03972_),
    .ZN(_04201_));
 XOR2_X2 _13302_ (.A(_03931_),
    .B(_04201_),
    .Z(_04202_));
 OAI21_X1 _13303_ (.A(_03978_),
    .B1(_04080_),
    .B2(_04081_),
    .ZN(_04203_));
 NAND2_X1 _13304_ (.A1(net6),
    .A2(_04173_),
    .ZN(_04204_));
 OAI21_X2 _13305_ (.A(_04203_),
    .B1(_04204_),
    .B2(_04165_),
    .ZN(_04205_));
 OR2_X1 _13306_ (.A1(_04202_),
    .A2(_04205_),
    .ZN(_04206_));
 NAND3_X1 _13307_ (.A1(_04086_),
    .A2(_04005_),
    .A3(_04018_),
    .ZN(_04207_));
 NOR2_X2 _13308_ (.A1(_04163_),
    .A2(_04207_),
    .ZN(_04208_));
 AOI21_X1 _13309_ (.A(_09231_),
    .B1(_09234_),
    .B2(_04005_),
    .ZN(_04209_));
 INV_X1 _13310_ (.A(_04209_),
    .ZN(_04210_));
 AOI21_X2 _13311_ (.A(_09228_),
    .B1(_04086_),
    .B2(_04210_),
    .ZN(_04211_));
 INV_X1 _13312_ (.A(_04211_),
    .ZN(_04212_));
 NOR2_X1 _13313_ (.A1(_04208_),
    .A2(_04212_),
    .ZN(_04213_));
 NAND2_X1 _13314_ (.A1(_04092_),
    .A2(_04213_),
    .ZN(_04214_));
 NAND2_X1 _13315_ (.A1(_03790_),
    .A2(_04213_),
    .ZN(_04215_));
 MUX2_X2 _13316_ (.A(_04214_),
    .B(_04215_),
    .S(_04070_),
    .Z(_04216_));
 NOR3_X4 _13317_ (.A1(_04200_),
    .A2(_04206_),
    .A3(_04216_),
    .ZN(_04217_));
 XOR2_X2 _13318_ (.A(_04199_),
    .B(_04217_),
    .Z(_04218_));
 OR4_X2 _13319_ (.A1(_04026_),
    .A2(_04025_),
    .A3(_04028_),
    .A4(_04215_),
    .ZN(_04219_));
 OAI21_X4 _13320_ (.A(_04219_),
    .B1(_04214_),
    .B2(_04070_),
    .ZN(_04220_));
 NAND2_X1 _13321_ (.A1(net8),
    .A2(_04173_),
    .ZN(_04221_));
 OAI221_X2 _13322_ (.A(_04202_),
    .B1(_04220_),
    .B2(_04192_),
    .C1(_04221_),
    .C2(_03978_),
    .ZN(_04222_));
 INV_X1 _13323_ (.A(_04202_),
    .ZN(_04223_));
 NAND4_X1 _13324_ (.A1(net6),
    .A2(net8),
    .A3(_04173_),
    .A4(_04223_),
    .ZN(_04224_));
 NOR3_X1 _13325_ (.A1(net408),
    .A2(_04204_),
    .A3(_04223_),
    .ZN(_04225_));
 NOR2_X1 _13326_ (.A1(_04202_),
    .A2(_04203_),
    .ZN(_04226_));
 OAI21_X1 _13327_ (.A(_04216_),
    .B1(_04225_),
    .B2(_04226_),
    .ZN(_04227_));
 NAND3_X2 _13328_ (.A1(_04222_),
    .A2(_04224_),
    .A3(_04227_),
    .ZN(_04228_));
 MUX2_X2 _13329_ (.A(_09200_),
    .B(_04174_),
    .S(net8),
    .Z(_04229_));
 XNOR2_X2 _13330_ (.A(_04090_),
    .B(_04229_),
    .ZN(_04230_));
 INV_X2 _13331_ (.A(_09260_),
    .ZN(_04231_));
 INV_X1 _13332_ (.A(_09261_),
    .ZN(_04232_));
 AOI21_X4 _13333_ (.A(_09254_),
    .B1(_09255_),
    .B2(_04147_),
    .ZN(_04233_));
 OAI21_X4 _13334_ (.A(_04231_),
    .B1(_04233_),
    .B2(_04232_),
    .ZN(_04234_));
 INV_X1 _13335_ (.A(_09234_),
    .ZN(_04235_));
 INV_X1 _13336_ (.A(_04018_),
    .ZN(_04236_));
 OAI21_X1 _13337_ (.A(_04235_),
    .B1(_04163_),
    .B2(_04236_),
    .ZN(_04237_));
 AOI21_X2 _13338_ (.A(_09231_),
    .B1(_04237_),
    .B2(_04005_),
    .ZN(_04238_));
 XNOR2_X2 _13339_ (.A(_04086_),
    .B(_04238_),
    .ZN(_04239_));
 NOR3_X2 _13340_ (.A1(_04230_),
    .A2(_04234_),
    .A3(_04239_),
    .ZN(_04240_));
 NOR3_X4 _13341_ (.A1(_04234_),
    .A2(_03822_),
    .A3(net408),
    .ZN(_04241_));
 NOR3_X4 _13342_ (.A1(_04234_),
    .A2(net8),
    .A3(_09203_),
    .ZN(_04242_));
 NOR2_X4 _13343_ (.A1(_04241_),
    .A2(_04242_),
    .ZN(_04243_));
 NOR2_X4 _13344_ (.A1(_04243_),
    .A2(_04229_),
    .ZN(_04244_));
 NOR2_X4 _13345_ (.A1(_04096_),
    .A2(_04133_),
    .ZN(_04245_));
 AOI21_X4 _13346_ (.A(_04240_),
    .B1(_04244_),
    .B2(_04245_),
    .ZN(_04246_));
 NOR2_X4 _13347_ (.A1(_04228_),
    .A2(_04246_),
    .ZN(_04247_));
 NAND3_X4 _13348_ (.A1(_04197_),
    .A2(_04218_),
    .A3(_04247_),
    .ZN(_04248_));
 NAND2_X1 _13349_ (.A1(_03831_),
    .A2(_03924_),
    .ZN(_04249_));
 OAI211_X4 _13350_ (.A(_04024_),
    .B(_04110_),
    .C1(_04025_),
    .C2(_04026_),
    .ZN(_04250_));
 AOI21_X2 _13351_ (.A(_03896_),
    .B1(_04249_),
    .B2(_04250_),
    .ZN(_04251_));
 XNOR2_X2 _13352_ (.A(_03911_),
    .B(_04251_),
    .ZN(_04252_));
 OAI21_X4 _13353_ (.A(_04027_),
    .B1(_04034_),
    .B2(_04035_),
    .ZN(_04253_));
 INV_X1 _13354_ (.A(_04129_),
    .ZN(_04254_));
 NOR4_X1 _13355_ (.A1(_04077_),
    .A2(_04030_),
    .A3(_04079_),
    .A4(_04082_),
    .ZN(_04255_));
 OAI21_X1 _13356_ (.A(_04254_),
    .B1(_04255_),
    .B2(net12),
    .ZN(_04256_));
 NOR3_X2 _13357_ (.A1(_04253_),
    .A2(_04069_),
    .A3(_04256_),
    .ZN(_04257_));
 NAND2_X1 _13358_ (.A1(_04092_),
    .A2(_04211_),
    .ZN(_04258_));
 NAND2_X1 _13359_ (.A1(_03790_),
    .A2(_04211_),
    .ZN(_04259_));
 MUX2_X1 _13360_ (.A(_04258_),
    .B(_04259_),
    .S(_04070_),
    .Z(_04260_));
 NAND2_X2 _13361_ (.A1(_03925_),
    .A2(_04112_),
    .ZN(_04261_));
 XNOR2_X2 _13362_ (.A(_04021_),
    .B(_03921_),
    .ZN(_04262_));
 NAND3_X2 _13363_ (.A1(_04261_),
    .A2(_04250_),
    .A3(_04262_),
    .ZN(_04263_));
 NOR2_X1 _13364_ (.A1(net6),
    .A2(_03970_),
    .ZN(_04264_));
 OAI33_X1 _13365_ (.A1(_03875_),
    .A2(_03920_),
    .A3(_04071_),
    .B1(_04074_),
    .B2(_04264_),
    .B3(_03973_),
    .ZN(_04265_));
 NAND2_X1 _13366_ (.A1(_03790_),
    .A2(_04265_),
    .ZN(_04266_));
 NOR4_X4 _13367_ (.A1(_04026_),
    .A2(_04025_),
    .A3(_04028_),
    .A4(_04266_),
    .ZN(_04267_));
 NOR2_X2 _13368_ (.A1(_04079_),
    .A2(_04189_),
    .ZN(_04268_));
 OR2_X1 _13369_ (.A1(_04267_),
    .A2(_04268_),
    .ZN(_04269_));
 AOI211_X2 _13370_ (.A(_04260_),
    .B(_04263_),
    .C1(_04269_),
    .C2(_04208_),
    .ZN(_04270_));
 OAI211_X2 _13371_ (.A(_04257_),
    .B(_04270_),
    .C1(_04096_),
    .C2(_04133_),
    .ZN(_04271_));
 XNOR2_X2 _13372_ (.A(_04252_),
    .B(_04271_),
    .ZN(_04272_));
 INV_X1 _13373_ (.A(_04263_),
    .ZN(_04273_));
 XOR2_X2 _13374_ (.A(_04250_),
    .B(_04262_),
    .Z(_04274_));
 NAND4_X1 _13375_ (.A1(_04014_),
    .A2(_04008_),
    .A3(_09220_),
    .A4(_09223_),
    .ZN(_04275_));
 OR4_X1 _13376_ (.A1(_04016_),
    .A2(_01097_),
    .A3(_04207_),
    .A4(_04275_),
    .ZN(_04276_));
 INV_X1 _13377_ (.A(_04276_),
    .ZN(_04277_));
 AND3_X1 _13378_ (.A1(_04067_),
    .A2(_04068_),
    .A3(_04277_),
    .ZN(_04278_));
 OAI211_X4 _13379_ (.A(_04038_),
    .B(_04278_),
    .C1(_04268_),
    .C2(_04267_),
    .ZN(_04279_));
 NAND4_X4 _13380_ (.A1(_04104_),
    .A2(_04118_),
    .A3(_04126_),
    .A4(_04279_),
    .ZN(_04280_));
 NAND3_X4 _13381_ (.A1(_04185_),
    .A2(_04132_),
    .A3(_04280_),
    .ZN(_04281_));
 MUX2_X1 _13382_ (.A(_04273_),
    .B(_04274_),
    .S(_04281_),
    .Z(_04282_));
 NAND2_X2 _13383_ (.A1(_04261_),
    .A2(_04250_),
    .ZN(_04283_));
 INV_X1 _13384_ (.A(_04274_),
    .ZN(_04284_));
 NAND2_X1 _13385_ (.A1(_04283_),
    .A2(_04284_),
    .ZN(_04285_));
 OR4_X2 _13386_ (.A1(_04253_),
    .A2(_04069_),
    .A3(_04216_),
    .A4(_04256_),
    .ZN(_04286_));
 OR3_X1 _13387_ (.A1(_04200_),
    .A2(_04285_),
    .A3(_04286_),
    .ZN(_04287_));
 AND2_X1 _13388_ (.A1(_04261_),
    .A2(_04250_),
    .ZN(_04288_));
 OAI21_X1 _13389_ (.A(_04288_),
    .B1(_04200_),
    .B2(_04286_),
    .ZN(_04289_));
 AOI211_X4 _13390_ (.A(_04272_),
    .B(_04282_),
    .C1(_04287_),
    .C2(_04289_),
    .ZN(_04290_));
 NAND3_X2 _13391_ (.A1(net12),
    .A2(_04101_),
    .A3(_04099_),
    .ZN(_04291_));
 AOI21_X1 _13392_ (.A(net408),
    .B1(_04291_),
    .B2(_04101_),
    .ZN(_04292_));
 AND2_X1 _13393_ (.A1(_04292_),
    .A2(_04100_),
    .ZN(_04293_));
 AOI21_X1 _13394_ (.A(_04293_),
    .B1(_04187_),
    .B2(_04185_),
    .ZN(_04294_));
 NAND3_X1 _13395_ (.A1(_04118_),
    .A2(_04220_),
    .A3(_04257_),
    .ZN(_04295_));
 MUX2_X2 _13396_ (.A(_04294_),
    .B(_04293_),
    .S(_04295_),
    .Z(_04296_));
 NAND2_X2 _13397_ (.A1(_04111_),
    .A2(_04113_),
    .ZN(_04297_));
 NOR2_X1 _13398_ (.A1(_04116_),
    .A2(_04283_),
    .ZN(_04298_));
 NAND4_X4 _13399_ (.A1(_04185_),
    .A2(_04298_),
    .A3(_04132_),
    .A4(_04280_),
    .ZN(_04299_));
 XNOR2_X2 _13400_ (.A(_04297_),
    .B(_04299_),
    .ZN(_04300_));
 NOR2_X4 _13401_ (.A1(_04296_),
    .A2(_04300_),
    .ZN(_04301_));
 NAND4_X4 _13402_ (.A1(_03910_),
    .A2(_03926_),
    .A3(_03938_),
    .A4(_03955_),
    .ZN(_04302_));
 NOR3_X2 _13403_ (.A1(_03951_),
    .A2(_03964_),
    .A3(_03986_),
    .ZN(_04303_));
 AOI21_X4 _13404_ (.A(_04047_),
    .B1(_04302_),
    .B2(_04303_),
    .ZN(_04304_));
 NOR2_X1 _13405_ (.A1(_04196_),
    .A2(_04304_),
    .ZN(_04305_));
 OAI33_X1 _13406_ (.A1(_04026_),
    .A2(_04025_),
    .A3(_04028_),
    .B1(_04077_),
    .B2(_04079_),
    .B3(_04082_),
    .ZN(_04306_));
 NAND3_X1 _13407_ (.A1(_04306_),
    .A2(_04220_),
    .A3(_04304_),
    .ZN(_04307_));
 AND2_X1 _13408_ (.A1(_04066_),
    .A2(_04063_),
    .ZN(_04308_));
 AOI21_X2 _13409_ (.A(_04308_),
    .B1(_04302_),
    .B2(_03987_),
    .ZN(_04309_));
 INV_X1 _13410_ (.A(_04309_),
    .ZN(_04310_));
 AOI21_X2 _13411_ (.A(_04305_),
    .B1(_04307_),
    .B2(_04310_),
    .ZN(_04311_));
 NAND2_X1 _13412_ (.A1(_04196_),
    .A2(_04304_),
    .ZN(_04312_));
 NOR2_X1 _13413_ (.A1(_04084_),
    .A2(_04216_),
    .ZN(_04313_));
 MUX2_X1 _13414_ (.A(_04312_),
    .B(_04310_),
    .S(_04313_),
    .Z(_04314_));
 OAI21_X4 _13415_ (.A(_04311_),
    .B1(_04314_),
    .B2(_04245_),
    .ZN(_04315_));
 NOR3_X2 _13416_ (.A1(_04069_),
    .A2(_04084_),
    .A3(_04216_),
    .ZN(_04316_));
 OAI21_X2 _13417_ (.A(_04316_),
    .B1(_04133_),
    .B2(_04096_),
    .ZN(_04317_));
 NOR4_X2 _13418_ (.A1(_04253_),
    .A2(_04069_),
    .A3(_04084_),
    .A4(_04095_),
    .ZN(_04318_));
 NAND2_X1 _13419_ (.A1(_04031_),
    .A2(_04091_),
    .ZN(_04319_));
 OAI21_X2 _13420_ (.A(_04318_),
    .B1(_04319_),
    .B2(_04133_),
    .ZN(_04320_));
 AND2_X1 _13421_ (.A1(_04067_),
    .A2(_04306_),
    .ZN(_04321_));
 AOI22_X4 _13422_ (.A1(_04038_),
    .A2(_04068_),
    .B1(_04220_),
    .B2(_04321_),
    .ZN(_04322_));
 OR3_X1 _13423_ (.A1(_04069_),
    .A2(_04084_),
    .A3(_04095_),
    .ZN(_04323_));
 AOI21_X2 _13424_ (.A(_04322_),
    .B1(_04323_),
    .B2(_04253_),
    .ZN(_04324_));
 NAND3_X4 _13425_ (.A1(_04317_),
    .A2(_04320_),
    .A3(_04324_),
    .ZN(_04325_));
 OR2_X1 _13426_ (.A1(_04185_),
    .A2(_04132_),
    .ZN(_04326_));
 NOR4_X1 _13427_ (.A1(_04253_),
    .A2(_04069_),
    .A3(_04084_),
    .A4(_04216_),
    .ZN(_04327_));
 MUX2_X1 _13428_ (.A(_04027_),
    .B(net12),
    .S(_04030_),
    .Z(_04328_));
 OR2_X1 _13429_ (.A1(_04327_),
    .A2(_04328_),
    .ZN(_04329_));
 NAND3_X2 _13430_ (.A1(_04281_),
    .A2(_04326_),
    .A3(_04329_),
    .ZN(_04330_));
 NOR3_X4 _13431_ (.A1(_04315_),
    .A2(_04325_),
    .A3(_04330_),
    .ZN(_04331_));
 NOR2_X1 _13432_ (.A1(_04165_),
    .A2(_04121_),
    .ZN(_04332_));
 NOR3_X1 _13433_ (.A1(_03880_),
    .A2(_04291_),
    .A3(_04332_),
    .ZN(_04333_));
 NAND2_X1 _13434_ (.A1(_04126_),
    .A2(_04279_),
    .ZN(_04334_));
 NAND4_X4 _13435_ (.A1(_04185_),
    .A2(_04186_),
    .A3(_04132_),
    .A4(_04334_),
    .ZN(_04335_));
 NOR3_X1 _13436_ (.A1(_03880_),
    .A2(_04103_),
    .A3(_04121_),
    .ZN(_04336_));
 NOR3_X1 _13437_ (.A1(_03880_),
    .A2(_04103_),
    .A3(_04124_),
    .ZN(_04337_));
 AND3_X1 _13438_ (.A1(_04185_),
    .A2(_04186_),
    .A3(_04132_),
    .ZN(_04338_));
 AOI221_X2 _13439_ (.A(_04333_),
    .B1(_04335_),
    .B2(_04336_),
    .C1(_04337_),
    .C2(_04338_),
    .ZN(_04339_));
 NAND3_X2 _13440_ (.A1(_03867_),
    .A2(_04103_),
    .A3(_04124_),
    .ZN(_04340_));
 OAI21_X2 _13441_ (.A(_03873_),
    .B1(_03880_),
    .B2(_04340_),
    .ZN(_04341_));
 AOI21_X1 _13442_ (.A(_03880_),
    .B1(net8),
    .B2(_04103_),
    .ZN(_04342_));
 NAND2_X1 _13443_ (.A1(_03867_),
    .A2(_04342_),
    .ZN(_04343_));
 OR3_X1 _13444_ (.A1(_03867_),
    .A2(_03880_),
    .A3(_04291_),
    .ZN(_04344_));
 AOI21_X2 _13445_ (.A(_04286_),
    .B1(_04343_),
    .B2(_04344_),
    .ZN(_04345_));
 NAND3_X2 _13446_ (.A1(_04104_),
    .A2(_04118_),
    .A3(_04124_),
    .ZN(_04346_));
 AOI21_X2 _13447_ (.A(_04346_),
    .B1(_04187_),
    .B2(_04185_),
    .ZN(_04347_));
 AOI21_X4 _13448_ (.A(_04341_),
    .B1(_04345_),
    .B2(_04347_),
    .ZN(_04348_));
 AOI211_X2 _13449_ (.A(_04286_),
    .B(_04346_),
    .C1(_04184_),
    .C2(_04187_),
    .ZN(_04349_));
 NAND2_X1 _13450_ (.A1(_04103_),
    .A2(_04124_),
    .ZN(_04350_));
 NOR2_X1 _13451_ (.A1(_04165_),
    .A2(_04350_),
    .ZN(_04351_));
 MUX2_X1 _13452_ (.A(_04350_),
    .B(_04351_),
    .S(_03867_),
    .Z(_04352_));
 XOR2_X2 _13453_ (.A(_04349_),
    .B(_04352_),
    .Z(_04353_));
 NOR3_X2 _13454_ (.A1(_04339_),
    .A2(_04348_),
    .A3(_04353_),
    .ZN(_04354_));
 NAND4_X4 _13455_ (.A1(_04290_),
    .A2(_04301_),
    .A3(_04331_),
    .A4(_04354_),
    .ZN(_04355_));
 NOR2_X4 _13456_ (.A1(_04248_),
    .A2(_04355_),
    .ZN(_04356_));
 BUF_X4 _13457_ (.A(_04356_),
    .Z(_04357_));
 MUX2_X2 _13458_ (.A(_04148_),
    .B(_09253_),
    .S(net26),
    .Z(_09279_));
 INV_X1 _13459_ (.A(_04348_),
    .ZN(_04358_));
 NOR2_X2 _13460_ (.A1(_04339_),
    .A2(_04353_),
    .ZN(_04359_));
 NAND4_X2 _13461_ (.A1(_04290_),
    .A2(_04301_),
    .A3(_04358_),
    .A4(_04359_),
    .ZN(_04360_));
 AND4_X1 _13462_ (.A1(_04197_),
    .A2(_04218_),
    .A3(_04247_),
    .A4(_04331_),
    .ZN(_04361_));
 OR2_X2 _13463_ (.A1(_04245_),
    .A2(_04286_),
    .ZN(_04362_));
 OR2_X1 _13464_ (.A1(_04285_),
    .A2(_04362_),
    .ZN(_04363_));
 XNOR2_X1 _13465_ (.A(_04284_),
    .B(_04281_),
    .ZN(_04364_));
 NAND3_X1 _13466_ (.A1(_04288_),
    .A2(_04362_),
    .A3(_04364_),
    .ZN(_04365_));
 NAND2_X1 _13467_ (.A1(_04363_),
    .A2(_04365_),
    .ZN(_04366_));
 NAND3_X1 _13468_ (.A1(_04360_),
    .A2(_04361_),
    .A3(_04366_),
    .ZN(_04367_));
 XNOR2_X2 _13469_ (.A(_04272_),
    .B(_04367_),
    .ZN(_04368_));
 AND2_X1 _13470_ (.A1(_04273_),
    .A2(_04281_),
    .ZN(_04369_));
 NAND4_X4 _13471_ (.A1(_04197_),
    .A2(_04218_),
    .A3(net404),
    .A4(_04331_),
    .ZN(_04370_));
 AND4_X1 _13472_ (.A1(_04290_),
    .A2(_04301_),
    .A3(_04358_),
    .A4(_04359_),
    .ZN(_04371_));
 OAI21_X1 _13473_ (.A(_04369_),
    .B1(_04370_),
    .B2(_04371_),
    .ZN(_04372_));
 INV_X1 _13474_ (.A(_04362_),
    .ZN(_04373_));
 NOR3_X1 _13475_ (.A1(_04263_),
    .A2(_04281_),
    .A3(_04373_),
    .ZN(_04374_));
 OAI21_X1 _13476_ (.A(_04374_),
    .B1(_04370_),
    .B2(_04371_),
    .ZN(_04375_));
 NOR2_X1 _13477_ (.A1(_04166_),
    .A2(_04182_),
    .ZN(_04376_));
 NAND2_X1 _13478_ (.A1(net408),
    .A2(_04181_),
    .ZN(_04377_));
 NOR2_X2 _13479_ (.A1(_04090_),
    .A2(_04229_),
    .ZN(_04378_));
 NAND2_X1 _13480_ (.A1(_04306_),
    .A2(_04378_),
    .ZN(_04379_));
 OAI221_X2 _13481_ (.A(_04376_),
    .B1(_04200_),
    .B2(_04377_),
    .C1(_04245_),
    .C2(_04379_),
    .ZN(_04380_));
 AND3_X1 _13482_ (.A1(_04222_),
    .A2(_04224_),
    .A3(_04227_),
    .ZN(_04381_));
 NOR2_X1 _13483_ (.A1(_04202_),
    .A2(_04205_),
    .ZN(_04382_));
 AOI222_X2 _13484_ (.A1(net426),
    .A2(net14),
    .B1(_04378_),
    .B2(_04382_),
    .C1(_04198_),
    .C2(net23),
    .ZN(_04383_));
 OAI21_X4 _13485_ (.A(_04381_),
    .B1(_04383_),
    .B2(_04245_),
    .ZN(_04384_));
 OAI21_X2 _13486_ (.A(_04378_),
    .B1(_04096_),
    .B2(_04133_),
    .ZN(_04385_));
 NAND2_X1 _13487_ (.A1(_04090_),
    .A2(_04229_),
    .ZN(_04386_));
 NAND2_X4 _13488_ (.A1(_04385_),
    .A2(_04386_),
    .ZN(_04387_));
 NOR4_X4 _13489_ (.A1(_04380_),
    .A2(_04315_),
    .A3(_04384_),
    .A4(_04387_),
    .ZN(_04388_));
 NAND4_X4 _13490_ (.A1(_09227_),
    .A2(_04185_),
    .A3(_04186_),
    .A4(_04187_),
    .ZN(_04389_));
 OAI21_X4 _13491_ (.A(_04239_),
    .B1(_04133_),
    .B2(net407),
    .ZN(_04390_));
 INV_X1 _13492_ (.A(_09254_),
    .ZN(_04391_));
 INV_X1 _13493_ (.A(_09248_),
    .ZN(_04392_));
 AOI21_X1 _13494_ (.A(_09239_),
    .B1(_02103_),
    .B2(_09240_),
    .ZN(_04393_));
 INV_X1 _13495_ (.A(_09246_),
    .ZN(_04394_));
 OAI21_X1 _13496_ (.A(_04139_),
    .B1(_04393_),
    .B2(_04394_),
    .ZN(_04395_));
 AND2_X1 _13497_ (.A1(_09243_),
    .A2(_04395_),
    .ZN(_04396_));
 OR2_X1 _13498_ (.A1(_09242_),
    .A2(_04396_),
    .ZN(_04397_));
 AOI21_X1 _13499_ (.A(_09251_),
    .B1(_04397_),
    .B2(_09252_),
    .ZN(_04398_));
 INV_X1 _13500_ (.A(_09249_),
    .ZN(_04399_));
 OAI21_X1 _13501_ (.A(_04392_),
    .B1(_04398_),
    .B2(_04399_),
    .ZN(_04400_));
 AOI21_X1 _13502_ (.A(_09257_),
    .B1(_04400_),
    .B2(_09258_),
    .ZN(_04401_));
 OAI21_X1 _13503_ (.A(_04391_),
    .B1(_04401_),
    .B2(_04136_),
    .ZN(_04402_));
 NAND2_X1 _13504_ (.A1(_09261_),
    .A2(_04402_),
    .ZN(_04403_));
 NAND4_X4 _13505_ (.A1(_04231_),
    .A2(_04389_),
    .A3(_04390_),
    .A4(_04403_),
    .ZN(_04404_));
 NOR3_X2 _13506_ (.A1(_04325_),
    .A2(_04330_),
    .A3(_04404_),
    .ZN(_04405_));
 NAND2_X1 _13507_ (.A1(_04388_),
    .A2(_04405_),
    .ZN(_04406_));
 AND4_X1 _13508_ (.A1(_04290_),
    .A2(_04301_),
    .A3(_04331_),
    .A4(_04354_),
    .ZN(_04407_));
 BUF_X4 _13509_ (.A(_04407_),
    .Z(_04408_));
 XNOR2_X2 _13510_ (.A(_04199_),
    .B(_04217_),
    .ZN(_04409_));
 OAI33_X1 _13511_ (.A1(_04230_),
    .A2(_04234_),
    .A3(_04239_),
    .B1(_04243_),
    .B2(_04229_),
    .B3(_04134_),
    .ZN(_04410_));
 NAND2_X2 _13512_ (.A1(_04381_),
    .A2(net374),
    .ZN(_04411_));
 NOR3_X4 _13513_ (.A1(_04380_),
    .A2(_04409_),
    .A3(_04411_),
    .ZN(_04412_));
 AOI21_X2 _13514_ (.A(_04406_),
    .B1(_04408_),
    .B2(_04412_),
    .ZN(_04413_));
 MUX2_X1 _13515_ (.A(_04372_),
    .B(_04375_),
    .S(_04413_),
    .Z(_04414_));
 NOR2_X1 _13516_ (.A1(_04371_),
    .A2(_04370_),
    .ZN(_04415_));
 NAND3_X1 _13517_ (.A1(_04283_),
    .A2(_04284_),
    .A3(_04362_),
    .ZN(_04416_));
 INV_X1 _13518_ (.A(_04416_),
    .ZN(_04417_));
 AOI21_X1 _13519_ (.A(_04363_),
    .B1(_04361_),
    .B2(_04360_),
    .ZN(_04418_));
 AND2_X1 _13520_ (.A1(_04388_),
    .A2(_04405_),
    .ZN(_04419_));
 OAI21_X1 _13521_ (.A(_04419_),
    .B1(_04355_),
    .B2(net406),
    .ZN(_04420_));
 AOI22_X2 _13522_ (.A1(_04415_),
    .A2(_04417_),
    .B1(_04418_),
    .B2(_04420_),
    .ZN(_04421_));
 NAND2_X1 _13523_ (.A1(_04360_),
    .A2(_04361_),
    .ZN(_04422_));
 OR3_X1 _13524_ (.A1(_04283_),
    .A2(_04284_),
    .A3(_04281_),
    .ZN(_04423_));
 OR3_X1 _13525_ (.A1(_04422_),
    .A2(_04362_),
    .A3(_04423_),
    .ZN(_04424_));
 NOR2_X1 _13526_ (.A1(_04373_),
    .A2(_04423_),
    .ZN(_04425_));
 OAI21_X1 _13527_ (.A(_04425_),
    .B1(_04370_),
    .B2(_04371_),
    .ZN(_04426_));
 AND3_X1 _13528_ (.A1(_04288_),
    .A2(_04274_),
    .A3(_04281_),
    .ZN(_04427_));
 OAI21_X1 _13529_ (.A(_04427_),
    .B1(_04370_),
    .B2(_04371_),
    .ZN(_04428_));
 MUX2_X1 _13530_ (.A(_04426_),
    .B(_04428_),
    .S(_04413_),
    .Z(_04429_));
 NAND4_X4 _13531_ (.A1(_04414_),
    .A2(_04421_),
    .A3(_04424_),
    .A4(_04429_),
    .ZN(_04430_));
 XNOR2_X1 _13532_ (.A(_04232_),
    .B(_04402_),
    .ZN(_04431_));
 NAND2_X2 _13533_ (.A1(_04389_),
    .A2(_04390_),
    .ZN(_04432_));
 XNOR2_X1 _13534_ (.A(_04234_),
    .B(_04432_),
    .ZN(_04433_));
 XNOR2_X1 _13535_ (.A(_04387_),
    .B(_04404_),
    .ZN(_04434_));
 AND2_X2 _13536_ (.A1(_04385_),
    .A2(_04386_),
    .ZN(_04435_));
 NOR3_X1 _13537_ (.A1(_09227_),
    .A2(_09230_),
    .A3(net40),
    .ZN(_04436_));
 NOR3_X1 _13538_ (.A1(_04245_),
    .A2(_04020_),
    .A3(_04239_),
    .ZN(_04437_));
 OAI21_X1 _13539_ (.A(_04435_),
    .B1(_04436_),
    .B2(_04437_),
    .ZN(_04438_));
 OAI33_X1 _13540_ (.A1(_04431_),
    .A2(_04433_),
    .A3(_04434_),
    .B1(_04438_),
    .B2(_04248_),
    .B3(_04355_),
    .ZN(_04439_));
 CLKBUF_X3 _13541_ (.A(_09281_),
    .Z(_04440_));
 INV_X1 _13542_ (.A(_09283_),
    .ZN(_04441_));
 INV_X1 _13543_ (.A(_09271_),
    .ZN(_04442_));
 INV_X1 _13544_ (.A(_09277_),
    .ZN(_04443_));
 INV_X1 _13545_ (.A(_09265_),
    .ZN(_04444_));
 OAI21_X1 _13546_ (.A(_09266_),
    .B1(_09285_),
    .B2(\butterfly_count[1] ),
    .ZN(_04445_));
 NAND2_X1 _13547_ (.A1(_04444_),
    .A2(_04445_),
    .ZN(_04446_));
 NAND2_X2 clone5 (.A1(_03788_),
    .A2(_03749_),
    .ZN(net5));
 AOI21_X1 _13549_ (.A(_09263_),
    .B1(_04446_),
    .B2(_09264_),
    .ZN(_04448_));
 INV_X1 _13550_ (.A(_09278_),
    .ZN(_04449_));
 OAI21_X1 _13551_ (.A(_04443_),
    .B1(_04448_),
    .B2(_04449_),
    .ZN(_04450_));
 AOI21_X1 _13552_ (.A(_09274_),
    .B1(_04450_),
    .B2(_09275_),
    .ZN(_04451_));
 INV_X1 _13553_ (.A(_09272_),
    .ZN(_04452_));
 OAI21_X2 _13554_ (.A(_04442_),
    .B1(_04451_),
    .B2(_04452_),
    .ZN(_04453_));
 AOI21_X2 _13555_ (.A(_09268_),
    .B1(_04453_),
    .B2(_09269_),
    .ZN(_04454_));
 INV_X2 _13556_ (.A(_09284_),
    .ZN(_04455_));
 OAI21_X4 _13557_ (.A(_04441_),
    .B1(_04454_),
    .B2(_04455_),
    .ZN(_04456_));
 AOI21_X4 _13558_ (.A(_09280_),
    .B1(_04440_),
    .B2(_04456_),
    .ZN(_04457_));
 NAND2_X4 _13559_ (.A1(net373),
    .A2(_04457_),
    .ZN(_04458_));
 NAND2_X1 _13560_ (.A1(_04327_),
    .A2(_04328_),
    .ZN(_04459_));
 OAI21_X2 _13561_ (.A(_04329_),
    .B1(_04459_),
    .B2(_04245_),
    .ZN(_04460_));
 OR4_X1 _13562_ (.A1(_04248_),
    .A2(_04315_),
    .A3(_04325_),
    .A4(_04408_),
    .ZN(_04461_));
 XOR2_X2 _13563_ (.A(_04460_),
    .B(_04461_),
    .Z(_04462_));
 AND2_X1 _13564_ (.A1(_04281_),
    .A2(_04326_),
    .ZN(_04463_));
 NOR3_X1 _13565_ (.A1(_04325_),
    .A2(_04404_),
    .A3(_04460_),
    .ZN(_04464_));
 NAND2_X1 _13566_ (.A1(_04388_),
    .A2(_04464_),
    .ZN(_04465_));
 AOI21_X4 _13567_ (.A(_04465_),
    .B1(_04408_),
    .B2(_04412_),
    .ZN(_04466_));
 XOR2_X2 _13568_ (.A(_04463_),
    .B(_04466_),
    .Z(_04467_));
 NOR3_X2 _13569_ (.A1(_04380_),
    .A2(_04384_),
    .A3(_04387_),
    .ZN(_04468_));
 NOR2_X2 _13570_ (.A1(_04387_),
    .A2(_04404_),
    .ZN(_04469_));
 NAND2_X1 _13571_ (.A1(_04181_),
    .A2(_04134_),
    .ZN(_04470_));
 AOI21_X1 _13572_ (.A(_04202_),
    .B1(_04082_),
    .B2(net14),
    .ZN(_04471_));
 NOR2_X1 _13573_ (.A1(_04225_),
    .A2(_04471_),
    .ZN(_04472_));
 XNOR2_X2 _13574_ (.A(_04470_),
    .B(_04472_),
    .ZN(_04473_));
 AOI21_X2 _13575_ (.A(_04205_),
    .B1(_04220_),
    .B2(_04188_),
    .ZN(_04474_));
 AND3_X1 _13576_ (.A1(_04188_),
    .A2(_04205_),
    .A3(_04220_),
    .ZN(_04475_));
 OR2_X1 _13577_ (.A1(_04474_),
    .A2(_04475_),
    .ZN(_04476_));
 NAND4_X1 _13578_ (.A1(_04246_),
    .A2(_04469_),
    .A3(_04473_),
    .A4(_04476_),
    .ZN(_04477_));
 OAI21_X1 _13579_ (.A(_04199_),
    .B1(_04206_),
    .B2(_04095_),
    .ZN(_04478_));
 AOI21_X2 _13580_ (.A(_04228_),
    .B1(_04478_),
    .B2(net40),
    .ZN(_04479_));
 NAND4_X1 _13581_ (.A1(_04197_),
    .A2(net374),
    .A3(_04479_),
    .A4(_04435_),
    .ZN(_04480_));
 OR3_X1 _13582_ (.A1(_04410_),
    .A2(_04387_),
    .A3(_04404_),
    .ZN(_04481_));
 OAI21_X2 _13583_ (.A(net374),
    .B1(_04474_),
    .B2(_04475_),
    .ZN(_04482_));
 OR3_X2 _13584_ (.A1(_04410_),
    .A2(_04474_),
    .A3(_04475_),
    .ZN(_04483_));
 NAND4_X1 _13585_ (.A1(_04480_),
    .A2(_04481_),
    .A3(_04482_),
    .A4(_04483_),
    .ZN(_04484_));
 OAI222_X2 _13586_ (.A1(net405),
    .A2(_04355_),
    .B1(_04468_),
    .B2(_04477_),
    .C1(_04484_),
    .C2(_04473_),
    .ZN(_04485_));
 XNOR2_X2 _13587_ (.A(_04218_),
    .B(_04247_),
    .ZN(_04486_));
 AOI21_X4 _13588_ (.A(_04197_),
    .B1(_04479_),
    .B2(_04469_),
    .ZN(_04487_));
 OAI21_X2 _13589_ (.A(_04197_),
    .B1(_04218_),
    .B2(_04247_),
    .ZN(_04488_));
 OAI22_X4 _13590_ (.A1(_04486_),
    .A2(_04487_),
    .B1(_04488_),
    .B2(_04355_),
    .ZN(_04489_));
 NAND2_X2 _13591_ (.A1(_04134_),
    .A2(_04309_),
    .ZN(_04490_));
 MUX2_X2 _13592_ (.A(_04309_),
    .B(_04490_),
    .S(_04313_),
    .Z(_04491_));
 NOR3_X2 _13593_ (.A1(_04248_),
    .A2(_04408_),
    .A3(_04491_),
    .ZN(_04492_));
 INV_X1 _13594_ (.A(_04491_),
    .ZN(_04493_));
 AOI21_X2 _13595_ (.A(_04493_),
    .B1(_04355_),
    .B2(_04412_),
    .ZN(_04494_));
 OAI211_X4 _13596_ (.A(_04485_),
    .B(_04489_),
    .C1(_04492_),
    .C2(_04494_),
    .ZN(_04495_));
 NOR2_X1 _13597_ (.A1(_04379_),
    .A2(_04310_),
    .ZN(_04496_));
 OAI22_X4 _13598_ (.A1(_04312_),
    .A2(_04490_),
    .B1(_04496_),
    .B2(_04304_),
    .ZN(_04497_));
 NAND2_X1 _13599_ (.A1(_04231_),
    .A2(_04403_),
    .ZN(_04498_));
 NOR2_X2 _13600_ (.A1(_04432_),
    .A2(_04498_),
    .ZN(_04499_));
 AND3_X1 _13601_ (.A1(_04499_),
    .A2(_04468_),
    .A3(_04491_),
    .ZN(_04500_));
 OAI21_X2 _13602_ (.A(_04500_),
    .B1(_04355_),
    .B2(_04248_),
    .ZN(_04501_));
 XNOR2_X2 _13603_ (.A(_04497_),
    .B(_04501_),
    .ZN(_04502_));
 AOI21_X2 _13604_ (.A(_04322_),
    .B1(_04316_),
    .B2(net40),
    .ZN(_04503_));
 NOR4_X1 _13605_ (.A1(_04380_),
    .A2(_04409_),
    .A3(_04411_),
    .A4(_04315_),
    .ZN(_04504_));
 OR2_X1 _13606_ (.A1(_04503_),
    .A2(_04504_),
    .ZN(_04505_));
 NAND2_X1 _13607_ (.A1(_04503_),
    .A2(_04504_),
    .ZN(_04506_));
 OAI21_X4 _13608_ (.A(_04505_),
    .B1(_04506_),
    .B2(net399),
    .ZN(_04507_));
 NAND2_X1 _13609_ (.A1(_04253_),
    .A2(_04323_),
    .ZN(_04508_));
 AND2_X1 _13610_ (.A1(_04320_),
    .A2(_04508_),
    .ZN(_04509_));
 NAND3_X2 _13611_ (.A1(_04503_),
    .A2(_04388_),
    .A3(_04499_),
    .ZN(_04510_));
 AOI21_X4 _13612_ (.A(_04510_),
    .B1(_04408_),
    .B2(_04412_),
    .ZN(_04511_));
 XNOR2_X2 _13613_ (.A(_04509_),
    .B(_04511_),
    .ZN(_04512_));
 NOR4_X4 _13614_ (.A1(_04495_),
    .A2(_04502_),
    .A3(_04507_),
    .A4(_04512_),
    .ZN(_04513_));
 NAND3_X1 _13615_ (.A1(_04462_),
    .A2(_04467_),
    .A3(_04513_),
    .ZN(_04514_));
 NOR3_X4 _13616_ (.A1(_04495_),
    .A2(_04502_),
    .A3(_04507_),
    .ZN(_04515_));
 XOR2_X2 _13617_ (.A(_04509_),
    .B(_04511_),
    .Z(_04516_));
 AND2_X2 _13618_ (.A1(_04462_),
    .A2(_04516_),
    .ZN(_04517_));
 XNOR2_X2 _13619_ (.A(_04463_),
    .B(_04466_),
    .ZN(_04518_));
 NOR2_X2 _13620_ (.A1(_04368_),
    .A2(_04518_),
    .ZN(_04519_));
 AND4_X4 _13621_ (.A1(_04430_),
    .A2(_04515_),
    .A3(_04517_),
    .A4(_04519_),
    .ZN(_04520_));
 BUF_X8 _13622_ (.A(_04520_),
    .Z(_04521_));
 XOR2_X2 _13623_ (.A(_04297_),
    .B(_04299_),
    .Z(_04522_));
 AOI21_X2 _13624_ (.A(_04432_),
    .B1(_04408_),
    .B2(_04412_),
    .ZN(_04523_));
 AND3_X1 _13625_ (.A1(_04290_),
    .A2(_04331_),
    .A3(_04468_),
    .ZN(_04524_));
 OAI21_X1 _13626_ (.A(_04498_),
    .B1(_04491_),
    .B2(_09260_),
    .ZN(_04525_));
 NAND3_X2 _13627_ (.A1(_04523_),
    .A2(_04524_),
    .A3(_04525_),
    .ZN(_04526_));
 XNOR2_X2 _13628_ (.A(_04522_),
    .B(_04526_),
    .ZN(_04527_));
 AOI21_X2 _13629_ (.A(_04351_),
    .B1(_04121_),
    .B2(_04291_),
    .ZN(_04528_));
 XNOR2_X2 _13630_ (.A(_04335_),
    .B(_04528_),
    .ZN(_04529_));
 NOR2_X1 _13631_ (.A1(_04325_),
    .A2(_04330_),
    .ZN(_04530_));
 NAND4_X1 _13632_ (.A1(_04290_),
    .A2(_04301_),
    .A3(_04530_),
    .A4(_04388_),
    .ZN(_04531_));
 AOI211_X2 _13633_ (.A(_04404_),
    .B(_04531_),
    .C1(_04412_),
    .C2(_04408_),
    .ZN(_04532_));
 XNOR2_X2 _13634_ (.A(_04529_),
    .B(_04532_),
    .ZN(_04533_));
 AND4_X1 _13635_ (.A1(_04290_),
    .A2(_04522_),
    .A3(_04360_),
    .A4(_04361_),
    .ZN(_04534_));
 XOR2_X2 _13636_ (.A(_04296_),
    .B(_04534_),
    .Z(_04535_));
 XOR2_X1 _13637_ (.A(_04335_),
    .B(_04528_),
    .Z(_04536_));
 NOR4_X1 _13638_ (.A1(_04296_),
    .A2(_04300_),
    .A3(_04353_),
    .A4(_04536_),
    .ZN(_04537_));
 NAND4_X1 _13639_ (.A1(_04290_),
    .A2(_04388_),
    .A3(_04405_),
    .A4(_04537_),
    .ZN(_04538_));
 AOI21_X1 _13640_ (.A(_04538_),
    .B1(_04408_),
    .B2(_04412_),
    .ZN(_04539_));
 NAND2_X1 _13641_ (.A1(_03880_),
    .A2(_04340_),
    .ZN(_04540_));
 OAI221_X2 _13642_ (.A(_03873_),
    .B1(_03878_),
    .B2(_03879_),
    .C1(_03875_),
    .C2(_03788_),
    .ZN(_04541_));
 OAI21_X1 _13643_ (.A(_04540_),
    .B1(_04541_),
    .B2(_04340_),
    .ZN(_04542_));
 OAI21_X1 _13644_ (.A(_03867_),
    .B1(_03881_),
    .B2(_04103_),
    .ZN(_04543_));
 OR2_X1 _13645_ (.A1(_03867_),
    .A2(_04103_),
    .ZN(_04544_));
 AND4_X1 _13646_ (.A1(_04124_),
    .A2(_04338_),
    .A3(_04543_),
    .A4(_04544_),
    .ZN(_04545_));
 XNOR2_X2 _13647_ (.A(_04542_),
    .B(_04545_),
    .ZN(_04546_));
 XNOR2_X2 _13648_ (.A(_04539_),
    .B(_04546_),
    .ZN(_04547_));
 NOR4_X4 _13649_ (.A1(_04353_),
    .A2(_04533_),
    .A3(_04535_),
    .A4(_04547_),
    .ZN(_04548_));
 AND2_X1 _13650_ (.A1(_04290_),
    .A2(_04301_),
    .ZN(_04549_));
 NAND3_X1 _13651_ (.A1(_04549_),
    .A2(_04331_),
    .A3(_04359_),
    .ZN(_04550_));
 OAI21_X2 _13652_ (.A(_04348_),
    .B1(_04550_),
    .B2(net406),
    .ZN(_04551_));
 INV_X1 _13653_ (.A(_09268_),
    .ZN(_04552_));
 INV_X1 _13654_ (.A(_09274_),
    .ZN(_04553_));
 INV_X1 _13655_ (.A(_09263_),
    .ZN(_04554_));
 OAI21_X2 _13656_ (.A(_09264_),
    .B1(_09266_),
    .B2(_09265_),
    .ZN(_04555_));
 NAND2_X2 _13657_ (.A1(_04555_),
    .A2(_04554_),
    .ZN(_04556_));
 AOI21_X2 _13658_ (.A(_09277_),
    .B1(_04556_),
    .B2(_09278_),
    .ZN(_04557_));
 INV_X1 _13659_ (.A(_09275_),
    .ZN(_04558_));
 OAI21_X4 _13660_ (.A(_04553_),
    .B1(_04558_),
    .B2(_04557_),
    .ZN(_04559_));
 AOI21_X4 _13661_ (.A(_09271_),
    .B1(_09272_),
    .B2(_04559_),
    .ZN(_04560_));
 INV_X1 _13662_ (.A(_09269_),
    .ZN(_04561_));
 OAI21_X4 _13663_ (.A(_04552_),
    .B1(_04560_),
    .B2(_04561_),
    .ZN(_04562_));
 AOI21_X4 _13664_ (.A(_09283_),
    .B1(_04562_),
    .B2(_09284_),
    .ZN(_04563_));
 INV_X2 _13665_ (.A(_04563_),
    .ZN(_04564_));
 AOI21_X4 _13666_ (.A(_09280_),
    .B1(_04440_),
    .B2(_04564_),
    .ZN(_04565_));
 AND3_X4 _13667_ (.A1(_04565_),
    .A2(_04551_),
    .A3(net373),
    .ZN(_04566_));
 AND3_X4 _13668_ (.A1(_04527_),
    .A2(_04548_),
    .A3(_04566_),
    .ZN(_04567_));
 BUF_X8 _13669_ (.A(_04567_),
    .Z(_04568_));
 AOI211_X2 _13670_ (.A(_04458_),
    .B(_04514_),
    .C1(_04521_),
    .C2(net34),
    .ZN(_04569_));
 NAND2_X1 _13671_ (.A1(_04430_),
    .A2(_04569_),
    .ZN(_04570_));
 XNOR2_X2 _13672_ (.A(_04368_),
    .B(_04570_),
    .ZN(_04571_));
 NAND2_X1 _13673_ (.A1(_04462_),
    .A2(_04513_),
    .ZN(_04572_));
 NAND2_X4 _13674_ (.A1(_04439_),
    .A2(_04565_),
    .ZN(_04573_));
 AOI211_X2 _13675_ (.A(_04572_),
    .B(_04573_),
    .C1(_04521_),
    .C2(_04568_),
    .ZN(_04574_));
 XNOR2_X2 _13676_ (.A(_04518_),
    .B(_04574_),
    .ZN(_04575_));
 INV_X1 _13677_ (.A(_04495_),
    .ZN(_04576_));
 XOR2_X2 _13678_ (.A(_04497_),
    .B(_04501_),
    .Z(_04577_));
 NOR3_X1 _13679_ (.A1(_04577_),
    .A2(_04507_),
    .A3(_04573_),
    .ZN(_04578_));
 NAND3_X4 _13680_ (.A1(_04527_),
    .A2(_04548_),
    .A3(net413),
    .ZN(_04579_));
 NAND4_X4 _13681_ (.A1(_04430_),
    .A2(_04515_),
    .A3(_04517_),
    .A4(_04519_),
    .ZN(_04580_));
 OAI211_X2 _13682_ (.A(_04576_),
    .B(_04578_),
    .C1(_04579_),
    .C2(_04580_),
    .ZN(_04581_));
 AND2_X1 _13683_ (.A1(net373),
    .A2(_04457_),
    .ZN(_04582_));
 NOR2_X1 _13684_ (.A1(_04507_),
    .A2(_04582_),
    .ZN(_04583_));
 AND2_X1 _13685_ (.A1(_04507_),
    .A2(_04582_),
    .ZN(_04584_));
 AOI21_X1 _13686_ (.A(_04583_),
    .B1(_04584_),
    .B2(_04576_),
    .ZN(_04585_));
 NAND2_X1 _13687_ (.A1(_04577_),
    .A2(_04573_),
    .ZN(_04586_));
 AOI21_X1 _13688_ (.A(_04495_),
    .B1(_04521_),
    .B2(net34),
    .ZN(_04587_));
 OR2_X1 _13689_ (.A1(_04502_),
    .A2(_04507_),
    .ZN(_04588_));
 OAI221_X2 _13690_ (.A(_04581_),
    .B1(_04585_),
    .B2(_04586_),
    .C1(_04587_),
    .C2(_04588_),
    .ZN(_04589_));
 INV_X1 _13691_ (.A(_04573_),
    .ZN(_04590_));
 AND3_X1 _13692_ (.A1(_04462_),
    .A2(_04512_),
    .A3(_04590_),
    .ZN(_04591_));
 OAI21_X2 _13693_ (.A(_04515_),
    .B1(_04580_),
    .B2(_04579_),
    .ZN(_04592_));
 MUX2_X2 _13694_ (.A(_04591_),
    .B(_04517_),
    .S(_04592_),
    .Z(_04593_));
 NAND3_X1 _13695_ (.A1(_04517_),
    .A2(_04458_),
    .A3(_04573_),
    .ZN(_04594_));
 OR4_X1 _13696_ (.A1(_04462_),
    .A2(_04512_),
    .A3(_04458_),
    .A4(_04590_),
    .ZN(_04595_));
 OAI21_X2 _13697_ (.A(_04594_),
    .B1(_04595_),
    .B2(_04592_),
    .ZN(_04596_));
 OAI211_X4 _13698_ (.A(_04575_),
    .B(_04589_),
    .C1(_04593_),
    .C2(_04596_),
    .ZN(_04597_));
 NAND2_X1 _13699_ (.A1(_04413_),
    .A2(_04362_),
    .ZN(_04598_));
 XNOR2_X1 _13700_ (.A(_04281_),
    .B(_04598_),
    .ZN(_04599_));
 NAND2_X1 _13701_ (.A1(_04274_),
    .A2(_04599_),
    .ZN(_04600_));
 AOI21_X1 _13702_ (.A(_04274_),
    .B1(_04413_),
    .B2(_04373_),
    .ZN(_04601_));
 OAI221_X2 _13703_ (.A(_04600_),
    .B1(_04601_),
    .B2(_04288_),
    .C1(_04263_),
    .C2(_04599_),
    .ZN(_04602_));
 XNOR2_X1 _13704_ (.A(_04283_),
    .B(_04362_),
    .ZN(_04603_));
 XNOR2_X2 _13705_ (.A(_04422_),
    .B(_04603_),
    .ZN(_04604_));
 INV_X1 _13706_ (.A(_04604_),
    .ZN(_04605_));
 NAND4_X1 _13707_ (.A1(_04462_),
    .A2(_04467_),
    .A3(_04513_),
    .A4(_04605_),
    .ZN(_04606_));
 AOI211_X2 _13708_ (.A(_04573_),
    .B(_04606_),
    .C1(_04521_),
    .C2(net34),
    .ZN(_04607_));
 XNOR2_X2 _13709_ (.A(_04602_),
    .B(_04607_),
    .ZN(_04608_));
 XNOR2_X2 _13710_ (.A(_04569_),
    .B(_04604_),
    .ZN(_04609_));
 NAND2_X1 _13711_ (.A1(_04608_),
    .A2(_04609_),
    .ZN(_04610_));
 NOR3_X4 _13712_ (.A1(_04571_),
    .A2(_04597_),
    .A3(_04610_),
    .ZN(_04611_));
 XNOR2_X1 _13713_ (.A(_04146_),
    .B(_04400_),
    .ZN(_04612_));
 XNOR2_X1 _13714_ (.A(_02757_),
    .B(_02796_),
    .ZN(_04613_));
 OR4_X1 _13715_ (.A1(_02103_),
    .A2(_03003_),
    .A3(_04613_),
    .A4(_03100_),
    .ZN(_04614_));
 NAND2_X1 _13716_ (.A1(_03048_),
    .A2(_04614_),
    .ZN(_04615_));
 AOI21_X1 _13717_ (.A(_02103_),
    .B1(_02796_),
    .B2(_03100_),
    .ZN(_04616_));
 OAI21_X1 _13718_ (.A(_02757_),
    .B1(_02796_),
    .B2(_03100_),
    .ZN(_04617_));
 NAND2_X1 _13719_ (.A1(_04616_),
    .A2(_04617_),
    .ZN(_04618_));
 AOI21_X2 _13720_ (.A(_04615_),
    .B1(_04618_),
    .B2(_03003_),
    .ZN(_04619_));
 NAND3_X4 _13721_ (.A1(_03773_),
    .A2(_04619_),
    .A3(_03552_),
    .ZN(_04620_));
 XOR2_X2 _13722_ (.A(_03049_),
    .B(_04614_),
    .Z(_04621_));
 XOR2_X2 _13723_ (.A(_04621_),
    .B(_04620_),
    .Z(_09145_));
 NOR2_X2 _13724_ (.A1(_03354_),
    .A2(_09145_),
    .ZN(_04622_));
 AOI21_X2 _13725_ (.A(_04622_),
    .B1(_03354_),
    .B2(_09147_),
    .ZN(_09165_));
 XOR2_X1 _13726_ (.A(_09167_),
    .B(_03996_),
    .Z(_04623_));
 MUX2_X1 _13727_ (.A(_09165_),
    .B(_04623_),
    .S(_03524_),
    .Z(_09183_));
 NAND2_X1 _13728_ (.A1(_03543_),
    .A2(_03554_),
    .ZN(_04624_));
 XNOR2_X1 _13729_ (.A(_03568_),
    .B(_04624_),
    .ZN(_04625_));
 MUX2_X1 _13730_ (.A(_09183_),
    .B(_04625_),
    .S(_03791_),
    .Z(_09212_));
 OR3_X1 _13731_ (.A1(_09214_),
    .A2(_09193_),
    .A3(_03815_),
    .ZN(_04626_));
 AND2_X1 _13732_ (.A1(_03816_),
    .A2(_04626_),
    .ZN(_04627_));
 MUX2_X1 _13733_ (.A(_09212_),
    .B(_04627_),
    .S(_03991_),
    .Z(_09236_));
 XNOR2_X1 _13734_ (.A(_09238_),
    .B(_04015_),
    .ZN(_04628_));
 MUX2_X1 _13735_ (.A(_09236_),
    .B(_04628_),
    .S(_04135_),
    .Z(_09256_));
 MUX2_X1 _13736_ (.A(_04612_),
    .B(_09256_),
    .S(net26),
    .Z(_09282_));
 OR3_X2 _13737_ (.A1(_04580_),
    .A2(_04579_),
    .A3(_09282_),
    .ZN(_04629_));
 XNOR2_X1 _13738_ (.A(_04455_),
    .B(_04562_),
    .ZN(_04630_));
 INV_X1 _13739_ (.A(_04630_),
    .ZN(_04631_));
 OAI21_X4 _13740_ (.A(_04631_),
    .B1(_04579_),
    .B2(_04580_),
    .ZN(_04632_));
 AOI21_X4 _13741_ (.A(_08819_),
    .B1(_04629_),
    .B2(_04632_),
    .ZN(_04633_));
 AND3_X2 _13742_ (.A1(_08819_),
    .A2(_04629_),
    .A3(_04632_),
    .ZN(_04634_));
 INV_X1 _13743_ (.A(_09301_),
    .ZN(_04635_));
 INV_X1 _13744_ (.A(_09305_),
    .ZN(_04636_));
 INV_X1 _13745_ (.A(_09307_),
    .ZN(_04637_));
 INV_X1 _13746_ (.A(_09293_),
    .ZN(_04638_));
 INV_X1 _13747_ (.A(_09295_),
    .ZN(_04639_));
 OAI21_X2 _13748_ (.A(_09296_),
    .B1(_09288_),
    .B2(_09289_),
    .ZN(_04640_));
 AOI21_X4 _13749_ (.A(_04638_),
    .B1(_04640_),
    .B2(_04639_),
    .ZN(_04641_));
 OAI21_X4 _13750_ (.A(_09308_),
    .B1(_09292_),
    .B2(_04641_),
    .ZN(_04642_));
 AOI21_X4 _13751_ (.A(_04636_),
    .B1(_04637_),
    .B2(_04642_),
    .ZN(_04643_));
 OAI21_X4 _13752_ (.A(_09302_),
    .B1(_04643_),
    .B2(_09304_),
    .ZN(_04644_));
 NAND2_X4 _13753_ (.A1(_04635_),
    .A2(_04644_),
    .ZN(_04645_));
 BUF_X2 _13754_ (.A(_09299_),
    .Z(_04646_));
 AOI21_X4 _13755_ (.A(_09298_),
    .B1(_04645_),
    .B2(_04646_),
    .ZN(_04647_));
 NOR3_X4 _13756_ (.A1(_04647_),
    .A2(_04633_),
    .A3(_04634_),
    .ZN(_04648_));
 NOR2_X2 _13757_ (.A1(net26),
    .A2(_04404_),
    .ZN(_04649_));
 OR2_X1 _13758_ (.A1(_04431_),
    .A2(_04433_),
    .ZN(_04650_));
 INV_X1 _13759_ (.A(_04565_),
    .ZN(_04651_));
 AOI211_X2 _13760_ (.A(_04650_),
    .B(_04651_),
    .C1(net410),
    .C2(_04520_),
    .ZN(_04652_));
 OAI21_X2 _13761_ (.A(_04435_),
    .B1(_04649_),
    .B2(_04652_),
    .ZN(_04653_));
 OR3_X2 _13762_ (.A1(_04435_),
    .A2(_04649_),
    .A3(_04652_),
    .ZN(_04654_));
 NAND3_X2 _13763_ (.A1(_02573_),
    .A2(_04629_),
    .A3(_04632_),
    .ZN(_04655_));
 INV_X1 _13764_ (.A(_04457_),
    .ZN(_04656_));
 NAND3_X1 _13765_ (.A1(_04234_),
    .A2(_04389_),
    .A3(_04390_),
    .ZN(_04657_));
 OAI21_X1 _13766_ (.A(_04657_),
    .B1(_04523_),
    .B2(_04234_),
    .ZN(_04658_));
 MUX2_X2 _13767_ (.A(_04431_),
    .B(_09259_),
    .S(_04356_),
    .Z(_04659_));
 OR4_X1 _13768_ (.A1(net412),
    .A2(_04656_),
    .A3(_04658_),
    .A4(_04659_),
    .ZN(_04660_));
 AND2_X1 _13769_ (.A1(_04651_),
    .A2(_04659_),
    .ZN(_04661_));
 OAI21_X1 _13770_ (.A(_04658_),
    .B1(_04659_),
    .B2(_04656_),
    .ZN(_04662_));
 OAI21_X1 _13771_ (.A(_04660_),
    .B1(_04661_),
    .B2(_04662_),
    .ZN(_04663_));
 XNOR2_X2 _13772_ (.A(_04440_),
    .B(_04456_),
    .ZN(_04664_));
 OAI211_X2 _13773_ (.A(_04663_),
    .B(_04664_),
    .C1(_04580_),
    .C2(_04579_),
    .ZN(_04665_));
 NAND2_X4 _13774_ (.A1(_04568_),
    .A2(_04521_),
    .ZN(_04666_));
 OAI21_X2 _13775_ (.A(_04665_),
    .B1(net37),
    .B2(_09279_),
    .ZN(_04667_));
 NAND4_X4 _13776_ (.A1(_04653_),
    .A2(_04654_),
    .A3(_04655_),
    .A4(_04667_),
    .ZN(_04668_));
 NOR2_X1 _13777_ (.A1(_04494_),
    .A2(_04492_),
    .ZN(_04669_));
 NAND2_X1 _13778_ (.A1(_04485_),
    .A2(_04489_),
    .ZN(_04670_));
 AOI211_X2 _13779_ (.A(_04458_),
    .B(_04670_),
    .C1(_04521_),
    .C2(_04568_),
    .ZN(_04671_));
 XNOR2_X2 _13780_ (.A(_04669_),
    .B(_04671_),
    .ZN(_04672_));
 NAND2_X1 _13781_ (.A1(_04409_),
    .A2(_04411_),
    .ZN(_04673_));
 NAND2_X1 _13782_ (.A1(_04218_),
    .A2(_04247_),
    .ZN(_04674_));
 OAI21_X2 _13783_ (.A(_04673_),
    .B1(net401),
    .B2(_04674_),
    .ZN(_04675_));
 XNOR2_X1 _13784_ (.A(_04469_),
    .B(_04473_),
    .ZN(_04676_));
 AND2_X1 _13785_ (.A1(_04246_),
    .A2(_04476_),
    .ZN(_04677_));
 NOR2_X1 _13786_ (.A1(_04473_),
    .A2(_04476_),
    .ZN(_04678_));
 AOI221_X2 _13787_ (.A(net400),
    .B1(_04676_),
    .B2(_04677_),
    .C1(_04678_),
    .C2(_04410_),
    .ZN(_04679_));
 OR2_X1 _13788_ (.A1(_04675_),
    .A2(_04679_),
    .ZN(_04680_));
 AOI211_X2 _13789_ (.A(_04573_),
    .B(_04680_),
    .C1(_04520_),
    .C2(_04568_),
    .ZN(_04681_));
 NAND2_X1 _13790_ (.A1(_04435_),
    .A2(_04499_),
    .ZN(_04682_));
 NOR4_X2 _13791_ (.A1(_04380_),
    .A2(net26),
    .A3(_04384_),
    .A4(_04682_),
    .ZN(_04683_));
 NOR2_X2 _13792_ (.A1(_04487_),
    .A2(_04683_),
    .ZN(_04684_));
 XOR2_X2 _13793_ (.A(_04681_),
    .B(_04684_),
    .Z(_04685_));
 AOI21_X4 _13794_ (.A(_04458_),
    .B1(net423),
    .B2(_04520_),
    .ZN(_04686_));
 OAI21_X4 _13795_ (.A(_04483_),
    .B1(_04482_),
    .B2(net26),
    .ZN(_04687_));
 XNOR2_X2 _13796_ (.A(_04686_),
    .B(_04687_),
    .ZN(_04688_));
 NAND3_X1 _13797_ (.A1(_04435_),
    .A2(_04476_),
    .A3(_04649_),
    .ZN(_04689_));
 XOR2_X2 _13798_ (.A(_04473_),
    .B(_04689_),
    .Z(_04690_));
 INV_X1 _13799_ (.A(_04690_),
    .ZN(_04691_));
 NOR2_X2 _13800_ (.A1(_04675_),
    .A2(_04691_),
    .ZN(_04692_));
 NAND4_X4 _13801_ (.A1(_04672_),
    .A2(_04685_),
    .A3(_04688_),
    .A4(_04692_),
    .ZN(_04693_));
 NOR3_X4 _13802_ (.A1(_04648_),
    .A2(_04668_),
    .A3(_04693_),
    .ZN(_04694_));
 XNOR2_X2 _13803_ (.A(_04300_),
    .B(_04526_),
    .ZN(_04695_));
 NOR4_X4 _13804_ (.A1(_04580_),
    .A2(_04695_),
    .A3(net34),
    .A4(_04458_),
    .ZN(_04696_));
 NAND2_X1 _13805_ (.A1(_04548_),
    .A2(_04696_),
    .ZN(_04697_));
 XNOR2_X2 _13806_ (.A(_04551_),
    .B(_04697_),
    .ZN(_04698_));
 NAND2_X1 _13807_ (.A1(_04521_),
    .A2(_04590_),
    .ZN(_04699_));
 NAND4_X1 _13808_ (.A1(net409),
    .A2(_09272_),
    .A3(_09275_),
    .A4(_09278_),
    .ZN(_04700_));
 NAND3_X1 _13809_ (.A1(_09269_),
    .A2(_09266_),
    .A3(_04440_),
    .ZN(_04701_));
 NOR4_X2 _13810_ (.A1(_04455_),
    .A2(_01111_),
    .A3(_04700_),
    .A4(_04701_),
    .ZN(_04702_));
 NAND2_X1 _13811_ (.A1(_04439_),
    .A2(_04702_),
    .ZN(_04703_));
 AND3_X1 _13812_ (.A1(_04548_),
    .A2(_04551_),
    .A3(_04703_),
    .ZN(_04704_));
 OAI21_X2 _13813_ (.A(_04527_),
    .B1(_04699_),
    .B2(_04704_),
    .ZN(_04705_));
 NAND3_X2 _13814_ (.A1(_04521_),
    .A2(_04695_),
    .A3(_04590_),
    .ZN(_04706_));
 AND3_X1 _13815_ (.A1(_04549_),
    .A2(_04415_),
    .A3(_04529_),
    .ZN(_04707_));
 XOR2_X2 _13816_ (.A(_04353_),
    .B(_04707_),
    .Z(_04708_));
 INV_X1 _13817_ (.A(_04708_),
    .ZN(_04709_));
 NAND4_X1 _13818_ (.A1(_04521_),
    .A2(_04527_),
    .A3(_04579_),
    .A4(_04582_),
    .ZN(_04710_));
 OR2_X1 _13819_ (.A1(_04533_),
    .A2(_04535_),
    .ZN(_04711_));
 OAI21_X2 _13820_ (.A(_04709_),
    .B1(_04710_),
    .B2(_04711_),
    .ZN(_04712_));
 OR3_X1 _13821_ (.A1(_04711_),
    .A2(_04710_),
    .A3(_04709_),
    .ZN(_04713_));
 AOI22_X4 _13822_ (.A1(_04705_),
    .A2(_04706_),
    .B1(_04712_),
    .B2(_04713_),
    .ZN(_04714_));
 NOR4_X2 _13823_ (.A1(_04695_),
    .A2(_04535_),
    .A3(_04699_),
    .A4(_04704_),
    .ZN(_04715_));
 XNOR2_X2 _13824_ (.A(_04533_),
    .B(_04715_),
    .ZN(_04716_));
 XNOR2_X2 _13825_ (.A(_04535_),
    .B(_04696_),
    .ZN(_04717_));
 NOR2_X2 _13826_ (.A1(_04580_),
    .A2(_04579_),
    .ZN(_04718_));
 OR4_X1 _13827_ (.A1(_04580_),
    .A2(_04695_),
    .A3(_04711_),
    .A4(_04708_),
    .ZN(_04719_));
 NOR3_X1 _13828_ (.A1(_04718_),
    .A2(_04573_),
    .A3(_04719_),
    .ZN(_04720_));
 XNOR2_X1 _13829_ (.A(_04547_),
    .B(_04720_),
    .ZN(_04721_));
 AND4_X1 _13830_ (.A1(_04714_),
    .A2(_04716_),
    .A3(_04717_),
    .A4(_04721_),
    .ZN(_04722_));
 NAND4_X4 _13831_ (.A1(_04611_),
    .A2(_04694_),
    .A3(_04698_),
    .A4(_04722_),
    .ZN(_04723_));
 BUF_X8 _13832_ (.A(_04723_),
    .Z(_04724_));
 BUF_X8 _13833_ (.A(_04724_),
    .Z(_04725_));
 XNOR2_X1 _13834_ (.A(_04646_),
    .B(_04645_),
    .ZN(_04726_));
 NAND2_X1 _13835_ (.A1(_04725_),
    .A2(_04726_),
    .ZN(_04727_));
 XNOR2_X1 _13836_ (.A(_04399_),
    .B(_04144_),
    .ZN(_04728_));
 NOR2_X1 _13837_ (.A1(_09149_),
    .A2(_03506_),
    .ZN(_09168_));
 NOR2_X1 _13838_ (.A1(_09173_),
    .A2(_09172_),
    .ZN(_04729_));
 XNOR2_X1 _13839_ (.A(_09170_),
    .B(_04729_),
    .ZN(_04730_));
 MUX2_X1 _13840_ (.A(_09168_),
    .B(_04730_),
    .S(_03791_),
    .Z(_09192_));
 XOR2_X1 _13841_ (.A(_09194_),
    .B(_03814_),
    .Z(_04731_));
 MUX2_X1 _13842_ (.A(_09192_),
    .B(_04731_),
    .S(_03991_),
    .Z(_09215_));
 XNOR2_X1 _13843_ (.A(_04014_),
    .B(_04160_),
    .ZN(_04732_));
 MUX2_X1 _13844_ (.A(_09215_),
    .B(_04732_),
    .S(_04135_),
    .Z(_09247_));
 MUX2_X1 _13845_ (.A(_04728_),
    .B(_09247_),
    .S(_04357_),
    .Z(_09267_));
 XNOR2_X1 _13846_ (.A(_04561_),
    .B(_04453_),
    .ZN(_04733_));
 MUX2_X1 _13847_ (.A(_09267_),
    .B(_04733_),
    .S(net37),
    .Z(_09297_));
 OAI21_X1 _13848_ (.A(_04727_),
    .B1(net44),
    .B2(_09297_),
    .ZN(_09310_));
 INV_X1 _13849_ (.A(_09302_),
    .ZN(_04734_));
 INV_X1 _13850_ (.A(_09296_),
    .ZN(_04735_));
 OAI21_X1 _13851_ (.A(_04639_),
    .B1(_09287_),
    .B2(_04735_),
    .ZN(_04736_));
 AOI21_X2 _13852_ (.A(_09292_),
    .B1(_04736_),
    .B2(_09293_),
    .ZN(_04737_));
 INV_X1 _13853_ (.A(_09308_),
    .ZN(_04738_));
 OAI21_X1 _13854_ (.A(_04637_),
    .B1(_04737_),
    .B2(_04738_),
    .ZN(_04739_));
 AOI21_X2 _13855_ (.A(_09304_),
    .B1(_04739_),
    .B2(_09305_),
    .ZN(_04740_));
 XNOR2_X1 _13856_ (.A(_04734_),
    .B(_04740_),
    .ZN(_04741_));
 NAND2_X1 _13857_ (.A1(_04725_),
    .A2(_04741_),
    .ZN(_04742_));
 XNOR2_X1 _13858_ (.A(_04143_),
    .B(_04397_),
    .ZN(_04743_));
 NOR2_X2 _13859_ (.A1(_01929_),
    .A2(_03506_),
    .ZN(_04744_));
 OAI21_X1 _13860_ (.A(_03552_),
    .B1(_03773_),
    .B2(_04744_),
    .ZN(_04745_));
 XOR2_X2 _13861_ (.A(_04619_),
    .B(_04745_),
    .Z(_09171_));
 NOR2_X1 _13862_ (.A1(_01929_),
    .A2(_03553_),
    .ZN(_04746_));
 XNOR2_X1 _13863_ (.A(_09173_),
    .B(_04746_),
    .ZN(_04747_));
 MUX2_X1 _13864_ (.A(_09171_),
    .B(_04747_),
    .S(_03791_),
    .Z(_09195_));
 OR3_X1 _13865_ (.A1(_09199_),
    .A2(_09197_),
    .A3(_09198_),
    .ZN(_04748_));
 AND2_X1 _13866_ (.A1(_03813_),
    .A2(_04748_),
    .ZN(_04749_));
 MUX2_X1 _13867_ (.A(_09195_),
    .B(_04749_),
    .S(_03991_),
    .Z(_09218_));
 XNOR2_X1 _13868_ (.A(_09220_),
    .B(_04011_),
    .ZN(_04750_));
 MUX2_X1 _13869_ (.A(_09218_),
    .B(_04750_),
    .S(_04135_),
    .Z(_09250_));
 MUX2_X1 _13870_ (.A(_04743_),
    .B(_09250_),
    .S(_04357_),
    .Z(_09270_));
 XNOR2_X1 _13871_ (.A(_04452_),
    .B(_04559_),
    .ZN(_04751_));
 MUX2_X1 _13872_ (.A(_09270_),
    .B(_04751_),
    .S(_04666_),
    .Z(_09300_));
 OAI21_X1 _13873_ (.A(_04742_),
    .B1(_09300_),
    .B2(net44),
    .ZN(_09314_));
 AND3_X1 _13874_ (.A1(_04636_),
    .A2(_04637_),
    .A3(_04642_),
    .ZN(_04752_));
 OAI21_X1 _13875_ (.A(_04725_),
    .B1(_04752_),
    .B2(_04643_),
    .ZN(_04753_));
 XOR2_X1 _13876_ (.A(_09243_),
    .B(_04141_),
    .Z(_04754_));
 NOR2_X1 _13877_ (.A1(_09199_),
    .A2(_04165_),
    .ZN(_09221_));
 OR3_X1 _13878_ (.A1(_04008_),
    .A2(_09223_),
    .A3(_09225_),
    .ZN(_04755_));
 AND2_X1 _13879_ (.A1(_04158_),
    .A2(_04755_),
    .ZN(_04756_));
 MUX2_X1 _13880_ (.A(_09221_),
    .B(_04756_),
    .S(_04135_),
    .Z(_09241_));
 MUX2_X1 _13881_ (.A(_04754_),
    .B(_09241_),
    .S(_04357_),
    .Z(_09273_));
 XNOR2_X1 _13882_ (.A(_04558_),
    .B(_04450_),
    .ZN(_04757_));
 MUX2_X1 _13883_ (.A(_09273_),
    .B(_04757_),
    .S(_04666_),
    .Z(_09303_));
 OAI21_X2 _13884_ (.A(_04753_),
    .B1(_09303_),
    .B2(net44),
    .ZN(_09318_));
 XNOR2_X1 _13885_ (.A(_04738_),
    .B(_04737_),
    .ZN(_04758_));
 NAND2_X1 _13886_ (.A1(_04725_),
    .A2(_04758_),
    .ZN(_04759_));
 XNOR2_X1 _13887_ (.A(_09246_),
    .B(_04393_),
    .ZN(_04760_));
 AOI21_X1 _13888_ (.A(_03773_),
    .B1(_03889_),
    .B2(_01150_),
    .ZN(_04761_));
 AOI21_X2 _13889_ (.A(_04761_),
    .B1(_04744_),
    .B2(net23),
    .ZN(_04762_));
 XNOR2_X2 _13890_ (.A(_03552_),
    .B(_04762_),
    .ZN(_09224_));
 XNOR2_X1 _13891_ (.A(_04008_),
    .B(_01710_),
    .ZN(_04763_));
 MUX2_X1 _13892_ (.A(_09224_),
    .B(_04763_),
    .S(_04135_),
    .Z(_09244_));
 MUX2_X1 _13893_ (.A(_04760_),
    .B(_09244_),
    .S(_04357_),
    .Z(_09276_));
 XNOR2_X1 _13894_ (.A(_04449_),
    .B(_04556_),
    .ZN(_04764_));
 MUX2_X1 _13895_ (.A(_09276_),
    .B(_04764_),
    .S(_04666_),
    .Z(_09306_));
 OAI21_X1 _13896_ (.A(_04759_),
    .B1(_09306_),
    .B2(net44),
    .ZN(_09322_));
 AND3_X1 _13897_ (.A1(_04638_),
    .A2(_04639_),
    .A3(_04640_),
    .ZN(_04765_));
 OAI21_X2 _13898_ (.A(_04725_),
    .B1(_04765_),
    .B2(_04641_),
    .ZN(_04766_));
 NOR2_X1 _13899_ (.A1(_09240_),
    .A2(_04357_),
    .ZN(_09262_));
 XOR2_X1 _13900_ (.A(_09264_),
    .B(_04446_),
    .Z(_04767_));
 MUX2_X1 _13901_ (.A(_09262_),
    .B(_04767_),
    .S(_04666_),
    .Z(_09291_));
 OAI21_X2 _13902_ (.A(_04766_),
    .B1(_09291_),
    .B2(net44),
    .ZN(_09326_));
 MUX2_X1 _13903_ (.A(_01095_),
    .B(_09266_),
    .S(_04666_),
    .Z(_04768_));
 INV_X2 _13904_ (.A(_04768_),
    .ZN(_09294_));
 NAND2_X1 _13905_ (.A1(_00860_),
    .A2(net87),
    .ZN(_04769_));
 INV_X1 _13906_ (.A(_09382_),
    .ZN(_04770_));
 INV_X1 _13907_ (.A(net86),
    .ZN(_04771_));
 OAI21_X1 _13908_ (.A(_00853_),
    .B1(_04770_),
    .B2(_04771_),
    .ZN(_04772_));
 AOI21_X1 _13909_ (.A(_00845_),
    .B1(_04769_),
    .B2(_04772_),
    .ZN(_00012_));
 NAND3_X1 _13910_ (.A1(_00848_),
    .A2(_00849_),
    .A3(_00850_),
    .ZN(_04773_));
 AND2_X1 _13911_ (.A1(_09343_),
    .A2(_04773_),
    .ZN(_04774_));
 AND3_X1 _13912_ (.A1(_09374_),
    .A2(\group[0] ),
    .A3(_04774_),
    .ZN(_09348_));
 INV_X2 _13913_ (.A(_00846_),
    .ZN(_04775_));
 NOR2_X4 _13914_ (.A1(_04775_),
    .A2(_01109_),
    .ZN(_04776_));
 AND3_X1 _13915_ (.A1(_00842_),
    .A2(_00851_),
    .A3(_04776_),
    .ZN(_04777_));
 BUF_X4 _13916_ (.A(_04777_),
    .Z(_04778_));
 BUF_X4 _13917_ (.A(_04778_),
    .Z(_04779_));
 MUX2_X1 _13918_ (.A(\idx1[0] ),
    .B(_00042_),
    .S(_04779_),
    .Z(_00013_));
 AND3_X1 _13919_ (.A1(_09374_),
    .A2(\group[1] ),
    .A3(_04774_),
    .ZN(_09350_));
 AND3_X1 _13920_ (.A1(\group[0] ),
    .A2(_09365_),
    .A3(_04774_),
    .ZN(_09353_));
 MUX2_X1 _13921_ (.A(\idx1[1] ),
    .B(_00043_),
    .S(_04779_),
    .Z(_00014_));
 XOR2_X1 _13922_ (.A(_09354_),
    .B(_09356_),
    .Z(_04780_));
 XNOR2_X1 _13923_ (.A(\butterfly_in_group[2] ),
    .B(_09351_),
    .ZN(_04781_));
 XNOR2_X1 _13924_ (.A(_04780_),
    .B(_04781_),
    .ZN(_04782_));
 NAND2_X1 _13925_ (.A1(_09374_),
    .A2(\group[2] ),
    .ZN(_04783_));
 NAND2_X1 _13926_ (.A1(\group[0] ),
    .A2(_09371_),
    .ZN(_04784_));
 NAND2_X1 _13927_ (.A1(\group[1] ),
    .A2(_09365_),
    .ZN(_04785_));
 XOR2_X1 _13928_ (.A(_04784_),
    .B(_04785_),
    .Z(_04786_));
 XNOR2_X1 _13929_ (.A(_04783_),
    .B(_04786_),
    .ZN(_04787_));
 NAND2_X1 _13930_ (.A1(_04774_),
    .A2(_04787_),
    .ZN(_04788_));
 XNOR2_X2 _13931_ (.A(_04782_),
    .B(_04788_),
    .ZN(_04789_));
 MUX2_X1 _13932_ (.A(\idx1[2] ),
    .B(_04789_),
    .S(_04779_),
    .Z(_00015_));
 BUF_X4 _13933_ (.A(\idx2[0] ),
    .Z(_04790_));
 MUX2_X1 _13934_ (.A(_04790_),
    .B(_00044_),
    .S(_04779_),
    .Z(_00016_));
 BUF_X4 _13935_ (.A(\idx2[1] ),
    .Z(_04791_));
 NAND3_X4 _13936_ (.A1(_00842_),
    .A2(_00851_),
    .A3(_04776_),
    .ZN(_04792_));
 NAND2_X1 _13937_ (.A1(_04791_),
    .A2(_04792_),
    .ZN(_04793_));
 OAI21_X1 _13938_ (.A(_04793_),
    .B1(_04792_),
    .B2(_07366_),
    .ZN(_00017_));
 BUF_X4 _13939_ (.A(\idx2[2] ),
    .Z(_04794_));
 XNOR2_X1 _13940_ (.A(_07365_),
    .B(_09329_),
    .ZN(_04795_));
 XNOR2_X1 _13941_ (.A(_04789_),
    .B(_04795_),
    .ZN(_04796_));
 MUX2_X1 _13942_ (.A(_04794_),
    .B(_04796_),
    .S(_04779_),
    .Z(_00018_));
 NAND2_X1 _13943_ (.A1(\twiddle_idx[0] ),
    .A2(_04792_),
    .ZN(_04797_));
 INV_X1 _13944_ (.A(_00849_),
    .ZN(_04798_));
 AND4_X1 _13945_ (.A1(_00848_),
    .A2(_04798_),
    .A3(\butterfly_in_group[2] ),
    .A4(_09362_),
    .ZN(_04799_));
 MUX2_X1 _13946_ (.A(\butterfly_in_group[0] ),
    .B(\butterfly_in_group[1] ),
    .S(_00849_),
    .Z(_04800_));
 NOR2_X2 _13947_ (.A1(_00848_),
    .A2(_09362_),
    .ZN(_04801_));
 AOI21_X4 _13948_ (.A(_04799_),
    .B1(_04800_),
    .B2(_04801_),
    .ZN(_04802_));
 OAI21_X4 _13949_ (.A(_04797_),
    .B1(_04802_),
    .B2(_04792_),
    .ZN(_00006_));
 MUX2_X1 _13950_ (.A(\butterfly_in_group[0] ),
    .B(\butterfly_in_group[2] ),
    .S(_00850_),
    .Z(_04803_));
 NAND2_X1 _13951_ (.A1(_00849_),
    .A2(_04803_),
    .ZN(_04804_));
 NAND3_X1 _13952_ (.A1(_04798_),
    .A2(_00850_),
    .A3(\butterfly_in_group[1] ),
    .ZN(_04805_));
 NAND2_X1 _13953_ (.A1(_04804_),
    .A2(_04805_),
    .ZN(_04806_));
 MUX2_X2 _13954_ (.A(\twiddle_idx[1] ),
    .B(_04806_),
    .S(_04778_),
    .Z(_00019_));
 XNOR2_X1 _13955_ (.A(_00006_),
    .B(_00019_),
    .ZN(_00007_));
 INV_X1 _13956_ (.A(_00019_),
    .ZN(_00008_));
 CLKBUF_X3 _13957_ (.A(_00033_),
    .Z(_04807_));
 CLKBUF_X3 _13958_ (.A(_04807_),
    .Z(_04808_));
 BUF_X4 _13959_ (.A(_00005_),
    .Z(_04809_));
 BUF_X4 _13960_ (.A(_00003_),
    .Z(_04810_));
 BUF_X4 clone52 (.A(_04812_),
    .Z(net52));
 BUF_X16 _13962_ (.A(_00004_),
    .Z(_04812_));
 MUX2_X1 _13963_ (.A(\samples_imag[0][0] ),
    .B(\samples_imag[2][0] ),
    .S(net51),
    .Z(_04813_));
 NOR2_X1 _13964_ (.A1(_04810_),
    .A2(_04813_),
    .ZN(_04814_));
 INV_X2 _13965_ (.A(_00003_),
    .ZN(_04815_));
 MUX2_X1 _13966_ (.A(\samples_imag[1][0] ),
    .B(\samples_imag[3][0] ),
    .S(_00004_),
    .Z(_04816_));
 NOR2_X1 _13967_ (.A1(_04815_),
    .A2(_04816_),
    .ZN(_04817_));
 NOR3_X2 _13968_ (.A1(_04809_),
    .A2(_04814_),
    .A3(_04817_),
    .ZN(_04818_));
 MUX2_X1 _13969_ (.A(\samples_imag[4][0] ),
    .B(\samples_imag[6][0] ),
    .S(net51),
    .Z(_04819_));
 MUX2_X1 _13970_ (.A(\samples_imag[5][0] ),
    .B(\samples_imag[7][0] ),
    .S(net51),
    .Z(_04820_));
 MUX2_X1 _13971_ (.A(_04819_),
    .B(_04820_),
    .S(_04810_),
    .Z(_04821_));
 AOI21_X4 _13972_ (.A(_04818_),
    .B1(_04821_),
    .B2(_04809_),
    .ZN(_04822_));
 OR2_X1 _13973_ (.A1(_04808_),
    .A2(_04822_),
    .ZN(_07701_));
 INV_X2 _13974_ (.A(_07701_),
    .ZN(_09384_));
 BUF_X4 _13975_ (.A(_00032_),
    .Z(_04823_));
 BUF_X4 _13976_ (.A(_04823_),
    .Z(_04824_));
 BUF_X8 _13977_ (.A(_04824_),
    .Z(_04825_));
 BUF_X8 _13978_ (.A(_04812_),
    .Z(_04826_));
 BUF_X8 _13979_ (.A(_04826_),
    .Z(_04827_));
 MUX2_X1 _13980_ (.A(\samples_real[0][13] ),
    .B(\samples_real[2][13] ),
    .S(_04827_),
    .Z(_04828_));
 MUX2_X1 _13981_ (.A(\samples_real[1][13] ),
    .B(\samples_real[3][13] ),
    .S(_04827_),
    .Z(_04829_));
 BUF_X4 _13982_ (.A(_04810_),
    .Z(_04830_));
 MUX2_X1 _13983_ (.A(_04828_),
    .B(_04829_),
    .S(_04830_),
    .Z(_04831_));
 MUX2_X1 _13984_ (.A(\samples_real[4][13] ),
    .B(\samples_real[6][13] ),
    .S(_04827_),
    .Z(_04832_));
 MUX2_X1 _13985_ (.A(\samples_real[5][13] ),
    .B(\samples_real[7][13] ),
    .S(_04827_),
    .Z(_04833_));
 BUF_X4 _13986_ (.A(_04810_),
    .Z(_04834_));
 MUX2_X1 _13987_ (.A(_04832_),
    .B(_04833_),
    .S(_04834_),
    .Z(_04835_));
 BUF_X8 _13988_ (.A(_04809_),
    .Z(_04836_));
 BUF_X8 _13989_ (.A(_04836_),
    .Z(_04837_));
 MUX2_X2 _13990_ (.A(_04831_),
    .B(_04835_),
    .S(_04837_),
    .Z(_04838_));
 INV_X1 _13991_ (.A(_04838_),
    .ZN(_04839_));
 NOR2_X1 _13992_ (.A1(_04825_),
    .A2(_04839_),
    .ZN(_09385_));
 BUF_X16 _13993_ (.A(_04812_),
    .Z(_04840_));
 MUX2_X1 _13994_ (.A(\samples_imag[0][1] ),
    .B(\samples_imag[2][1] ),
    .S(_04840_),
    .Z(_04841_));
 MUX2_X1 _13995_ (.A(\samples_imag[1][1] ),
    .B(\samples_imag[3][1] ),
    .S(_04840_),
    .Z(_04842_));
 MUX2_X1 _13996_ (.A(_04841_),
    .B(_04842_),
    .S(_04830_),
    .Z(_04843_));
 MUX2_X1 _13997_ (.A(\samples_imag[4][1] ),
    .B(\samples_imag[6][1] ),
    .S(_04840_),
    .Z(_04844_));
 MUX2_X1 _13998_ (.A(\samples_imag[5][1] ),
    .B(\samples_imag[7][1] ),
    .S(_04840_),
    .Z(_04845_));
 MUX2_X1 _13999_ (.A(_04844_),
    .B(_04845_),
    .S(_04830_),
    .Z(_04846_));
 BUF_X8 _14000_ (.A(_04836_),
    .Z(_04847_));
 MUX2_X2 _14001_ (.A(_04843_),
    .B(_04846_),
    .S(_04847_),
    .Z(_04848_));
 INV_X2 _14002_ (.A(_04848_),
    .ZN(_04849_));
 NOR2_X4 _14003_ (.A1(_04807_),
    .A2(_04849_),
    .ZN(_07377_));
 CLKBUF_X3 _14004_ (.A(_00035_),
    .Z(_04850_));
 BUF_X4 _14005_ (.A(_04810_),
    .Z(_04851_));
 BUF_X8 _14006_ (.A(_04812_),
    .Z(_04852_));
 MUX2_X1 _14007_ (.A(\samples_imag[0][2] ),
    .B(\samples_imag[2][2] ),
    .S(_04852_),
    .Z(_04853_));
 NOR2_X1 _14008_ (.A1(_04851_),
    .A2(_04853_),
    .ZN(_04854_));
 CLKBUF_X3 _14009_ (.A(_04815_),
    .Z(_04855_));
 MUX2_X1 _14010_ (.A(\samples_imag[1][2] ),
    .B(\samples_imag[3][2] ),
    .S(_04852_),
    .Z(_04856_));
 NOR2_X1 _14011_ (.A1(_04855_),
    .A2(_04856_),
    .ZN(_04857_));
 NOR3_X2 _14012_ (.A1(_04836_),
    .A2(_04854_),
    .A3(_04857_),
    .ZN(_04858_));
 BUF_X4 _14013_ (.A(net51),
    .Z(_04859_));
 MUX2_X1 _14014_ (.A(\samples_imag[4][2] ),
    .B(\samples_imag[6][2] ),
    .S(_04859_),
    .Z(_04860_));
 MUX2_X1 _14015_ (.A(\samples_imag[5][2] ),
    .B(\samples_imag[7][2] ),
    .S(_04859_),
    .Z(_04861_));
 BUF_X4 _14016_ (.A(_04810_),
    .Z(_04862_));
 MUX2_X1 _14017_ (.A(_04860_),
    .B(_04861_),
    .S(_04862_),
    .Z(_04863_));
 AOI21_X4 _14018_ (.A(_04858_),
    .B1(_04863_),
    .B2(_04847_),
    .ZN(_04864_));
 OR2_X4 _14019_ (.A1(_04850_),
    .A2(_04864_),
    .ZN(_07702_));
 INV_X2 _14020_ (.A(_07702_),
    .ZN(_07443_));
 INV_X1 _14021_ (.A(_00023_),
    .ZN(_04865_));
 NOR2_X4 _14022_ (.A1(_04865_),
    .A2(_04849_),
    .ZN(_07372_));
 INV_X2 _14023_ (.A(_07372_),
    .ZN(_07498_));
 OR2_X1 _14024_ (.A1(_04808_),
    .A2(_04864_),
    .ZN(_07499_));
 INV_X2 _14025_ (.A(_07499_),
    .ZN(_07373_));
 BUF_X8 _14026_ (.A(_04837_),
    .Z(_04866_));
 BUF_X4 _14027_ (.A(_04830_),
    .Z(_04867_));
 BUF_X4 _14028_ (.A(_04867_),
    .Z(_04868_));
 BUF_X16 _14029_ (.A(_04812_),
    .Z(_04869_));
 BUF_X16 _14030_ (.A(_04869_),
    .Z(_04870_));
 BUF_X16 _14031_ (.A(_04870_),
    .Z(_04871_));
 MUX2_X1 _14032_ (.A(\samples_imag[0][3] ),
    .B(\samples_imag[2][3] ),
    .S(_04871_),
    .Z(_04872_));
 NOR2_X2 _14033_ (.A1(_04868_),
    .A2(_04872_),
    .ZN(_04873_));
 CLKBUF_X3 _14034_ (.A(_04855_),
    .Z(_04874_));
 BUF_X8 _14035_ (.A(_04840_),
    .Z(_04875_));
 MUX2_X1 _14036_ (.A(\samples_imag[1][3] ),
    .B(\samples_imag[3][3] ),
    .S(_04875_),
    .Z(_04876_));
 NOR2_X1 _14037_ (.A1(_04874_),
    .A2(_04876_),
    .ZN(_04877_));
 NOR3_X2 _14038_ (.A1(_04866_),
    .A2(_04873_),
    .A3(_04877_),
    .ZN(_04878_));
 MUX2_X1 _14039_ (.A(\samples_imag[4][3] ),
    .B(\samples_imag[6][3] ),
    .S(_04871_),
    .Z(_04879_));
 MUX2_X1 _14040_ (.A(\samples_imag[5][3] ),
    .B(\samples_imag[7][3] ),
    .S(_04871_),
    .Z(_04880_));
 MUX2_X1 _14041_ (.A(_04879_),
    .B(_04880_),
    .S(_04868_),
    .Z(_04881_));
 AOI21_X4 _14042_ (.A(_04878_),
    .B1(_04881_),
    .B2(_04866_),
    .ZN(_04882_));
 NOR2_X2 _14043_ (.A1(_04808_),
    .A2(_04882_),
    .ZN(_07374_));
 BUF_X16 _14044_ (.A(_04812_),
    .Z(_04883_));
 BUF_X8 _14045_ (.A(_04883_),
    .Z(_04884_));
 MUX2_X1 _14046_ (.A(\samples_imag[0][4] ),
    .B(\samples_imag[2][4] ),
    .S(_04884_),
    .Z(_04885_));
 NOR2_X1 _14047_ (.A1(_04867_),
    .A2(_04885_),
    .ZN(_04886_));
 MUX2_X1 _14048_ (.A(\samples_imag[1][4] ),
    .B(\samples_imag[3][4] ),
    .S(_04884_),
    .Z(_04887_));
 NOR2_X1 _14049_ (.A1(_04874_),
    .A2(_04887_),
    .ZN(_04888_));
 NOR3_X2 _14050_ (.A1(_04837_),
    .A2(_04886_),
    .A3(_04888_),
    .ZN(_04889_));
 MUX2_X1 _14051_ (.A(\samples_imag[4][4] ),
    .B(\samples_imag[6][4] ),
    .S(net53),
    .Z(_04890_));
 MUX2_X1 _14052_ (.A(\samples_imag[5][4] ),
    .B(\samples_imag[7][4] ),
    .S(_04870_),
    .Z(_04891_));
 MUX2_X1 _14053_ (.A(_04890_),
    .B(_04891_),
    .S(_04867_),
    .Z(_04892_));
 BUF_X8 _14054_ (.A(_04847_),
    .Z(_04893_));
 AOI21_X4 _14055_ (.A(_04889_),
    .B1(_04892_),
    .B2(_04893_),
    .ZN(_04894_));
 NOR2_X2 _14056_ (.A1(_04808_),
    .A2(_04894_),
    .ZN(_07409_));
 BUF_X4 _14057_ (.A(_04850_),
    .Z(_04895_));
 BUF_X4 _14058_ (.A(net51),
    .Z(_04896_));
 MUX2_X1 _14059_ (.A(\samples_imag[0][5] ),
    .B(\samples_imag[2][5] ),
    .S(_04896_),
    .Z(_04897_));
 NOR2_X1 _14060_ (.A1(_04862_),
    .A2(_04897_),
    .ZN(_04898_));
 MUX2_X1 _14061_ (.A(\samples_imag[1][5] ),
    .B(\samples_imag[3][5] ),
    .S(_04896_),
    .Z(_04899_));
 NOR2_X1 _14062_ (.A1(_04815_),
    .A2(_04899_),
    .ZN(_04900_));
 NOR3_X2 _14063_ (.A1(_04836_),
    .A2(_04898_),
    .A3(_04900_),
    .ZN(_04901_));
 MUX2_X1 _14064_ (.A(\samples_imag[4][5] ),
    .B(\samples_imag[6][5] ),
    .S(_04826_),
    .Z(_04902_));
 MUX2_X1 _14065_ (.A(\samples_imag[5][5] ),
    .B(\samples_imag[7][5] ),
    .S(_04826_),
    .Z(_04903_));
 MUX2_X1 _14066_ (.A(_04902_),
    .B(_04903_),
    .S(_04810_),
    .Z(_04904_));
 BUF_X8 _14067_ (.A(_04809_),
    .Z(_04905_));
 AOI21_X4 _14068_ (.A(_04901_),
    .B1(_04904_),
    .B2(_04905_),
    .ZN(_04906_));
 NOR2_X4 _14069_ (.A1(_04895_),
    .A2(_04906_),
    .ZN(_07410_));
 BUF_X4 _14070_ (.A(_04895_),
    .Z(_04907_));
 NOR2_X4 _14071_ (.A1(_04907_),
    .A2(_04894_),
    .ZN(_07381_));
 NOR2_X1 _14072_ (.A1(_04808_),
    .A2(_04906_),
    .ZN(_07382_));
 MUX2_X1 _14073_ (.A(\samples_imag[0][6] ),
    .B(\samples_imag[2][6] ),
    .S(_04871_),
    .Z(_04908_));
 MUX2_X1 _14074_ (.A(\samples_imag[1][6] ),
    .B(\samples_imag[3][6] ),
    .S(_04871_),
    .Z(_04909_));
 MUX2_X1 _14075_ (.A(_04908_),
    .B(_04909_),
    .S(_04868_),
    .Z(_04910_));
 BUF_X16 _14076_ (.A(_04871_),
    .Z(_04911_));
 MUX2_X1 _14077_ (.A(\samples_imag[4][6] ),
    .B(\samples_imag[6][6] ),
    .S(_04911_),
    .Z(_04912_));
 MUX2_X1 _14078_ (.A(\samples_imag[5][6] ),
    .B(\samples_imag[7][6] ),
    .S(_04911_),
    .Z(_04913_));
 MUX2_X1 _14079_ (.A(_04912_),
    .B(_04913_),
    .S(_04868_),
    .Z(_04914_));
 MUX2_X2 _14080_ (.A(_04910_),
    .B(_04914_),
    .S(_04866_),
    .Z(_04915_));
 INV_X4 _14081_ (.A(_04915_),
    .ZN(_04916_));
 NOR2_X4 _14082_ (.A1(_04916_),
    .A2(_04907_),
    .ZN(_07383_));
 OR2_X2 _14083_ (.A1(_04907_),
    .A2(_04822_),
    .ZN(_07853_));
 INV_X4 _14084_ (.A(_07853_),
    .ZN(_07378_));
 MUX2_X1 _14085_ (.A(\samples_real[0][12] ),
    .B(\samples_real[2][12] ),
    .S(_04896_),
    .Z(_04917_));
 NOR2_X1 _14086_ (.A1(_04862_),
    .A2(_04917_),
    .ZN(_04918_));
 MUX2_X1 _14087_ (.A(\samples_real[1][12] ),
    .B(\samples_real[3][12] ),
    .S(_04896_),
    .Z(_04919_));
 NOR2_X1 _14088_ (.A1(_04815_),
    .A2(_04919_),
    .ZN(_04920_));
 NOR3_X2 _14089_ (.A1(_04836_),
    .A2(_04918_),
    .A3(_04920_),
    .ZN(_04921_));
 MUX2_X1 _14090_ (.A(\samples_real[4][12] ),
    .B(\samples_real[6][12] ),
    .S(_04852_),
    .Z(_04922_));
 MUX2_X1 _14091_ (.A(\samples_real[5][12] ),
    .B(\samples_real[7][12] ),
    .S(_04852_),
    .Z(_04923_));
 MUX2_X1 _14092_ (.A(_04922_),
    .B(_04923_),
    .S(_04810_),
    .Z(_04924_));
 AOI21_X4 _14093_ (.A(_04921_),
    .B1(_04924_),
    .B2(_04905_),
    .ZN(_04925_));
 NOR2_X2 _14094_ (.A1(_04825_),
    .A2(_04925_),
    .ZN(_07481_));
 OR2_X2 _14095_ (.A1(_04907_),
    .A2(_04882_),
    .ZN(_07500_));
 INV_X2 _14096_ (.A(_07500_),
    .ZN(_07411_));
 AND2_X1 _14097_ (.A1(_00024_),
    .A2(_04915_),
    .ZN(_09390_));
 INV_X1 _14098_ (.A(_09390_),
    .ZN(_07422_));
 MUX2_X1 _14099_ (.A(\samples_imag[0][7] ),
    .B(\samples_imag[2][7] ),
    .S(_04827_),
    .Z(_04926_));
 NOR2_X1 _14100_ (.A1(_04834_),
    .A2(_04926_),
    .ZN(_04927_));
 MUX2_X1 _14101_ (.A(\samples_imag[1][7] ),
    .B(\samples_imag[3][7] ),
    .S(_04840_),
    .Z(_04928_));
 NOR2_X1 _14102_ (.A1(_04855_),
    .A2(_04928_),
    .ZN(_04929_));
 NOR3_X2 _14103_ (.A1(_04837_),
    .A2(_04927_),
    .A3(_04929_),
    .ZN(_04930_));
 MUX2_X1 _14104_ (.A(\samples_imag[4][7] ),
    .B(\samples_imag[6][7] ),
    .S(_04884_),
    .Z(_04931_));
 MUX2_X1 _14105_ (.A(\samples_imag[5][7] ),
    .B(\samples_imag[7][7] ),
    .S(_04884_),
    .Z(_04932_));
 MUX2_X1 _14106_ (.A(_04931_),
    .B(_04932_),
    .S(_04834_),
    .Z(_04933_));
 AOI21_X4 _14107_ (.A(_04930_),
    .B1(_04933_),
    .B2(_04893_),
    .ZN(_04934_));
 OR2_X2 _14108_ (.A1(_04907_),
    .A2(_04934_),
    .ZN(_07423_));
 INV_X2 _14109_ (.A(_07423_),
    .ZN(_07449_));
 INV_X1 _14110_ (.A(_04934_),
    .ZN(_04935_));
 NAND2_X1 _14111_ (.A1(_00024_),
    .A2(_04935_),
    .ZN(_07396_));
 MUX2_X1 _14112_ (.A(\samples_imag[0][8] ),
    .B(\samples_imag[2][8] ),
    .S(_04870_),
    .Z(_04936_));
 NOR2_X1 _14113_ (.A1(_04867_),
    .A2(_04936_),
    .ZN(_04937_));
 MUX2_X1 _14114_ (.A(\samples_imag[1][8] ),
    .B(\samples_imag[3][8] ),
    .S(_04870_),
    .Z(_04938_));
 NOR2_X1 _14115_ (.A1(_04874_),
    .A2(_04938_),
    .ZN(_04939_));
 NOR3_X2 _14116_ (.A1(_04893_),
    .A2(_04937_),
    .A3(_04939_),
    .ZN(_04940_));
 MUX2_X1 _14117_ (.A(\samples_imag[4][8] ),
    .B(\samples_imag[6][8] ),
    .S(_04875_),
    .Z(_04941_));
 MUX2_X1 _14118_ (.A(\samples_imag[5][8] ),
    .B(\samples_imag[7][8] ),
    .S(_04875_),
    .Z(_04942_));
 MUX2_X1 _14119_ (.A(_04941_),
    .B(_04942_),
    .S(_04867_),
    .Z(_04943_));
 AOI21_X4 _14120_ (.A(_04940_),
    .B1(_04943_),
    .B2(_04893_),
    .ZN(_04944_));
 OR2_X2 _14121_ (.A1(_04907_),
    .A2(_04944_),
    .ZN(_07397_));
 INV_X1 _14122_ (.A(_07397_),
    .ZN(_07552_));
 MUX2_X1 _14123_ (.A(\samples_imag[0][9] ),
    .B(\samples_imag[2][9] ),
    .S(_04871_),
    .Z(_04945_));
 NOR2_X1 _14124_ (.A1(_04868_),
    .A2(_04945_),
    .ZN(_04946_));
 MUX2_X1 _14125_ (.A(\samples_imag[1][9] ),
    .B(\samples_imag[3][9] ),
    .S(_04871_),
    .Z(_04947_));
 NOR2_X1 _14126_ (.A1(_04874_),
    .A2(_04947_),
    .ZN(_04948_));
 NOR3_X2 _14127_ (.A1(_04866_),
    .A2(_04946_),
    .A3(_04948_),
    .ZN(_04949_));
 MUX2_X1 _14128_ (.A(\samples_imag[4][9] ),
    .B(\samples_imag[6][9] ),
    .S(_04911_),
    .Z(_04950_));
 MUX2_X1 _14129_ (.A(\samples_imag[5][9] ),
    .B(\samples_imag[7][9] ),
    .S(_04911_),
    .Z(_04951_));
 MUX2_X1 _14130_ (.A(_04950_),
    .B(_04951_),
    .S(_04868_),
    .Z(_04952_));
 AOI21_X4 _14131_ (.A(_04949_),
    .B1(_04952_),
    .B2(_04866_),
    .ZN(_04953_));
 OR2_X2 _14132_ (.A1(_04907_),
    .A2(_04953_),
    .ZN(_07398_));
 INV_X1 _14133_ (.A(_07398_),
    .ZN(_07391_));
 MUX2_X1 _14134_ (.A(\samples_imag[0][10] ),
    .B(\samples_imag[2][10] ),
    .S(_04871_),
    .Z(_04954_));
 NOR2_X1 _14135_ (.A1(_04868_),
    .A2(_04954_),
    .ZN(_04955_));
 MUX2_X1 _14136_ (.A(\samples_imag[1][10] ),
    .B(\samples_imag[3][10] ),
    .S(_04871_),
    .Z(_04956_));
 NOR2_X1 _14137_ (.A1(_04874_),
    .A2(_04956_),
    .ZN(_04957_));
 NOR3_X2 _14138_ (.A1(_04866_),
    .A2(_04955_),
    .A3(_04957_),
    .ZN(_04958_));
 MUX2_X1 _14139_ (.A(\samples_imag[4][10] ),
    .B(\samples_imag[6][10] ),
    .S(_04911_),
    .Z(_04959_));
 MUX2_X1 _14140_ (.A(\samples_imag[5][10] ),
    .B(\samples_imag[7][10] ),
    .S(_04911_),
    .Z(_04960_));
 MUX2_X1 _14141_ (.A(_04959_),
    .B(_04960_),
    .S(_04868_),
    .Z(_04961_));
 AOI21_X4 _14142_ (.A(_04958_),
    .B1(_04866_),
    .B2(_04961_),
    .ZN(_04962_));
 OR2_X1 _14143_ (.A1(_04907_),
    .A2(_04962_),
    .ZN(_07451_));
 INV_X1 _14144_ (.A(_07451_),
    .ZN(_07392_));
 MUX2_X1 _14145_ (.A(\samples_imag[0][11] ),
    .B(\samples_imag[2][11] ),
    .S(_04911_),
    .Z(_04963_));
 NOR2_X1 _14146_ (.A1(_04868_),
    .A2(_04963_),
    .ZN(_04964_));
 MUX2_X1 _14147_ (.A(\samples_imag[1][11] ),
    .B(\samples_imag[3][11] ),
    .S(_04911_),
    .Z(_04965_));
 NOR2_X1 _14148_ (.A1(_04874_),
    .A2(_04965_),
    .ZN(_04966_));
 NOR3_X2 _14149_ (.A1(_04866_),
    .A2(_04964_),
    .A3(_04966_),
    .ZN(_04967_));
 MUX2_X1 _14150_ (.A(\samples_imag[4][11] ),
    .B(\samples_imag[6][11] ),
    .S(_04911_),
    .Z(_04968_));
 MUX2_X1 _14151_ (.A(\samples_imag[5][11] ),
    .B(\samples_imag[7][11] ),
    .S(_04911_),
    .Z(_04969_));
 MUX2_X1 _14152_ (.A(_04968_),
    .B(_04969_),
    .S(_04868_),
    .Z(_04970_));
 AOI21_X4 _14153_ (.A(_04967_),
    .B1(_04970_),
    .B2(_04866_),
    .ZN(_04971_));
 NOR2_X1 _14154_ (.A1(_04907_),
    .A2(_04971_),
    .ZN(_07393_));
 MUX2_X1 _14155_ (.A(\samples_imag[0][12] ),
    .B(\samples_imag[2][12] ),
    .S(_04884_),
    .Z(_04972_));
 NOR2_X1 _14156_ (.A1(_04867_),
    .A2(_04972_),
    .ZN(_04973_));
 MUX2_X1 _14157_ (.A(\samples_imag[1][12] ),
    .B(\samples_imag[3][12] ),
    .S(_04884_),
    .Z(_04974_));
 NOR2_X1 _14158_ (.A1(_04874_),
    .A2(_04974_),
    .ZN(_04975_));
 NOR3_X2 _14159_ (.A1(_04837_),
    .A2(_04973_),
    .A3(_04975_),
    .ZN(_04976_));
 MUX2_X1 _14160_ (.A(\samples_imag[4][12] ),
    .B(\samples_imag[6][12] ),
    .S(net53),
    .Z(_04977_));
 MUX2_X1 _14161_ (.A(\samples_imag[5][12] ),
    .B(\samples_imag[7][12] ),
    .S(net53),
    .Z(_04978_));
 MUX2_X1 _14162_ (.A(_04977_),
    .B(_04978_),
    .S(_04834_),
    .Z(_04979_));
 AOI21_X4 _14163_ (.A(_04976_),
    .B1(_04979_),
    .B2(_04893_),
    .ZN(_04980_));
 NOR2_X1 _14164_ (.A1(_04895_),
    .A2(_04980_),
    .ZN(_07401_));
 INV_X4 _14165_ (.A(_04823_),
    .ZN(_04981_));
 MUX2_X1 _14166_ (.A(\samples_real[0][11] ),
    .B(\samples_real[2][11] ),
    .S(_04896_),
    .Z(_04982_));
 NOR2_X1 _14167_ (.A1(_04810_),
    .A2(_04982_),
    .ZN(_04983_));
 MUX2_X1 _14168_ (.A(\samples_real[1][11] ),
    .B(\samples_real[3][11] ),
    .S(_04896_),
    .Z(_04984_));
 NOR2_X1 _14169_ (.A1(_04815_),
    .A2(_04984_),
    .ZN(_04985_));
 NOR3_X2 _14170_ (.A1(_04836_),
    .A2(_04983_),
    .A3(_04985_),
    .ZN(_04986_));
 MUX2_X1 _14171_ (.A(\samples_real[4][11] ),
    .B(\samples_real[6][11] ),
    .S(_04852_),
    .Z(_04987_));
 MUX2_X1 _14172_ (.A(\samples_real[5][11] ),
    .B(\samples_real[7][11] ),
    .S(_04826_),
    .Z(_04988_));
 MUX2_X1 _14173_ (.A(_04987_),
    .B(_04988_),
    .S(_04810_),
    .Z(_04989_));
 AOI21_X2 _14174_ (.A(_04986_),
    .B1(_04989_),
    .B2(_04905_),
    .ZN(_04990_));
 INV_X1 _14175_ (.A(_04990_),
    .ZN(_04991_));
 NAND2_X1 _14176_ (.A1(_04981_),
    .A2(_04991_),
    .ZN(_07471_));
 INV_X1 _14177_ (.A(_07471_),
    .ZN(_07529_));
 CLKBUF_X3 _14178_ (.A(_00036_),
    .Z(_04992_));
 MUX2_X1 _14179_ (.A(\samples_imag[0][13] ),
    .B(\samples_imag[2][13] ),
    .S(_04827_),
    .Z(_04993_));
 NOR2_X1 _14180_ (.A1(_04834_),
    .A2(_04993_),
    .ZN(_04994_));
 MUX2_X1 _14181_ (.A(\samples_imag[1][13] ),
    .B(\samples_imag[3][13] ),
    .S(_04827_),
    .Z(_04995_));
 NOR2_X1 _14182_ (.A1(_04874_),
    .A2(_04995_),
    .ZN(_04996_));
 NOR3_X2 _14183_ (.A1(_04837_),
    .A2(_04994_),
    .A3(_04996_),
    .ZN(_04997_));
 MUX2_X1 _14184_ (.A(\samples_imag[4][13] ),
    .B(\samples_imag[6][13] ),
    .S(net53),
    .Z(_04998_));
 MUX2_X1 _14185_ (.A(\samples_imag[5][13] ),
    .B(\samples_imag[7][13] ),
    .S(net53),
    .Z(_04999_));
 MUX2_X1 _14186_ (.A(_04998_),
    .B(_04999_),
    .S(_04834_),
    .Z(_05000_));
 AOI21_X4 _14187_ (.A(_04997_),
    .B1(_05000_),
    .B2(_04893_),
    .ZN(_05001_));
 NOR2_X1 _14188_ (.A1(_04992_),
    .A2(_05001_),
    .ZN(_09394_));
 MUX2_X1 _14189_ (.A(\samples_imag[0][14] ),
    .B(\samples_imag[2][14] ),
    .S(_04883_),
    .Z(_05002_));
 NOR2_X1 _14190_ (.A1(_04830_),
    .A2(_05002_),
    .ZN(_05003_));
 MUX2_X1 _14191_ (.A(\samples_imag[1][14] ),
    .B(\samples_imag[3][14] ),
    .S(_04883_),
    .Z(_05004_));
 NOR2_X1 _14192_ (.A1(_04855_),
    .A2(_05004_),
    .ZN(_05005_));
 NOR3_X2 _14193_ (.A1(_04905_),
    .A2(_05003_),
    .A3(_05005_),
    .ZN(_05006_));
 MUX2_X1 _14194_ (.A(\samples_imag[4][14] ),
    .B(\samples_imag[6][14] ),
    .S(net52),
    .Z(_05007_));
 MUX2_X1 _14195_ (.A(\samples_imag[5][14] ),
    .B(\samples_imag[7][14] ),
    .S(_04869_),
    .Z(_05008_));
 MUX2_X1 _14196_ (.A(_05007_),
    .B(_05008_),
    .S(_04830_),
    .Z(_05009_));
 AOI21_X4 _14197_ (.A(_05006_),
    .B1(_05009_),
    .B2(_04837_),
    .ZN(_05010_));
 NOR2_X1 _14198_ (.A1(_00037_),
    .A2(_05010_),
    .ZN(_09395_));
 MUX2_X1 _14199_ (.A(\samples_real[0][2] ),
    .B(\samples_real[2][2] ),
    .S(_04827_),
    .Z(_05011_));
 NOR2_X2 _14200_ (.A1(_04834_),
    .A2(_05011_),
    .ZN(_05012_));
 MUX2_X1 _14201_ (.A(\samples_real[1][2] ),
    .B(\samples_real[3][2] ),
    .S(_04827_),
    .Z(_05013_));
 NOR2_X2 _14202_ (.A1(_04874_),
    .A2(_05013_),
    .ZN(_05014_));
 NOR3_X2 _14203_ (.A1(_04837_),
    .A2(_05012_),
    .A3(_05014_),
    .ZN(_05015_));
 MUX2_X1 _14204_ (.A(\samples_real[4][2] ),
    .B(\samples_real[6][2] ),
    .S(_04884_),
    .Z(_05016_));
 MUX2_X1 _14205_ (.A(\samples_real[5][2] ),
    .B(\samples_real[7][2] ),
    .S(_04884_),
    .Z(_05017_));
 MUX2_X1 _14206_ (.A(_05016_),
    .B(_05017_),
    .S(_04834_),
    .Z(_05018_));
 AOI21_X4 _14207_ (.A(_05015_),
    .B1(_05018_),
    .B2(_04893_),
    .ZN(_05019_));
 NOR2_X4 _14208_ (.A1(_04823_),
    .A2(_05019_),
    .ZN(_07559_));
 MUX2_X1 _14209_ (.A(\samples_real[0][1] ),
    .B(\samples_real[2][1] ),
    .S(_04827_),
    .Z(_05020_));
 NOR2_X1 _14210_ (.A1(_04834_),
    .A2(_05020_),
    .ZN(_05021_));
 MUX2_X1 _14211_ (.A(\samples_real[1][1] ),
    .B(\samples_real[3][1] ),
    .S(_04840_),
    .Z(_05022_));
 NOR2_X1 _14212_ (.A1(_04855_),
    .A2(_05022_),
    .ZN(_05023_));
 NOR3_X2 _14213_ (.A1(_04837_),
    .A2(_05021_),
    .A3(_05023_),
    .ZN(_05024_));
 MUX2_X1 _14214_ (.A(\samples_real[4][1] ),
    .B(\samples_real[6][1] ),
    .S(_04884_),
    .Z(_05025_));
 MUX2_X1 _14215_ (.A(\samples_real[5][1] ),
    .B(\samples_real[7][1] ),
    .S(_04884_),
    .Z(_05026_));
 MUX2_X1 _14216_ (.A(_05025_),
    .B(_05026_),
    .S(_04834_),
    .Z(_05027_));
 AOI21_X4 _14217_ (.A(_05024_),
    .B1(_04893_),
    .B2(_05027_),
    .ZN(_05028_));
 NOR2_X4 _14218_ (.A1(_04825_),
    .A2(_05028_),
    .ZN(_07603_));
 MUX2_X1 _14219_ (.A(\samples_real[0][4] ),
    .B(\samples_real[2][4] ),
    .S(_04852_),
    .Z(_05029_));
 NOR2_X1 _14220_ (.A1(_04862_),
    .A2(_05029_),
    .ZN(_05030_));
 MUX2_X1 _14221_ (.A(\samples_real[1][4] ),
    .B(\samples_real[3][4] ),
    .S(_04896_),
    .Z(_05031_));
 NOR2_X1 _14222_ (.A1(_04815_),
    .A2(_05031_),
    .ZN(_05032_));
 NOR3_X2 _14223_ (.A1(_04836_),
    .A2(_05030_),
    .A3(_05032_),
    .ZN(_05033_));
 MUX2_X1 _14224_ (.A(\samples_real[4][4] ),
    .B(\samples_real[6][4] ),
    .S(_04859_),
    .Z(_05034_));
 MUX2_X1 _14225_ (.A(\samples_real[5][4] ),
    .B(\samples_real[7][4] ),
    .S(_04859_),
    .Z(_05035_));
 MUX2_X1 _14226_ (.A(_05034_),
    .B(_05035_),
    .S(_04862_),
    .Z(_05036_));
 AOI21_X4 _14227_ (.A(_05033_),
    .B1(_05036_),
    .B2(_04847_),
    .ZN(_05037_));
 NOR2_X4 _14228_ (.A1(_04825_),
    .A2(_05037_),
    .ZN(_07671_));
 MUX2_X1 _14229_ (.A(\samples_real[0][10] ),
    .B(\samples_real[2][10] ),
    .S(_04875_),
    .Z(_05038_));
 NOR2_X1 _14230_ (.A1(_04867_),
    .A2(_05038_),
    .ZN(_05039_));
 MUX2_X1 _14231_ (.A(\samples_real[1][10] ),
    .B(\samples_real[3][10] ),
    .S(_04870_),
    .Z(_05040_));
 NOR2_X1 _14232_ (.A1(_04874_),
    .A2(_05040_),
    .ZN(_05041_));
 NOR3_X2 _14233_ (.A1(_04893_),
    .A2(_05039_),
    .A3(_05041_),
    .ZN(_05042_));
 MUX2_X1 _14234_ (.A(\samples_real[4][10] ),
    .B(\samples_real[6][10] ),
    .S(_04875_),
    .Z(_05043_));
 MUX2_X1 _14235_ (.A(\samples_real[5][10] ),
    .B(\samples_real[7][10] ),
    .S(_04875_),
    .Z(_05044_));
 MUX2_X1 _14236_ (.A(_05043_),
    .B(_05044_),
    .S(_04867_),
    .Z(_05045_));
 AOI21_X4 _14237_ (.A(_05042_),
    .B1(_04866_),
    .B2(_05045_),
    .ZN(_05046_));
 NOR2_X4 _14238_ (.A1(_04825_),
    .A2(_05046_),
    .ZN(_07472_));
 MUX2_X1 _14239_ (.A(\samples_real[0][0] ),
    .B(\samples_real[2][0] ),
    .S(_04826_),
    .Z(_05047_));
 NOR2_X1 _14240_ (.A1(_04851_),
    .A2(_05047_),
    .ZN(_05048_));
 MUX2_X1 _14241_ (.A(\samples_real[1][0] ),
    .B(\samples_real[3][0] ),
    .S(_04826_),
    .Z(_05049_));
 NOR2_X1 _14242_ (.A1(_04855_),
    .A2(_05049_),
    .ZN(_05050_));
 NOR3_X2 _14243_ (.A1(_04905_),
    .A2(_05048_),
    .A3(_05050_),
    .ZN(_05051_));
 MUX2_X1 _14244_ (.A(\samples_real[4][0] ),
    .B(\samples_real[6][0] ),
    .S(_04883_),
    .Z(_05052_));
 MUX2_X1 _14245_ (.A(\samples_real[5][0] ),
    .B(\samples_real[7][0] ),
    .S(_04883_),
    .Z(_05053_));
 MUX2_X1 _14246_ (.A(_05052_),
    .B(_05053_),
    .S(_04851_),
    .Z(_05054_));
 AOI21_X4 _14247_ (.A(_05051_),
    .B1(_05054_),
    .B2(_04847_),
    .ZN(_05055_));
 NOR2_X4 _14248_ (.A1(_04823_),
    .A2(_05055_),
    .ZN(_07653_));
 MUX2_X1 _14249_ (.A(\samples_real[0][3] ),
    .B(\samples_real[2][3] ),
    .S(_04852_),
    .Z(_05056_));
 NOR2_X1 _14250_ (.A1(_04851_),
    .A2(_05056_),
    .ZN(_05057_));
 MUX2_X1 _14251_ (.A(\samples_real[1][3] ),
    .B(\samples_real[3][3] ),
    .S(_04896_),
    .Z(_05058_));
 NOR2_X1 _14252_ (.A1(_04855_),
    .A2(_05058_),
    .ZN(_05059_));
 NOR3_X2 _14253_ (.A1(_04836_),
    .A2(_05057_),
    .A3(_05059_),
    .ZN(_05060_));
 MUX2_X1 _14254_ (.A(\samples_real[4][3] ),
    .B(\samples_real[6][3] ),
    .S(_04859_),
    .Z(_05061_));
 MUX2_X1 _14255_ (.A(\samples_real[5][3] ),
    .B(\samples_real[7][3] ),
    .S(_04859_),
    .Z(_05062_));
 MUX2_X1 _14256_ (.A(_05061_),
    .B(_05062_),
    .S(_04862_),
    .Z(_05063_));
 AOI21_X4 _14257_ (.A(_05060_),
    .B1(_05063_),
    .B2(_04847_),
    .ZN(_05064_));
 NOR2_X4 _14258_ (.A1(_04825_),
    .A2(_05064_),
    .ZN(_07718_));
 MUX2_X1 _14259_ (.A(\samples_real[0][5] ),
    .B(\samples_real[2][5] ),
    .S(_04826_),
    .Z(_05065_));
 NOR2_X1 _14260_ (.A1(_04851_),
    .A2(_05065_),
    .ZN(_05066_));
 MUX2_X1 _14261_ (.A(\samples_real[1][5] ),
    .B(\samples_real[3][5] ),
    .S(_04852_),
    .Z(_05067_));
 NOR2_X1 _14262_ (.A1(_04855_),
    .A2(_05067_),
    .ZN(_05068_));
 NOR3_X2 _14263_ (.A1(_04905_),
    .A2(_05066_),
    .A3(_05068_),
    .ZN(_05069_));
 MUX2_X1 _14264_ (.A(\samples_real[4][5] ),
    .B(\samples_real[6][5] ),
    .S(_04883_),
    .Z(_05070_));
 MUX2_X1 _14265_ (.A(\samples_real[5][5] ),
    .B(\samples_real[7][5] ),
    .S(_04883_),
    .Z(_05071_));
 MUX2_X1 _14266_ (.A(_05070_),
    .B(_05071_),
    .S(_04851_),
    .Z(_05072_));
 AOI21_X4 _14267_ (.A(_05069_),
    .B1(_05072_),
    .B2(_04847_),
    .ZN(_05073_));
 NOR2_X4 _14268_ (.A1(_04825_),
    .A2(_05073_),
    .ZN(_07621_));
 MUX2_X1 _14269_ (.A(\samples_real[0][7] ),
    .B(\samples_real[2][7] ),
    .S(_04852_),
    .Z(_05074_));
 NOR2_X1 _14270_ (.A1(_04862_),
    .A2(_05074_),
    .ZN(_05075_));
 MUX2_X1 _14271_ (.A(\samples_real[1][7] ),
    .B(\samples_real[3][7] ),
    .S(_04896_),
    .Z(_05076_));
 NOR2_X1 _14272_ (.A1(_04815_),
    .A2(_05076_),
    .ZN(_05077_));
 NOR3_X2 _14273_ (.A1(_04836_),
    .A2(_05075_),
    .A3(_05077_),
    .ZN(_05078_));
 MUX2_X1 _14274_ (.A(\samples_real[4][7] ),
    .B(\samples_real[6][7] ),
    .S(_04826_),
    .Z(_05079_));
 MUX2_X1 _14275_ (.A(\samples_real[5][7] ),
    .B(\samples_real[7][7] ),
    .S(_04859_),
    .Z(_05080_));
 MUX2_X1 _14276_ (.A(_05079_),
    .B(_05080_),
    .S(_04862_),
    .Z(_05081_));
 AOI21_X4 _14277_ (.A(_05078_),
    .B1(_05081_),
    .B2(_04905_),
    .ZN(_05082_));
 NOR2_X4 _14278_ (.A1(_04825_),
    .A2(_05082_),
    .ZN(_07533_));
 MUX2_X1 _14279_ (.A(\samples_real[0][8] ),
    .B(\samples_real[2][8] ),
    .S(_04883_),
    .Z(_05083_));
 NOR2_X1 _14280_ (.A1(_04830_),
    .A2(_05083_),
    .ZN(_05084_));
 MUX2_X1 _14281_ (.A(\samples_real[1][8] ),
    .B(\samples_real[3][8] ),
    .S(_04859_),
    .Z(_05085_));
 NOR2_X1 _14282_ (.A1(_04855_),
    .A2(_05085_),
    .ZN(_05086_));
 NOR3_X2 _14283_ (.A1(_04905_),
    .A2(_05084_),
    .A3(_05086_),
    .ZN(_05087_));
 MUX2_X1 _14284_ (.A(\samples_real[4][8] ),
    .B(\samples_real[6][8] ),
    .S(_04869_),
    .Z(_05088_));
 MUX2_X1 _14285_ (.A(\samples_real[5][8] ),
    .B(\samples_real[7][8] ),
    .S(_04869_),
    .Z(_05089_));
 MUX2_X1 _14286_ (.A(_05088_),
    .B(_05089_),
    .S(_04851_),
    .Z(_05090_));
 AOI21_X4 _14287_ (.A(_05087_),
    .B1(_05090_),
    .B2(_04837_),
    .ZN(_05091_));
 NOR2_X4 _14288_ (.A1(_04825_),
    .A2(_05091_),
    .ZN(_07485_));
 MUX2_X1 _14289_ (.A(\samples_real[0][6] ),
    .B(\samples_real[2][6] ),
    .S(_04852_),
    .Z(_05092_));
 NOR2_X2 _14290_ (.A1(_04862_),
    .A2(_05092_),
    .ZN(_05093_));
 MUX2_X1 _14291_ (.A(\samples_real[1][6] ),
    .B(\samples_real[3][6] ),
    .S(_04896_),
    .Z(_05094_));
 NOR2_X2 _14292_ (.A1(_04815_),
    .A2(_05094_),
    .ZN(_05095_));
 NOR3_X4 _14293_ (.A1(_04836_),
    .A2(_05093_),
    .A3(_05095_),
    .ZN(_05096_));
 MUX2_X1 _14294_ (.A(\samples_real[4][6] ),
    .B(\samples_real[6][6] ),
    .S(_04826_),
    .Z(_05097_));
 MUX2_X1 _14295_ (.A(\samples_real[5][6] ),
    .B(\samples_real[7][6] ),
    .S(_04826_),
    .Z(_05098_));
 MUX2_X1 _14296_ (.A(_05097_),
    .B(_05098_),
    .S(_04862_),
    .Z(_05099_));
 AOI21_X4 _14297_ (.A(_05096_),
    .B1(_05099_),
    .B2(_04905_),
    .ZN(_05100_));
 NOR2_X4 _14298_ (.A1(_04825_),
    .A2(_05100_),
    .ZN(_07578_));
 MUX2_X1 _14299_ (.A(\samples_real[0][9] ),
    .B(\samples_real[2][9] ),
    .S(_04859_),
    .Z(_05101_));
 NOR2_X1 _14300_ (.A1(_04851_),
    .A2(_05101_),
    .ZN(_05102_));
 MUX2_X1 _14301_ (.A(\samples_real[1][9] ),
    .B(\samples_real[3][9] ),
    .S(_04859_),
    .Z(_05103_));
 NOR2_X1 _14302_ (.A1(_04855_),
    .A2(_05103_),
    .ZN(_05104_));
 NOR3_X4 _14303_ (.A1(_04905_),
    .A2(_05102_),
    .A3(_05104_),
    .ZN(_05105_));
 MUX2_X1 _14304_ (.A(\samples_real[4][9] ),
    .B(\samples_real[6][9] ),
    .S(_04883_),
    .Z(_05106_));
 MUX2_X1 _14305_ (.A(\samples_real[5][9] ),
    .B(\samples_real[7][9] ),
    .S(_04883_),
    .Z(_05107_));
 MUX2_X1 _14306_ (.A(_05106_),
    .B(_05107_),
    .S(_04851_),
    .Z(_05108_));
 AOI21_X4 _14307_ (.A(_05105_),
    .B1(_05108_),
    .B2(_04847_),
    .ZN(_05109_));
 NOR2_X4 _14308_ (.A1(_04824_),
    .A2(_05109_),
    .ZN(_07473_));
 AND2_X1 _14309_ (.A1(_09580_),
    .A2(_07653_),
    .ZN(_09581_));
 OR2_X4 _14310_ (.A1(_04823_),
    .A2(_04864_),
    .ZN(_08332_));
 INV_X2 _14311_ (.A(_08332_),
    .ZN(_08285_));
 NAND2_X4 _14312_ (.A1(_04981_),
    .A2(_04848_),
    .ZN(_08333_));
 INV_X4 _14313_ (.A(_08333_),
    .ZN(_08336_));
 OR2_X4 _14314_ (.A1(_04823_),
    .A2(_04906_),
    .ZN(_08105_));
 INV_X2 _14315_ (.A(_08105_),
    .ZN(_08108_));
 OR2_X2 _14316_ (.A1(_05046_),
    .A2(_04907_),
    .ZN(_08077_));
 INV_X1 _14317_ (.A(_08077_),
    .ZN(_07989_));
 OR2_X4 _14318_ (.A1(_04823_),
    .A2(_04822_),
    .ZN(_08424_));
 INV_X4 _14319_ (.A(_08424_),
    .ZN(_08426_));
 OR2_X4 _14320_ (.A1(_04824_),
    .A2(_04894_),
    .ZN(_08168_));
 INV_X2 _14321_ (.A(_08168_),
    .ZN(_07921_));
 NAND2_X4 _14322_ (.A1(_04981_),
    .A2(_04935_),
    .ZN(_07953_));
 INV_X1 _14323_ (.A(_07953_),
    .ZN(_07956_));
 NAND2_X4 _14324_ (.A1(_04981_),
    .A2(_04915_),
    .ZN(_08040_));
 INV_X2 _14325_ (.A(_08040_),
    .ZN(_08043_));
 OR2_X4 _14326_ (.A1(_04824_),
    .A2(_04944_),
    .ZN(_07928_));
 INV_X1 _14327_ (.A(_07928_),
    .ZN(_07933_));
 OR2_X4 _14328_ (.A1(_04953_),
    .A2(_04824_),
    .ZN(_07929_));
 INV_X2 _14329_ (.A(_07929_),
    .ZN(_07914_));
 OR2_X4 _14330_ (.A1(_04824_),
    .A2(_04962_),
    .ZN(_07930_));
 INV_X1 _14331_ (.A(_07930_),
    .ZN(_07915_));
 NOR2_X2 _14332_ (.A1(_04824_),
    .A2(_04971_),
    .ZN(_07916_));
 OR2_X4 _14333_ (.A1(_04824_),
    .A2(net437),
    .ZN(_08230_));
 INV_X2 _14334_ (.A(_08230_),
    .ZN(_08233_));
 NOR2_X2 _14335_ (.A1(_04824_),
    .A2(_04980_),
    .ZN(_09592_));
 NOR2_X1 _14336_ (.A1(_04824_),
    .A2(_05001_),
    .ZN(_09593_));
 OR2_X2 _14337_ (.A1(_05028_),
    .A2(_04807_),
    .ZN(_08126_));
 INV_X2 _14338_ (.A(_08126_),
    .ZN(_07967_));
 OR2_X2 _14339_ (.A1(_04895_),
    .A2(_05028_),
    .ZN(_08190_));
 INV_X2 _14340_ (.A(_08190_),
    .ZN(_08352_));
 OR2_X1 _14341_ (.A1(_04808_),
    .A2(_05055_),
    .ZN(_08191_));
 INV_X2 _14342_ (.A(_08191_),
    .ZN(_08054_));
 OR2_X4 _14343_ (.A1(_04850_),
    .A2(_05019_),
    .ZN(_08127_));
 INV_X2 _14344_ (.A(_08127_),
    .ZN(_08055_));
 OR2_X2 _14345_ (.A1(_04807_),
    .A2(_05064_),
    .ZN(_08004_));
 INV_X1 _14346_ (.A(_08004_),
    .ZN(_07939_));
 OR2_X4 _14347_ (.A1(_04808_),
    .A2(_05019_),
    .ZN(_08065_));
 INV_X1 _14348_ (.A(_08065_),
    .ZN(_07940_));
 OR2_X2 _14349_ (.A1(_04895_),
    .A2(_05037_),
    .ZN(_08005_));
 INV_X2 _14350_ (.A(_08005_),
    .ZN(_07941_));
 OR2_X2 _14351_ (.A1(_04850_),
    .A2(_05109_),
    .ZN(_08135_));
 INV_X1 _14352_ (.A(_08135_),
    .ZN(_07990_));
 OR2_X2 _14353_ (.A1(_04895_),
    .A2(_05055_),
    .ZN(_08536_));
 INV_X4 _14354_ (.A(_08536_),
    .ZN(_08234_));
 OR2_X2 _14355_ (.A1(_04895_),
    .A2(_05064_),
    .ZN(_08066_));
 INV_X2 _14356_ (.A(_08066_),
    .ZN(_07968_));
 OR2_X2 _14357_ (.A1(_04850_),
    .A2(_05073_),
    .ZN(_07985_));
 INV_X2 _14358_ (.A(_07985_),
    .ZN(_08133_));
 OR2_X2 _14359_ (.A1(_04850_),
    .A2(_05082_),
    .ZN(_08256_));
 INV_X2 _14360_ (.A(_08256_),
    .ZN(_08017_));
 OR2_X1 _14361_ (.A1(_05073_),
    .A2(_04808_),
    .ZN(_08006_));
 INV_X1 _14362_ (.A(_08006_),
    .ZN(_07976_));
 OR2_X2 _14363_ (.A1(_05100_),
    .A2(_04895_),
    .ZN(_08303_));
 INV_X2 _14364_ (.A(_08303_),
    .ZN(_07977_));
 NOR2_X1 _14365_ (.A1(_04808_),
    .A2(_05082_),
    .ZN(_07978_));
 OR2_X2 _14366_ (.A1(_04895_),
    .A2(_05091_),
    .ZN(_08198_));
 INV_X1 _14367_ (.A(_08198_),
    .ZN(_07991_));
 CLKBUF_X3 _14368_ (.A(_00022_),
    .Z(_05110_));
 MUX2_X1 _14369_ (.A(\samples_real[0][14] ),
    .B(\samples_real[2][14] ),
    .S(_04869_),
    .Z(_05111_));
 MUX2_X1 _14370_ (.A(\samples_real[1][14] ),
    .B(\samples_real[3][14] ),
    .S(_04840_),
    .Z(_05112_));
 MUX2_X1 _14371_ (.A(_05111_),
    .B(_05112_),
    .S(_04830_),
    .Z(_05113_));
 MUX2_X1 _14372_ (.A(\samples_real[4][14] ),
    .B(\samples_real[6][14] ),
    .S(_04840_),
    .Z(_05114_));
 MUX2_X1 _14373_ (.A(\samples_real[5][14] ),
    .B(\samples_real[7][14] ),
    .S(_04840_),
    .Z(_05115_));
 MUX2_X1 _14374_ (.A(_05114_),
    .B(_05115_),
    .S(_04830_),
    .Z(_05116_));
 MUX2_X1 _14375_ (.A(_05113_),
    .B(_05116_),
    .S(_04847_),
    .Z(_05117_));
 NAND2_X1 _14376_ (.A1(_05110_),
    .A2(_05117_),
    .ZN(_07995_));
 NAND2_X1 _14377_ (.A1(_05110_),
    .A2(_04838_),
    .ZN(_08020_));
 INV_X1 _14378_ (.A(_04925_),
    .ZN(_05118_));
 NAND2_X1 _14379_ (.A1(_05110_),
    .A2(_05118_),
    .ZN(_08078_));
 NAND2_X1 _14380_ (.A1(_05110_),
    .A2(_04991_),
    .ZN(_08136_));
 INV_X1 _14381_ (.A(_05046_),
    .ZN(_05119_));
 NAND2_X1 _14382_ (.A1(_05110_),
    .A2(_05119_),
    .ZN(_08199_));
 INV_X1 _14383_ (.A(_08242_),
    .ZN(_09637_));
 INV_X1 _14384_ (.A(_05109_),
    .ZN(_05120_));
 NAND2_X1 _14385_ (.A1(_05110_),
    .A2(_05120_),
    .ZN(_08257_));
 INV_X1 _14386_ (.A(_05091_),
    .ZN(_05121_));
 NAND2_X1 _14387_ (.A1(_05110_),
    .A2(_05121_),
    .ZN(_08304_));
 NOR2_X1 _14388_ (.A1(_04992_),
    .A2(_05100_),
    .ZN(_08355_));
 INV_X2 _14389_ (.A(_05110_),
    .ZN(_05122_));
 OR2_X1 _14390_ (.A1(_05122_),
    .A2(_05100_),
    .ZN(_08394_));
 INV_X1 _14391_ (.A(_05073_),
    .ZN(_05123_));
 NAND2_X1 _14392_ (.A1(_05110_),
    .A2(_05123_),
    .ZN(_08448_));
 NOR2_X1 _14393_ (.A1(_00037_),
    .A2(_05037_),
    .ZN(_08493_));
 NOR2_X1 _14394_ (.A1(_04992_),
    .A2(_05064_),
    .ZN(_08494_));
 OR2_X1 _14395_ (.A1(_05122_),
    .A2(_05064_),
    .ZN(_08515_));
 INV_X1 _14396_ (.A(_05019_),
    .ZN(_05124_));
 NAND2_X1 _14397_ (.A1(_05110_),
    .A2(_05124_),
    .ZN(_08537_));
 NOR3_X2 _14398_ (.A1(_00845_),
    .A2(_04775_),
    .A3(_00851_),
    .ZN(_00009_));
 INV_X1 _14399_ (.A(_09406_),
    .ZN(_07476_));
 INV_X1 _14400_ (.A(_09460_),
    .ZN(_07659_));
 INV_X1 _14401_ (.A(_09473_),
    .ZN(_07710_));
 INV_X1 _14402_ (.A(_09489_),
    .ZN(_07753_));
 INV_X1 _14403_ (.A(_09502_),
    .ZN(_07792_));
 INV_X1 _14404_ (.A(_09519_),
    .ZN(_07833_));
 INV_X1 _14405_ (.A(_07746_),
    .ZN(_07742_));
 INV_X1 _14406_ (.A(_09521_),
    .ZN(_07877_));
 OR2_X1 _14407_ (.A1(_04850_),
    .A2(_04925_),
    .ZN(_07994_));
 INV_X1 _14408_ (.A(_09600_),
    .ZN(_07999_));
 OR2_X2 _14409_ (.A1(_04807_),
    .A2(_05037_),
    .ZN(_07984_));
 INV_X1 _14410_ (.A(_08059_),
    .ZN(_08086_));
 INV_X1 _14411_ (.A(_08138_),
    .ZN(_08140_));
 INV_X1 _14412_ (.A(_08120_),
    .ZN(_08144_));
 INV_X1 _14413_ (.A(_08297_),
    .ZN(_08292_));
 INV_X1 _14414_ (.A(_08280_),
    .ZN(_08320_));
 INV_X1 _14415_ (.A(_08447_),
    .ZN(_08444_));
 INV_X1 _14416_ (.A(_08501_),
    .ZN(_08497_));
 INV_X1 _14417_ (.A(_08513_),
    .ZN(_08532_));
 INV_X1 _14418_ (.A(_08629_),
    .ZN(_07348_));
 INV_X1 _14419_ (.A(_08710_),
    .ZN(_07356_));
 INV_X1 _14420_ (.A(_09403_),
    .ZN(_07495_));
 INV_X1 _14421_ (.A(_09419_),
    .ZN(_07525_));
 INV_X1 _14422_ (.A(_09432_),
    .ZN(_07572_));
 INV_X1 _14423_ (.A(_09444_),
    .ZN(_07615_));
 INV_X1 _14424_ (.A(_09457_),
    .ZN(_07665_));
 INV_X1 _14425_ (.A(_09462_),
    .ZN(_07694_));
 INV_X1 _14426_ (.A(_09551_),
    .ZN(_07878_));
 INV_X1 _14427_ (.A(_09562_),
    .ZN(_07905_));
 INV_X1 _14428_ (.A(_07913_),
    .ZN(_07908_));
 INV_X1 _14429_ (.A(_09601_),
    .ZN(_08062_));
 INV_X1 _14430_ (.A(_09606_),
    .ZN(_08124_));
 INV_X1 _14431_ (.A(_08125_),
    .ZN(_08145_));
 INV_X1 _14432_ (.A(_09614_),
    .ZN(_08187_));
 INV_X1 _14433_ (.A(_09625_),
    .ZN(_08249_));
 INV_X1 _14434_ (.A(_08509_),
    .ZN(_08507_));
 INV_X1 _14435_ (.A(_08514_),
    .ZN(_08511_));
 INV_X1 _14436_ (.A(_08535_),
    .ZN(_08533_));
 INV_X1 _14437_ (.A(_08539_),
    .ZN(_08540_));
 INV_X1 _14438_ (.A(_08551_),
    .ZN(_08544_));
 INV_X1 _14439_ (.A(_09743_),
    .ZN(_08549_));
 INV_X2 _14440_ (.A(_08556_),
    .ZN(_07349_));
 INV_X2 _14441_ (.A(_08637_),
    .ZN(_07357_));
 INV_X1 _14442_ (.A(_09413_),
    .ZN(_07478_));
 INV_X1 _14443_ (.A(_09402_),
    .ZN(_07496_));
 INV_X1 _14444_ (.A(_09418_),
    .ZN(_07526_));
 INV_X1 _14445_ (.A(_09431_),
    .ZN(_07573_));
 INV_X1 _14446_ (.A(_09443_),
    .ZN(_07616_));
 INV_X1 _14447_ (.A(_09465_),
    .ZN(_07661_));
 INV_X1 _14448_ (.A(_09456_),
    .ZN(_07666_));
 INV_X1 _14449_ (.A(_09461_),
    .ZN(_07695_));
 INV_X1 _14450_ (.A(_09479_),
    .ZN(_07712_));
 INV_X1 _14451_ (.A(_07705_),
    .ZN(_07743_));
 INV_X1 _14452_ (.A(_09494_),
    .ZN(_07755_));
 INV_X1 _14453_ (.A(_09507_),
    .ZN(_07794_));
 INV_X1 _14454_ (.A(_09525_),
    .ZN(_07835_));
 INV_X1 _14455_ (.A(_09531_),
    .ZN(_07857_));
 INV_X1 _14456_ (.A(_09561_),
    .ZN(_07906_));
 OR2_X1 _14457_ (.A1(_04807_),
    .A2(_05100_),
    .ZN(_07986_));
 INV_X2 _14458_ (.A(_04992_),
    .ZN(_05125_));
 NAND2_X1 _14459_ (.A1(_05125_),
    .A2(_04838_),
    .ZN(_07996_));
 INV_X1 _14460_ (.A(_08011_),
    .ZN(_08001_));
 NAND2_X1 _14461_ (.A1(_05125_),
    .A2(_05118_),
    .ZN(_08021_));
 NAND2_X1 _14462_ (.A1(_05125_),
    .A2(_04991_),
    .ZN(_08079_));
 NAND2_X1 _14463_ (.A1(_05125_),
    .A2(_05119_),
    .ZN(_08137_));
 NAND2_X1 _14464_ (.A1(_05125_),
    .A2(_05120_),
    .ZN(_08200_));
 NAND2_X1 _14465_ (.A1(_05125_),
    .A2(_05121_),
    .ZN(_08258_));
 OR2_X1 _14466_ (.A1(_04992_),
    .A2(_05082_),
    .ZN(_08305_));
 NAND2_X1 _14467_ (.A1(_05125_),
    .A2(_05123_),
    .ZN(_08395_));
 OR2_X1 _14468_ (.A1(_04992_),
    .A2(_05037_),
    .ZN(_08449_));
 INV_X1 _14469_ (.A(_08502_),
    .ZN(_08498_));
 INV_X1 _14470_ (.A(_08500_),
    .ZN(_08512_));
 NAND2_X1 _14471_ (.A1(_05125_),
    .A2(_05124_),
    .ZN(_08516_));
 INV_X1 _14472_ (.A(_08519_),
    .ZN(_08524_));
 OR2_X1 _14473_ (.A1(_04992_),
    .A2(_05028_),
    .ZN(_08538_));
 INV_X1 _14474_ (.A(_08542_),
    .ZN(_08550_));
 INV_X1 _14475_ (.A(_07376_),
    .ZN(_09388_));
 INV_X1 _14476_ (.A(_07385_),
    .ZN(_07387_));
 INV_X1 _14477_ (.A(_07408_),
    .ZN(_07435_));
 INV_X1 _14478_ (.A(_07421_),
    .ZN(_07427_));
 INV_X1 _14479_ (.A(_07442_),
    .ZN(_07490_));
 INV_X1 _14480_ (.A(_07457_),
    .ZN(_07492_));
 INV_X1 _14481_ (.A(_07461_),
    .ZN(_07467_));
 INV_X1 _14482_ (.A(_07515_),
    .ZN(_07521_));
 INV_X1 _14483_ (.A(_07546_),
    .ZN(_07591_));
 INV_X1 _14484_ (.A(_07562_),
    .ZN(_07567_));
 INV_X1 _14485_ (.A(_07597_),
    .ZN(_07638_));
 INV_X1 _14486_ (.A(_07613_),
    .ZN(_07640_));
 INV_X1 _14487_ (.A(_07646_),
    .ZN(_07690_));
 INV_X1 _14488_ (.A(_07655_),
    .ZN(_07660_));
 INV_X1 _14489_ (.A(_07677_),
    .ZN(_07688_));
 INV_X1 _14490_ (.A(_07724_),
    .ZN(_07735_));
 INV_X1 _14491_ (.A(_07741_),
    .ZN(_07776_));
 INV_X1 _14492_ (.A(_07766_),
    .ZN(_07778_));
 INV_X1 _14493_ (.A(_07784_),
    .ZN(_07815_));
 INV_X1 _14494_ (.A(_07805_),
    .ZN(_07817_));
 INV_X1 _14495_ (.A(_07876_),
    .ZN(_07879_));
 INV_X1 _14496_ (.A(_07932_),
    .ZN(_07950_));
 INV_X1 _14497_ (.A(_07955_),
    .ZN(_08037_));
 INV_X1 _14498_ (.A(_07961_),
    .ZN(_07972_));
 INV_X1 _14499_ (.A(_07983_),
    .ZN(_08000_));
 INV_X1 _14500_ (.A(_08042_),
    .ZN(_08102_));
 INV_X1 _14501_ (.A(_08089_),
    .ZN(_08091_));
 INV_X1 _14502_ (.A(_08107_),
    .ZN(_08165_));
 INV_X1 _14503_ (.A(_08111_),
    .ZN(_08118_));
 INV_X1 _14504_ (.A(_08170_),
    .ZN(_08227_));
 INV_X1 _14505_ (.A(_08174_),
    .ZN(_08181_));
 INV_X1 _14506_ (.A(_08232_),
    .ZN(_09633_));
 INV_X1 _14507_ (.A(_08246_),
    .ZN(_08283_));
 INV_X1 _14508_ (.A(_08254_),
    .ZN(_08261_));
 INV_X1 _14509_ (.A(_08268_),
    .ZN(_08279_));
 INV_X1 _14510_ (.A(_08296_),
    .ZN(_08330_));
 INV_X1 _14511_ (.A(_08301_),
    .ZN(_08308_));
 INV_X1 _14512_ (.A(_08315_),
    .ZN(_08326_));
 INV_X2 _14513_ (.A(_08335_),
    .ZN(_09663_));
 INV_X1 _14514_ (.A(_08346_),
    .ZN(_08381_));
 INV_X1 _14515_ (.A(_08351_),
    .ZN(_08358_));
 INV_X1 _14516_ (.A(_08357_),
    .ZN(_08390_));
 INV_X1 _14517_ (.A(_08366_),
    .ZN(_08377_));
 INV_X1 _14518_ (.A(_08392_),
    .ZN(_08398_));
 INV_X1 _14519_ (.A(_08393_),
    .ZN(_08445_));
 INV_X1 _14520_ (.A(_08406_),
    .ZN(_08418_));
 INV_X1 _14521_ (.A(_08425_),
    .ZN(_09690_));
 INV_X1 _14522_ (.A(_08492_),
    .ZN(_08510_));
 INV_X1 _14523_ (.A(_07379_),
    .ZN(_07386_));
 INV_X1 _14524_ (.A(_07412_),
    .ZN(_07388_));
 INV_X1 _14525_ (.A(_07416_),
    .ZN(_07426_));
 INV_X1 _14526_ (.A(_07441_),
    .ZN(_07436_));
 INV_X1 _14527_ (.A(_07447_),
    .ZN(_07428_));
 INV_X1 _14528_ (.A(_07456_),
    .ZN(_07466_));
 INV_X1 _14529_ (.A(_07510_),
    .ZN(_07520_));
 INV_X1 _14530_ (.A(_07514_),
    .ZN(_07468_));
 INV_X1 _14531_ (.A(_07545_),
    .ZN(_07541_));
 INV_X1 _14532_ (.A(_07557_),
    .ZN(_07566_));
 INV_X1 _14533_ (.A(_07561_),
    .ZN(_07522_));
 INV_X1 _14534_ (.A(_07596_),
    .ZN(_07592_));
 INV_X1 _14535_ (.A(_07605_),
    .ZN(_07568_));
 INV_X1 _14536_ (.A(_07612_),
    .ZN(_07623_));
 INV_X1 _14537_ (.A(_07645_),
    .ZN(_07639_));
 INV_X1 _14538_ (.A(_07740_),
    .ZN(_07734_));
 INV_X1 _14539_ (.A(_07783_),
    .ZN(_07777_));
 INV_X1 _14540_ (.A(_07822_),
    .ZN(_07816_));
 INV_X1 _14541_ (.A(_07931_),
    .ZN(_07935_));
 INV_X1 _14542_ (.A(_07954_),
    .ZN(_07963_));
 INV_X1 _14543_ (.A(_07987_),
    .ZN(_07981_));
 INV_X1 _14544_ (.A(_08007_),
    .ZN(_08010_));
 INV_X1 _14545_ (.A(_08041_),
    .ZN(_08050_));
 INV_X1 _14546_ (.A(_08047_),
    .ZN(_07973_));
 INV_X1 _14547_ (.A(_08067_),
    .ZN(_08070_));
 INV_X1 _14548_ (.A(_08106_),
    .ZN(_08113_));
 INV_X1 _14549_ (.A(_08128_),
    .ZN(_09612_));
 INV_X1 _14550_ (.A(_08169_),
    .ZN(_08177_));
 INV_X1 _14551_ (.A(_08122_),
    .ZN(_08119_));
 INV_X1 _14552_ (.A(_08192_),
    .ZN(_09623_));
 INV_X1 _14553_ (.A(_08231_),
    .ZN(_08239_));
 INV_X1 _14554_ (.A(_08185_),
    .ZN(_08182_));
 INV_X1 _14555_ (.A(_08300_),
    .ZN(_08262_));
 INV_X1 _14556_ (.A(_08334_),
    .ZN(_08338_));
 INV_X1 _14557_ (.A(_08350_),
    .ZN(_08309_));
 INV_X1 _14558_ (.A(_08356_),
    .ZN(_08360_));
 INV_X1 _14559_ (.A(_08391_),
    .ZN(_08359_));
 INV_X1 _14560_ (.A(_08388_),
    .ZN(_08384_));
 INV_X1 _14561_ (.A(_08495_),
    .ZN(_08475_));
 INV_X1 _14562_ (.A(_07400_),
    .ZN(_07418_));
 INV_X1 _14563_ (.A(_07390_),
    .ZN(_07406_));
 INV_X1 _14564_ (.A(_07425_),
    .ZN(_07445_));
 INV_X2 _14565_ (.A(_00025_),
    .ZN(_05126_));
 CLKBUF_X3 _14566_ (.A(_05126_),
    .Z(_05127_));
 NOR2_X1 _14567_ (.A1(_05127_),
    .A2(_04980_),
    .ZN(_09397_));
 INV_X1 _14568_ (.A(_07452_),
    .ZN(_07462_));
 NOR2_X1 _14569_ (.A1(_05127_),
    .A2(_04971_),
    .ZN(_09404_));
 INV_X1 _14570_ (.A(_07502_),
    .ZN(_09420_));
 INV_X1 _14571_ (.A(_07497_),
    .ZN(_07543_));
 NOR2_X1 _14572_ (.A1(_05127_),
    .A2(_04962_),
    .ZN(_09423_));
 NOR2_X1 _14573_ (.A1(_05127_),
    .A2(_04953_),
    .ZN(_09435_));
 INV_X1 _14574_ (.A(_07581_),
    .ZN(_09445_));
 INV_X1 _14575_ (.A(_07540_),
    .ZN(_07583_));
 NOR2_X1 _14576_ (.A1(_05127_),
    .A2(_04944_),
    .ZN(_09448_));
 INV_X1 _14577_ (.A(_07625_),
    .ZN(_09458_));
 INV_X1 _14578_ (.A(_07590_),
    .ZN(_07631_));
 NOR2_X1 _14579_ (.A1(_05127_),
    .A2(_04934_),
    .ZN(_09463_));
 INV_X1 _14580_ (.A(_07662_),
    .ZN(_07673_));
 INV_X1 _14581_ (.A(_07637_),
    .ZN(_07682_));
 NOR2_X1 _14582_ (.A1(_05127_),
    .A2(_04916_),
    .ZN(_09477_));
 INV_X1 _14583_ (.A(_07696_),
    .ZN(_07737_));
 INV_X1 _14584_ (.A(_07713_),
    .ZN(_07720_));
 INV_X1 _14585_ (.A(_07689_),
    .ZN(_07729_));
 INV_X1 _14586_ (.A(_07714_),
    .ZN(_07739_));
 INV_X1 _14587_ (.A(_07745_),
    .ZN(_09487_));
 NOR2_X1 _14588_ (.A1(_05127_),
    .A2(_04906_),
    .ZN(_09492_));
 INV_X1 _14589_ (.A(_07785_),
    .ZN(_07787_));
 INV_X1 _14590_ (.A(_07756_),
    .ZN(_07762_));
 INV_X1 _14591_ (.A(_07736_),
    .ZN(_07771_));
 INV_X1 _14592_ (.A(_07757_),
    .ZN(_07782_));
 NOR2_X1 _14593_ (.A1(_05127_),
    .A2(_04894_),
    .ZN(_09505_));
 INV_X1 _14594_ (.A(_07854_),
    .ZN(_07824_));
 INV_X1 _14595_ (.A(_07795_),
    .ZN(_07801_));
 INV_X1 _14596_ (.A(_07814_),
    .ZN(_07810_));
 INV_X1 _14597_ (.A(_07796_),
    .ZN(_07821_));
 NOR2_X1 _14598_ (.A1(_05127_),
    .A2(net437),
    .ZN(_09515_));
 INV_X1 _14599_ (.A(_07836_),
    .ZN(_09526_));
 INV_X1 _14600_ (.A(_07818_),
    .ZN(_07842_));
 INV_X1 _14601_ (.A(_07837_),
    .ZN(_07847_));
 NOR2_X1 _14602_ (.A1(_05126_),
    .A2(_04864_),
    .ZN(_09532_));
 INV_X1 _14603_ (.A(_07859_),
    .ZN(_09542_));
 NOR2_X1 _14604_ (.A1(_05126_),
    .A2(_04849_),
    .ZN(_09547_));
 INV_X1 _14605_ (.A(_07880_),
    .ZN(_07887_));
 INV_X1 _14606_ (.A(_07881_),
    .ZN(_07890_));
 NOR2_X1 _14607_ (.A1(_05126_),
    .A2(_04822_),
    .ZN(_09578_));
 OR2_X2 _14608_ (.A1(_04850_),
    .A2(_04990_),
    .ZN(_08019_));
 INV_X1 _14609_ (.A(_07938_),
    .ZN(_07957_));
 INV_X1 _14610_ (.A(_07966_),
    .ZN(_08044_));
 INV_X1 _14611_ (.A(_07998_),
    .ZN(_08014_));
 INV_X1 _14612_ (.A(_08061_),
    .ZN(_08057_));
 INV_X1 _14613_ (.A(_08053_),
    .ZN(_08109_));
 INV_X1 _14614_ (.A(_08023_),
    .ZN(_08074_));
 INV_X1 _14615_ (.A(_08116_),
    .ZN(_08171_));
 INV_X1 _14616_ (.A(_08081_),
    .ZN(_08131_));
 INV_X1 _14617_ (.A(_08093_),
    .ZN(_08149_));
 INV_X1 _14618_ (.A(_08179_),
    .ZN(_08235_));
 INV_X1 _14619_ (.A(_08183_),
    .ZN(_08207_));
 INV_X1 _14620_ (.A(_08139_),
    .ZN(_08195_));
 INV_X1 _14621_ (.A(_08156_),
    .ZN(_08216_));
 INV_X1 _14622_ (.A(_08247_),
    .ZN(_08243_));
 INV_X1 _14623_ (.A(_08202_),
    .ZN(_08253_));
 INV_X1 _14624_ (.A(_08222_),
    .ZN(_08273_));
 INV_X1 _14625_ (.A(_08264_),
    .ZN(_09643_));
 INV_X1 _14626_ (.A(_08260_),
    .ZN(_08299_));
 INV_X1 _14627_ (.A(_08291_),
    .ZN(_09652_));
 INV_X1 _14628_ (.A(_08347_),
    .ZN(_08342_));
 INV_X1 _14629_ (.A(_08311_),
    .ZN(_09657_));
 INV_X1 _14630_ (.A(_08307_),
    .ZN(_08349_));
 BUF_X4 _14631_ (.A(_05122_),
    .Z(_05128_));
 NOR2_X1 _14632_ (.A1(_05128_),
    .A2(_05082_),
    .ZN(_08354_));
 INV_X1 _14633_ (.A(_08327_),
    .ZN(_08371_));
 INV_X1 _14634_ (.A(_08341_),
    .ZN(_09665_));
 INV_X1 _14635_ (.A(_08362_),
    .ZN(_09670_));
 INV_X1 _14636_ (.A(_08407_),
    .ZN(_08402_));
 INV_X1 _14637_ (.A(_08378_),
    .ZN(_08412_));
 INV_X1 _14638_ (.A(_08387_),
    .ZN(_09674_));
 INV_X1 _14639_ (.A(_09682_),
    .ZN(_09685_));
 INV_X1 _14640_ (.A(_08423_),
    .ZN(_08435_));
 INV_X1 _14641_ (.A(_08419_),
    .ZN(_08431_));
 INV_X1 _14642_ (.A(_09679_),
    .ZN(_09691_));
 INV_X1 _14643_ (.A(_08446_),
    .ZN(_08452_));
 INV_X1 _14644_ (.A(_09699_),
    .ZN(_09700_));
 INV_X1 _14645_ (.A(_08443_),
    .ZN(_08464_));
 INV_X1 _14646_ (.A(_09704_),
    .ZN(_08489_));
 INV_X1 _14647_ (.A(_08473_),
    .ZN(_09713_));
 INV_X1 _14648_ (.A(_08472_),
    .ZN(_08485_));
 INV_X1 _14649_ (.A(_08476_),
    .ZN(_08483_));
 INV_X1 _14650_ (.A(_08477_),
    .ZN(_08487_));
 INV_X1 _14651_ (.A(_09720_),
    .ZN(_09730_));
 INV_X1 _14652_ (.A(_08517_),
    .ZN(_08523_));
 NOR2_X1 _14653_ (.A1(_05128_),
    .A2(_05028_),
    .ZN(_09748_));
 INV_X1 _14654_ (.A(_08559_),
    .ZN(_08557_));
 NOR4_X1 _14655_ (.A1(_08599_),
    .A2(_08604_),
    .A3(_08609_),
    .A4(_08559_),
    .ZN(_05129_));
 NOR4_X1 _14656_ (.A1(_08614_),
    .A2(_08619_),
    .A3(_08624_),
    .A4(_08629_),
    .ZN(_05130_));
 NOR4_X1 _14657_ (.A1(_08561_),
    .A2(_08553_),
    .A3(_08569_),
    .A4(_08594_),
    .ZN(_05131_));
 NOR4_X1 _14658_ (.A1(_08574_),
    .A2(_08579_),
    .A3(_08584_),
    .A4(_08589_),
    .ZN(_05132_));
 NAND4_X1 _14659_ (.A1(_05129_),
    .A2(_05130_),
    .A3(_05131_),
    .A4(_05132_),
    .ZN(_08562_));
 INV_X1 _14660_ (.A(_08640_),
    .ZN(_08638_));
 NOR4_X1 _14661_ (.A1(_08680_),
    .A2(_08685_),
    .A3(_08690_),
    .A4(_08640_),
    .ZN(_05133_));
 NOR4_X1 _14662_ (.A1(_08695_),
    .A2(_08700_),
    .A3(_08705_),
    .A4(_08710_),
    .ZN(_05134_));
 NOR4_X1 _14663_ (.A1(_08642_),
    .A2(_08634_),
    .A3(_08650_),
    .A4(_08675_),
    .ZN(_05135_));
 NOR4_X1 _14664_ (.A1(_08655_),
    .A2(_08660_),
    .A3(_08665_),
    .A4(_08670_),
    .ZN(_05136_));
 NAND4_X1 _14665_ (.A1(_05133_),
    .A2(_05134_),
    .A3(_05135_),
    .A4(_05136_),
    .ZN(_08643_));
 MUX2_X1 _14666_ (.A(_08722_),
    .B(_01167_),
    .S(_01428_),
    .Z(_08731_));
 INV_X2 _14667_ (.A(_01429_),
    .ZN(_08734_));
 NAND3_X1 _14668_ (.A1(_01168_),
    .A2(_01180_),
    .A3(_01208_),
    .ZN(_08744_));
 AOI21_X2 _14669_ (.A(_01425_),
    .B1(_01429_),
    .B2(net3),
    .ZN(_08747_));
 NOR2_X1 _14670_ (.A1(_01228_),
    .A2(_01305_),
    .ZN(_08765_));
 NAND2_X1 _14671_ (.A1(_01419_),
    .A2(_08747_),
    .ZN(_05137_));
 NAND2_X1 _14672_ (.A1(_05137_),
    .A2(_01432_),
    .ZN(_08768_));
 INV_X1 _14673_ (.A(_01353_),
    .ZN(_08778_));
 INV_X1 _14674_ (.A(_01436_),
    .ZN(_08781_));
 INV_X1 _14675_ (.A(_01476_),
    .ZN(_08801_));
 AOI211_X4 _14676_ (.A(_01102_),
    .B(_01249_),
    .C1(_01105_),
    .C2(_01107_),
    .ZN(_08816_));
 MUX2_X1 _14677_ (.A(_01476_),
    .B(_01464_),
    .S(_01309_),
    .Z(_05138_));
 INV_X1 _14678_ (.A(_05138_),
    .ZN(_08823_));
 INV_X1 _14679_ (.A(_03366_),
    .ZN(_09150_));
 XOR2_X1 _14680_ (.A(_09296_),
    .B(_09287_),
    .Z(_05139_));
 MUX2_X1 _14681_ (.A(_04768_),
    .B(_05139_),
    .S(_04724_),
    .Z(_09330_));
 MUX2_X1 _14682_ (.A(_09285_),
    .B(_09288_),
    .S(_04724_),
    .Z(_05140_));
 INV_X1 _14683_ (.A(_05140_),
    .ZN(_07368_));
 INV_X1 _14684_ (.A(_09336_),
    .ZN(_07369_));
 INV_X1 _14685_ (.A(_07424_),
    .ZN(_07419_));
 NOR2_X1 _14686_ (.A1(_05128_),
    .A2(_05001_),
    .ZN(_09398_));
 INV_X1 _14687_ (.A(_07501_),
    .ZN(_09401_));
 NOR2_X1 _14688_ (.A1(_05128_),
    .A2(_04980_),
    .ZN(_09405_));
 INV_X1 _14689_ (.A(_07506_),
    .ZN(_07517_));
 NOR2_X1 _14690_ (.A1(_05128_),
    .A2(_04971_),
    .ZN(_09424_));
 NOR2_X1 _14691_ (.A1(_05128_),
    .A2(net438),
    .ZN(_09436_));
 INV_X1 _14692_ (.A(_07588_),
    .ZN(_07584_));
 NOR2_X1 _14693_ (.A1(_05128_),
    .A2(_04953_),
    .ZN(_09449_));
 INV_X1 _14694_ (.A(_07635_),
    .ZN(_07632_));
 INV_X1 _14695_ (.A(_07700_),
    .ZN(_07697_));
 NOR2_X1 _14696_ (.A1(_05128_),
    .A2(_04944_),
    .ZN(_09464_));
 INV_X1 _14697_ (.A(_07667_),
    .ZN(_07674_));
 INV_X1 _14698_ (.A(_07686_),
    .ZN(_07683_));
 INV_X1 _14699_ (.A(_07744_),
    .ZN(_09472_));
 NOR2_X1 _14700_ (.A1(_05128_),
    .A2(_04934_),
    .ZN(_09478_));
 INV_X1 _14701_ (.A(_07733_),
    .ZN(_07730_));
 NOR2_X1 _14702_ (.A1(_05128_),
    .A2(_04916_),
    .ZN(_09493_));
 INV_X1 _14703_ (.A(_07775_),
    .ZN(_07772_));
 NOR2_X1 _14704_ (.A1(_05122_),
    .A2(_04906_),
    .ZN(_09506_));
 INV_X1 _14705_ (.A(_07779_),
    .ZN(_07811_));
 INV_X1 _14706_ (.A(_07786_),
    .ZN(_09512_));
 NOR2_X1 _14707_ (.A1(_05122_),
    .A2(_04894_),
    .ZN(_09516_));
 INV_X1 _14708_ (.A(_07858_),
    .ZN(_09529_));
 NOR2_X1 _14709_ (.A1(_05122_),
    .A2(net437),
    .ZN(_09533_));
 INV_X1 _14710_ (.A(_07855_),
    .ZN(_09541_));
 NOR2_X1 _14711_ (.A1(_05122_),
    .A2(_04864_),
    .ZN(_09548_));
 INV_X1 _14712_ (.A(_07903_),
    .ZN(_07900_));
 INV_X1 _14713_ (.A(_07910_),
    .ZN(_09575_));
 NOR2_X1 _14714_ (.A1(_05122_),
    .A2(_04849_),
    .ZN(_09579_));
 INV_X1 _14715_ (.A(_07965_),
    .ZN(_07958_));
 INV_X1 _14716_ (.A(_08052_),
    .ZN(_08045_));
 INV_X1 _14717_ (.A(_08022_),
    .ZN(_08025_));
 INV_X1 _14718_ (.A(_08115_),
    .ZN(_08110_));
 INV_X1 _14719_ (.A(_08012_),
    .ZN(_09604_));
 INV_X1 _14720_ (.A(_08080_),
    .ZN(_08083_));
 INV_X1 _14721_ (.A(_08175_),
    .ZN(_08172_));
 INV_X1 _14722_ (.A(_08072_),
    .ZN(_09610_));
 INV_X1 _14723_ (.A(_08188_),
    .ZN(_08146_));
 INV_X1 _14724_ (.A(_08154_),
    .ZN(_08150_));
 INV_X1 _14725_ (.A(_08241_),
    .ZN(_08236_));
 INV_X1 _14726_ (.A(_08189_),
    .ZN(_08208_));
 INV_X1 _14727_ (.A(_08201_),
    .ZN(_08204_));
 INV_X1 _14728_ (.A(_08250_),
    .ZN(_08209_));
 INV_X1 _14729_ (.A(_08220_),
    .ZN(_08217_));
 INV_X1 _14730_ (.A(_08251_),
    .ZN(_08265_));
 INV_X1 _14731_ (.A(_08277_),
    .ZN(_08274_));
 INV_X1 _14732_ (.A(_08290_),
    .ZN(_09638_));
 INV_X1 _14733_ (.A(_08263_),
    .ZN(_09646_));
 INV_X1 _14734_ (.A(_08324_),
    .ZN(_08321_));
 INV_X1 _14735_ (.A(_08340_),
    .ZN(_09653_));
 INV_X1 _14736_ (.A(_08310_),
    .ZN(_09660_));
 INV_X1 _14737_ (.A(_08375_),
    .ZN(_08372_));
 INV_X1 _14738_ (.A(_08386_),
    .ZN(_09666_));
 INV_X1 _14739_ (.A(_09676_),
    .ZN(_09669_));
 INV_X1 _14740_ (.A(_08361_),
    .ZN(_09671_));
 INV_X1 _14741_ (.A(_08416_),
    .ZN(_08413_));
 INV_X1 _14742_ (.A(_09678_),
    .ZN(_09675_));
 INV_X1 _14743_ (.A(_09693_),
    .ZN(_09681_));
 INV_X1 _14744_ (.A(_08401_),
    .ZN(_09683_));
 INV_X1 _14745_ (.A(_08439_),
    .ZN(_08436_));
 INV_X1 _14746_ (.A(_08400_),
    .ZN(_09687_));
 INV_X1 _14747_ (.A(_09695_),
    .ZN(_09692_));
 INV_X1 _14748_ (.A(_08450_),
    .ZN(_08454_));
 INV_X1 _14749_ (.A(_08468_),
    .ZN(_08465_));
 INV_X1 _14750_ (.A(_09721_),
    .ZN(_08490_));
 INV_X1 _14751_ (.A(_08451_),
    .ZN(_09709_));
 INV_X1 _14752_ (.A(_09707_),
    .ZN(_09719_));
 INV_X1 _14753_ (.A(_09722_),
    .ZN(_09731_));
 INV_X1 _14754_ (.A(_08543_),
    .ZN(_09746_));
 NOR2_X1 _14755_ (.A1(_05126_),
    .A2(_05055_),
    .ZN(_09749_));
 INV_X1 _14756_ (.A(_09400_),
    .ZN(_07494_));
 INV_X1 _14757_ (.A(_09412_),
    .ZN(_07477_));
 INV_X1 _14758_ (.A(_09426_),
    .ZN(_07571_));
 INV_X1 _14759_ (.A(_09438_),
    .ZN(_07614_));
 INV_X1 _14760_ (.A(_09451_),
    .ZN(_07664_));
 INV_X1 _14761_ (.A(_09459_),
    .ZN(_07693_));
 INV_X1 _14762_ (.A(_09520_),
    .ZN(_07834_));
 INV_X1 _14763_ (.A(_09559_),
    .ZN(_07904_));
 INV_X1 _14764_ (.A(_09605_),
    .ZN(_08123_));
 INV_X1 _14765_ (.A(_09611_),
    .ZN(_08186_));
 INV_X1 _14766_ (.A(_09622_),
    .ZN(_08248_));
 INV_X1 _14767_ (.A(_09708_),
    .ZN(_08491_));
 INV_X1 _14768_ (.A(_09476_),
    .ZN(_07711_));
 INV_X1 _14769_ (.A(_09491_),
    .ZN(_07754_));
 INV_X1 _14770_ (.A(_09504_),
    .ZN(_07793_));
 INV_X1 _14771_ (.A(_07912_),
    .ZN(_07909_));
 INV_X1 _14772_ (.A(_09517_),
    .ZN(_07856_));
 INV_X1 _14773_ (.A(_08522_),
    .ZN(_08518_));
 INV_X1 _14774_ (.A(_09667_),
    .ZN(_09668_));
 INV_X1 _14775_ (.A(_09677_),
    .ZN(_09680_));
 INV_X1 _14776_ (.A(_09694_),
    .ZN(_09697_));
 INV_X1 _14777_ (.A(_09710_),
    .ZN(_08474_));
 INV_X1 _14778_ (.A(_09732_),
    .ZN(_09737_));
 NAND2_X1 _14779_ (.A1(\butterfly_in_group[0] ),
    .A2(_04792_),
    .ZN(_05141_));
 INV_X1 _14780_ (.A(_04589_),
    .ZN(_05142_));
 OR2_X1 _14781_ (.A1(_04668_),
    .A2(_04693_),
    .ZN(_05143_));
 NOR3_X1 _14782_ (.A1(_05142_),
    .A2(net22),
    .A3(_05143_),
    .ZN(_05144_));
 NOR2_X1 _14783_ (.A1(_04718_),
    .A2(_04573_),
    .ZN(_05145_));
 NAND2_X1 _14784_ (.A1(_04515_),
    .A2(_05145_),
    .ZN(_05146_));
 XNOR2_X1 _14785_ (.A(_04516_),
    .B(_05146_),
    .ZN(_05147_));
 AND2_X1 _14786_ (.A1(_04653_),
    .A2(_04654_),
    .ZN(_05148_));
 AND2_X1 _14787_ (.A1(_04655_),
    .A2(_04667_),
    .ZN(_05149_));
 OAI21_X1 _14788_ (.A(_04635_),
    .B1(_04740_),
    .B2(_04734_),
    .ZN(_05150_));
 AOI21_X2 _14789_ (.A(_09298_),
    .B1(_05150_),
    .B2(_04646_),
    .ZN(_05151_));
 OR3_X2 _14790_ (.A1(_04633_),
    .A2(_04634_),
    .A3(_05151_),
    .ZN(_05152_));
 NAND3_X1 _14791_ (.A1(_09279_),
    .A2(_04521_),
    .A3(net34),
    .ZN(_05153_));
 INV_X1 _14792_ (.A(_04664_),
    .ZN(_05154_));
 OAI21_X1 _14793_ (.A(_05154_),
    .B1(_04579_),
    .B2(_04580_),
    .ZN(_05155_));
 NAND2_X1 _14794_ (.A1(_05153_),
    .A2(_05155_),
    .ZN(_05156_));
 NOR2_X1 _14795_ (.A1(_04718_),
    .A2(_04663_),
    .ZN(_05157_));
 OR2_X1 _14796_ (.A1(_05156_),
    .A2(_05157_),
    .ZN(_05158_));
 OAI211_X2 _14797_ (.A(_05148_),
    .B(_05149_),
    .C1(_05152_),
    .C2(_05158_),
    .ZN(_05159_));
 NAND3_X1 _14798_ (.A1(_04685_),
    .A2(_04688_),
    .A3(_04692_),
    .ZN(_05160_));
 NAND2_X1 _14799_ (.A1(_04653_),
    .A2(_04654_),
    .ZN(_05161_));
 AOI21_X1 _14800_ (.A(_05161_),
    .B1(_05149_),
    .B2(_05152_),
    .ZN(_05162_));
 AND3_X1 _14801_ (.A1(_05161_),
    .A2(_05149_),
    .A3(_05152_),
    .ZN(_05163_));
 OAI221_X2 _14802_ (.A(_05147_),
    .B1(_05159_),
    .B2(_05160_),
    .C1(_05162_),
    .C2(_05163_),
    .ZN(_05164_));
 NAND2_X1 _14803_ (.A1(_04705_),
    .A2(_04706_),
    .ZN(_05165_));
 AND3_X1 _14804_ (.A1(_04611_),
    .A2(_04694_),
    .A3(_05165_),
    .ZN(_05166_));
 NOR3_X1 _14805_ (.A1(_05144_),
    .A2(_05164_),
    .A3(_05166_),
    .ZN(_05167_));
 XNOR2_X1 _14806_ (.A(_04681_),
    .B(_04684_),
    .ZN(_05168_));
 NOR2_X1 _14807_ (.A1(_05168_),
    .A2(net24),
    .ZN(_05169_));
 OAI21_X2 _14808_ (.A(_04717_),
    .B1(_05167_),
    .B2(_05169_),
    .ZN(_05170_));
 NAND3_X1 _14809_ (.A1(_04611_),
    .A2(_04694_),
    .A3(_05165_),
    .ZN(_05171_));
 OR4_X2 _14810_ (.A1(_04717_),
    .A2(_05144_),
    .A3(_05164_),
    .A4(_05171_),
    .ZN(_05172_));
 INV_X1 _14811_ (.A(_09288_),
    .ZN(_05173_));
 MUX2_X1 _14812_ (.A(\butterfly_count[1] ),
    .B(_05173_),
    .S(_04723_),
    .Z(_05174_));
 BUF_X1 _14813_ (.A(_09332_),
    .Z(_05175_));
 NAND2_X1 _14814_ (.A1(_09320_),
    .A2(_09324_),
    .ZN(_05176_));
 NAND3_X1 _14815_ (.A1(_09316_),
    .A2(_09312_),
    .A3(_09328_),
    .ZN(_05177_));
 NOR2_X2 _14816_ (.A1(_05177_),
    .A2(_05176_),
    .ZN(_05178_));
 NAND3_X1 _14817_ (.A1(_05175_),
    .A2(_07363_),
    .A3(_05178_),
    .ZN(_05179_));
 OR2_X1 _14818_ (.A1(_05174_),
    .A2(_05179_),
    .ZN(_05180_));
 AOI21_X1 _14819_ (.A(_09319_),
    .B1(_09320_),
    .B2(_09323_),
    .ZN(_05181_));
 INV_X1 _14820_ (.A(_09331_),
    .ZN(_05182_));
 NAND2_X1 _14821_ (.A1(_09334_),
    .A2(_05175_),
    .ZN(_05183_));
 OAI21_X1 _14822_ (.A(_05182_),
    .B1(_05183_),
    .B2(_09338_),
    .ZN(_05184_));
 AOI21_X1 _14823_ (.A(_09327_),
    .B1(_05184_),
    .B2(_09328_),
    .ZN(_05185_));
 OAI21_X1 _14824_ (.A(_05181_),
    .B1(_05185_),
    .B2(_05176_),
    .ZN(_05186_));
 AOI21_X1 _14825_ (.A(_09315_),
    .B1(_05186_),
    .B2(_09316_),
    .ZN(_05187_));
 INV_X1 _14826_ (.A(_05187_),
    .ZN(_05188_));
 AOI21_X1 _14827_ (.A(_09311_),
    .B1(_05188_),
    .B2(_09312_),
    .ZN(_05189_));
 AOI22_X2 _14828_ (.A1(_05170_),
    .A2(_05172_),
    .B1(_05180_),
    .B2(_05189_),
    .ZN(_05190_));
 NAND2_X1 _14829_ (.A1(_04688_),
    .A2(_04692_),
    .ZN(_05191_));
 OAI21_X1 _14830_ (.A(_05168_),
    .B1(_05191_),
    .B2(_05159_),
    .ZN(_05192_));
 NAND3_X1 _14831_ (.A1(_04576_),
    .A2(_04577_),
    .A3(_04686_),
    .ZN(_05193_));
 XOR2_X1 _14832_ (.A(_04507_),
    .B(_05193_),
    .Z(_05194_));
 NAND2_X1 _14833_ (.A1(_04576_),
    .A2(_05145_),
    .ZN(_05195_));
 XNOR2_X2 _14834_ (.A(_04502_),
    .B(_05195_),
    .ZN(_05196_));
 NOR3_X1 _14835_ (.A1(_04648_),
    .A2(_05143_),
    .A3(_05196_),
    .ZN(_05197_));
 OAI21_X1 _14836_ (.A(_04589_),
    .B1(_04593_),
    .B2(_04596_),
    .ZN(_05198_));
 OR2_X2 _14837_ (.A1(_04633_),
    .A2(_04634_),
    .ZN(_05199_));
 NOR2_X1 _14838_ (.A1(_04734_),
    .A2(_04740_),
    .ZN(_05200_));
 AND3_X1 _14839_ (.A1(_05200_),
    .A2(_05153_),
    .A3(_05155_),
    .ZN(_05201_));
 OAI21_X1 _14840_ (.A(_04646_),
    .B1(_09301_),
    .B2(_05201_),
    .ZN(_05202_));
 INV_X1 _14841_ (.A(_09298_),
    .ZN(_05203_));
 AOI21_X2 _14842_ (.A(_05199_),
    .B1(_05202_),
    .B2(_05203_),
    .ZN(_05204_));
 NOR3_X1 _14843_ (.A1(_05198_),
    .A2(_05143_),
    .A3(_05204_),
    .ZN(_05205_));
 OAI221_X1 _14844_ (.A(_05192_),
    .B1(_05194_),
    .B2(_05197_),
    .C1(_05205_),
    .C2(_04575_),
    .ZN(_05206_));
 NOR2_X1 _14845_ (.A1(_04597_),
    .A2(_04610_),
    .ZN(_05207_));
 NOR3_X1 _14846_ (.A1(_04648_),
    .A2(_04668_),
    .A3(_05160_),
    .ZN(_05208_));
 NAND3_X1 _14847_ (.A1(_05207_),
    .A2(_04672_),
    .A3(_05208_),
    .ZN(_05209_));
 XOR2_X1 _14848_ (.A(_04368_),
    .B(_04570_),
    .Z(_05210_));
 OAI21_X1 _14849_ (.A(_05210_),
    .B1(_04672_),
    .B2(_05208_),
    .ZN(_05211_));
 AND2_X1 _14850_ (.A1(_05209_),
    .A2(_05211_),
    .ZN(_05212_));
 NOR3_X2 _14851_ (.A1(_04718_),
    .A2(_04573_),
    .A3(_04687_),
    .ZN(_05213_));
 XNOR2_X2 _14852_ (.A(_04690_),
    .B(_05213_),
    .ZN(_05214_));
 XOR2_X2 _14853_ (.A(_04686_),
    .B(_04687_),
    .Z(_05215_));
 NOR2_X1 _14854_ (.A1(_04668_),
    .A2(_05215_),
    .ZN(_05216_));
 AND2_X1 _14855_ (.A1(_05203_),
    .A2(_05202_),
    .ZN(_05217_));
 OAI221_X1 _14856_ (.A(_05216_),
    .B1(_04693_),
    .B2(net22),
    .C1(_05199_),
    .C2(_05217_),
    .ZN(_05218_));
 AND2_X1 _14857_ (.A1(_05214_),
    .A2(_05218_),
    .ZN(_05219_));
 NOR4_X1 _14858_ (.A1(_04668_),
    .A2(_04672_),
    .A3(_05215_),
    .A4(_05214_),
    .ZN(_05220_));
 OAI21_X1 _14859_ (.A(_05220_),
    .B1(_05217_),
    .B2(_05199_),
    .ZN(_05221_));
 NAND4_X2 _14860_ (.A1(_05178_),
    .A2(_09334_),
    .A3(_09337_),
    .A4(_05175_),
    .ZN(_05222_));
 NOR3_X1 _14861_ (.A1(_04718_),
    .A2(_04656_),
    .A3(_04659_),
    .ZN(_05223_));
 XOR2_X1 _14862_ (.A(_04658_),
    .B(_05223_),
    .Z(_05224_));
 NAND2_X1 _14863_ (.A1(_04686_),
    .A2(_04513_),
    .ZN(_05225_));
 XNOR2_X1 _14864_ (.A(_04462_),
    .B(_05225_),
    .ZN(_05226_));
 AND4_X4 _14865_ (.A1(_05222_),
    .A2(_04608_),
    .A3(_05224_),
    .A4(_05226_),
    .ZN(_05227_));
 NAND3_X4 _14866_ (.A1(_04714_),
    .A2(_05221_),
    .A3(_05227_),
    .ZN(_05228_));
 NOR4_X4 _14867_ (.A1(_05228_),
    .A2(_05212_),
    .A3(_05219_),
    .A4(_05206_),
    .ZN(_05229_));
 AND4_X1 _14868_ (.A1(_04611_),
    .A2(_04694_),
    .A3(_04698_),
    .A4(_04722_),
    .ZN(_05230_));
 NOR4_X1 _14869_ (.A1(_04597_),
    .A2(_05230_),
    .A3(_05143_),
    .A4(_05204_),
    .ZN(_05231_));
 NOR2_X1 _14870_ (.A1(_04668_),
    .A2(_04693_),
    .ZN(_05232_));
 AND2_X1 _14871_ (.A1(_05165_),
    .A2(_04717_),
    .ZN(_05233_));
 OR2_X1 _14872_ (.A1(_05152_),
    .A2(_05156_),
    .ZN(_05234_));
 AND4_X1 _14873_ (.A1(_04611_),
    .A2(_05232_),
    .A3(_05233_),
    .A4(_05234_),
    .ZN(_05235_));
 AOI21_X1 _14874_ (.A(_04716_),
    .B1(net24),
    .B2(_05235_),
    .ZN(_05236_));
 AND3_X1 _14875_ (.A1(_04716_),
    .A2(_04723_),
    .A3(_05235_),
    .ZN(_05237_));
 NOR3_X1 _14876_ (.A1(_05231_),
    .A2(_05236_),
    .A3(_05237_),
    .ZN(_05238_));
 NAND2_X1 _14877_ (.A1(_04565_),
    .A2(net37),
    .ZN(_05239_));
 XNOR2_X2 _14878_ (.A(_05239_),
    .B(_04659_),
    .ZN(_05240_));
 AND2_X1 _14879_ (.A1(_04629_),
    .A2(_04632_),
    .ZN(_05241_));
 AOI21_X1 _14880_ (.A(_05156_),
    .B1(_05241_),
    .B2(_02573_),
    .ZN(_05242_));
 NAND3_X1 _14881_ (.A1(_05199_),
    .A2(_05151_),
    .A3(_05242_),
    .ZN(_05243_));
 NAND2_X1 _14882_ (.A1(_05240_),
    .A2(_05243_),
    .ZN(_05244_));
 XOR2_X1 _14883_ (.A(_05199_),
    .B(_05151_),
    .Z(_05245_));
 OAI22_X1 _14884_ (.A1(_05152_),
    .A2(_05217_),
    .B1(_05242_),
    .B2(_05245_),
    .ZN(_05246_));
 OAI21_X1 _14885_ (.A(_05244_),
    .B1(_05246_),
    .B2(_05240_),
    .ZN(_05247_));
 AOI21_X1 _14886_ (.A(_04648_),
    .B1(_05241_),
    .B2(_02573_),
    .ZN(_05248_));
 XOR2_X1 _14887_ (.A(_05156_),
    .B(_05248_),
    .Z(_05249_));
 OR2_X1 _14888_ (.A1(_04694_),
    .A2(_05249_),
    .ZN(_05250_));
 OAI21_X1 _14889_ (.A(_05216_),
    .B1(_05217_),
    .B2(_05199_),
    .ZN(_05251_));
 XNOR2_X1 _14890_ (.A(_05214_),
    .B(_05251_),
    .ZN(_05252_));
 OR2_X1 _14891_ (.A1(_05156_),
    .A2(_05240_),
    .ZN(_05253_));
 OAI33_X1 _14892_ (.A1(_05247_),
    .A2(_05250_),
    .A3(_05252_),
    .B1(_05253_),
    .B2(_05241_),
    .B3(_04724_),
    .ZN(_05254_));
 OR2_X1 _14893_ (.A1(net22),
    .A2(_04668_),
    .ZN(_05255_));
 NOR4_X1 _14894_ (.A1(_04597_),
    .A2(_04648_),
    .A3(_04668_),
    .A4(_04693_),
    .ZN(_05256_));
 XNOR2_X1 _14895_ (.A(_04609_),
    .B(_05256_),
    .ZN(_05257_));
 OR4_X1 _14896_ (.A1(_05255_),
    .A2(_04688_),
    .A3(_05230_),
    .A4(_05257_),
    .ZN(_05258_));
 NAND2_X1 _14897_ (.A1(_04609_),
    .A2(_04688_),
    .ZN(_05259_));
 NOR2_X1 _14898_ (.A1(_05255_),
    .A2(_05230_),
    .ZN(_05260_));
 OAI21_X1 _14899_ (.A(_05258_),
    .B1(_05259_),
    .B2(_05260_),
    .ZN(_05261_));
 AND4_X4 _14900_ (.A1(_05229_),
    .A2(_05238_),
    .A3(_05254_),
    .A4(_05261_),
    .ZN(_05262_));
 NAND2_X1 _14901_ (.A1(_05190_),
    .A2(_05262_),
    .ZN(_05263_));
 INV_X1 _14902_ (.A(\butterfly_count[0] ),
    .ZN(_05264_));
 NOR2_X1 _14903_ (.A1(net22),
    .A2(_04668_),
    .ZN(_05265_));
 NOR2_X1 _14904_ (.A1(_05145_),
    .A2(_04679_),
    .ZN(_05266_));
 NAND3_X1 _14905_ (.A1(_05265_),
    .A2(net24),
    .A3(_05266_),
    .ZN(_05267_));
 AND2_X1 _14906_ (.A1(_04675_),
    .A2(_05267_),
    .ZN(_05268_));
 NAND2_X1 _14907_ (.A1(_05265_),
    .A2(_04690_),
    .ZN(_05269_));
 OAI21_X1 _14908_ (.A(_04679_),
    .B1(_05230_),
    .B2(_05269_),
    .ZN(_05270_));
 NAND2_X1 _14909_ (.A1(_04686_),
    .A2(_05270_),
    .ZN(_05271_));
 NOR2_X1 _14910_ (.A1(_05143_),
    .A2(_05204_),
    .ZN(_05272_));
 AND3_X1 _14911_ (.A1(_04714_),
    .A2(_04716_),
    .A3(_04717_),
    .ZN(_05273_));
 AND4_X1 _14912_ (.A1(_04611_),
    .A2(_04698_),
    .A3(_05196_),
    .A4(_05273_),
    .ZN(_05274_));
 NAND3_X1 _14913_ (.A1(net24),
    .A2(_05272_),
    .A3(_05274_),
    .ZN(_05275_));
 NAND3_X1 _14914_ (.A1(_04611_),
    .A2(_04694_),
    .A3(_04722_),
    .ZN(_05276_));
 NAND2_X1 _14915_ (.A1(_04698_),
    .A2(_04721_),
    .ZN(_05277_));
 NAND2_X1 _14916_ (.A1(_05276_),
    .A2(_05277_),
    .ZN(_05278_));
 AOI21_X1 _14917_ (.A(_05196_),
    .B1(_05272_),
    .B2(_04724_),
    .ZN(_05279_));
 AND3_X1 _14918_ (.A1(_04723_),
    .A2(_05272_),
    .A3(_05196_),
    .ZN(_05280_));
 OAI21_X2 _14919_ (.A(_05278_),
    .B1(_05279_),
    .B2(_05280_),
    .ZN(_05281_));
 AOI22_X4 _14920_ (.A1(_05268_),
    .A2(_05271_),
    .B1(_05275_),
    .B2(_05281_),
    .ZN(_05282_));
 NAND2_X1 _14921_ (.A1(_05264_),
    .A2(_05282_),
    .ZN(_05283_));
 OAI21_X1 _14922_ (.A(_04779_),
    .B1(_05263_),
    .B2(_05283_),
    .ZN(_05284_));
 NAND3_X4 _14923_ (.A1(_05190_),
    .A2(_05262_),
    .A3(_05282_),
    .ZN(_05285_));
 AND2_X4 _14924_ (.A1(_09337_),
    .A2(_05285_),
    .ZN(_05286_));
 OAI21_X1 _14925_ (.A(_05141_),
    .B1(_05284_),
    .B2(_05286_),
    .ZN(_00058_));
 INV_X1 _14926_ (.A(_07371_),
    .ZN(_05287_));
 NAND3_X1 _14927_ (.A1(_05287_),
    .A2(_04779_),
    .A3(_05285_),
    .ZN(_05288_));
 NAND2_X1 _14928_ (.A1(_04778_),
    .A2(_05174_),
    .ZN(_05289_));
 INV_X1 _14929_ (.A(\butterfly_in_group[1] ),
    .ZN(_05290_));
 OAI221_X1 _14930_ (.A(_05288_),
    .B1(_05289_),
    .B2(_05285_),
    .C1(_04779_),
    .C2(_05290_),
    .ZN(_00059_));
 NAND2_X1 _14931_ (.A1(\butterfly_in_group[2] ),
    .A2(_04792_),
    .ZN(_05291_));
 NAND2_X1 _14932_ (.A1(_09330_),
    .A2(_05282_),
    .ZN(_05292_));
 OAI21_X1 _14933_ (.A(_04779_),
    .B1(_05263_),
    .B2(_05292_),
    .ZN(_05293_));
 XNOR2_X1 _14934_ (.A(_07370_),
    .B(_05175_),
    .ZN(_05294_));
 AND2_X2 _14935_ (.A1(_05285_),
    .A2(_05294_),
    .ZN(_05295_));
 OAI21_X1 _14936_ (.A(_05291_),
    .B1(_05293_),
    .B2(_05295_),
    .ZN(_00060_));
 MUX2_X1 _14937_ (.A(\group[0] ),
    .B(_05285_),
    .S(_04779_),
    .Z(_00319_));
 MUX2_X1 _14938_ (.A(\group[1] ),
    .B(net24),
    .S(_04778_),
    .Z(_00320_));
 MUX2_X1 _14939_ (.A(\group[2] ),
    .B(net37),
    .S(_04778_),
    .Z(_00321_));
 CLKBUF_X3 _14940_ (.A(_00030_),
    .Z(_05296_));
 NOR2_X4 _14941_ (.A1(_04794_),
    .A2(\idx2[1] ),
    .ZN(_05297_));
 AND2_X1 _14942_ (.A1(_05296_),
    .A2(_05297_),
    .ZN(_05298_));
 INV_X1 _14943_ (.A(_00041_),
    .ZN(_05299_));
 NOR3_X2 _14944_ (.A1(_00853_),
    .A2(_00860_),
    .A3(_05299_),
    .ZN(_05300_));
 NAND3_X2 _14945_ (.A1(_00841_),
    .A2(_00851_),
    .A3(_05300_),
    .ZN(_05301_));
 NOR2_X2 _14946_ (.A1(_01109_),
    .A2(_05301_),
    .ZN(_05302_));
 INV_X1 _14947_ (.A(_08570_),
    .ZN(_05303_));
 INV_X1 _14948_ (.A(_08581_),
    .ZN(_05304_));
 INV_X1 _14949_ (.A(_08585_),
    .ZN(_05305_));
 BUF_X2 _14950_ (.A(_08586_),
    .Z(_05306_));
 INV_X2 _14951_ (.A(_08591_),
    .ZN(_05307_));
 INV_X1 _14952_ (.A(_08595_),
    .ZN(_05308_));
 INV_X1 _14953_ (.A(_08601_),
    .ZN(_05309_));
 INV_X1 _14954_ (.A(_08605_),
    .ZN(_05310_));
 CLKBUF_X2 _14955_ (.A(_08606_),
    .Z(_05311_));
 INV_X2 _14956_ (.A(_08611_),
    .ZN(_05312_));
 INV_X1 _14957_ (.A(_08615_),
    .ZN(_05313_));
 INV_X1 _14958_ (.A(_08620_),
    .ZN(_05314_));
 INV_X1 _14959_ (.A(_08630_),
    .ZN(_05315_));
 INV_X1 _14960_ (.A(_08631_),
    .ZN(_05316_));
 OAI21_X1 _14961_ (.A(_05315_),
    .B1(_07352_),
    .B2(_05316_),
    .ZN(_05317_));
 BUF_X8 clone129 (.A(net475),
    .Z(net129));
 AOI21_X4 _14963_ (.A(_08625_),
    .B1(_05317_),
    .B2(net493),
    .ZN(_05319_));
 INV_X2 _14964_ (.A(_08621_),
    .ZN(_05320_));
 OAI21_X1 _14965_ (.A(_05314_),
    .B1(_05319_),
    .B2(_05320_),
    .ZN(_05321_));
 NAND2_X1 _14966_ (.A1(_08616_),
    .A2(_05321_),
    .ZN(_05322_));
 AOI21_X2 _14967_ (.A(_05312_),
    .B1(_05322_),
    .B2(_05313_),
    .ZN(_05323_));
 OAI21_X2 _14968_ (.A(_05311_),
    .B1(_08610_),
    .B2(_05323_),
    .ZN(_05324_));
 AOI21_X2 _14969_ (.A(_05309_),
    .B1(_05324_),
    .B2(_05310_),
    .ZN(_05325_));
 OAI21_X2 _14970_ (.A(_08596_),
    .B1(_08600_),
    .B2(_05325_),
    .ZN(_05326_));
 AOI21_X2 _14971_ (.A(_05307_),
    .B1(_05326_),
    .B2(_05308_),
    .ZN(_05327_));
 OAI21_X2 _14972_ (.A(_05306_),
    .B1(_08590_),
    .B2(_05327_),
    .ZN(_05328_));
 AOI21_X2 _14973_ (.A(_05304_),
    .B1(_05305_),
    .B2(_05328_),
    .ZN(_05329_));
 OAI21_X2 _14974_ (.A(_08576_),
    .B1(_08580_),
    .B2(_05329_),
    .ZN(_05330_));
 INV_X2 _14975_ (.A(_05330_),
    .ZN(_05331_));
 OAI21_X4 _14976_ (.A(_08571_),
    .B1(_08575_),
    .B2(_05331_),
    .ZN(_05332_));
 NAND2_X1 _14977_ (.A1(_05303_),
    .A2(_05332_),
    .ZN(_05333_));
 AOI21_X2 _14978_ (.A(_08554_),
    .B1(_05333_),
    .B2(_08566_),
    .ZN(_05334_));
 XNOR2_X1 _14979_ (.A(\temp_imag[0] ),
    .B(_08561_),
    .ZN(_05335_));
 XNOR2_X2 _14980_ (.A(_05334_),
    .B(_05335_),
    .ZN(_05336_));
 NAND3_X4 _14981_ (.A1(\temp_imag[0] ),
    .A2(_08564_),
    .A3(_05336_),
    .ZN(_05337_));
 AND2_X4 _14982_ (.A1(_05337_),
    .A2(_05302_),
    .ZN(_05338_));
 BUF_X16 clone132 (.A(_05657_),
    .Z(net132));
 INV_X4 _14984_ (.A(_05338_),
    .ZN(_05340_));
 OR2_X4 _14985_ (.A1(_01311_),
    .A2(_05301_),
    .ZN(_05341_));
 OAI21_X4 _14986_ (.A(_05340_),
    .B1(_05341_),
    .B2(_05337_),
    .ZN(_05342_));
 NAND2_X1 _14987_ (.A1(_05298_),
    .A2(net153),
    .ZN(_05343_));
 CLKBUF_X2 _14988_ (.A(_00038_),
    .Z(_05344_));
 BUF_X2 _14989_ (.A(_00026_),
    .Z(_05345_));
 BUF_X2 _14990_ (.A(_00028_),
    .Z(_05346_));
 NAND3_X2 _14991_ (.A1(_05344_),
    .A2(_05345_),
    .A3(_05346_),
    .ZN(_05347_));
 BUF_X2 _14992_ (.A(_00039_),
    .Z(_05348_));
 INV_X1 _14993_ (.A(_00029_),
    .ZN(_05349_));
 INV_X1 _14994_ (.A(\sample_count[2] ),
    .ZN(_05350_));
 AND2_X2 _14995_ (.A1(_05350_),
    .A2(_09378_),
    .ZN(_05351_));
 NOR2_X1 _14996_ (.A1(_00860_),
    .A2(_00846_),
    .ZN(_05352_));
 AND3_X2 _14997_ (.A1(net86),
    .A2(_00858_),
    .A3(_05352_),
    .ZN(_05353_));
 NAND2_X2 _14998_ (.A1(_00841_),
    .A2(_05353_),
    .ZN(_05354_));
 NOR3_X4 _14999_ (.A1(_05349_),
    .A2(_05351_),
    .A3(_05354_),
    .ZN(_05355_));
 NAND3_X2 _15000_ (.A1(_05348_),
    .A2(_00027_),
    .A3(_05355_),
    .ZN(_05356_));
 OR2_X1 _15001_ (.A1(_01109_),
    .A2(_05301_),
    .ZN(_05357_));
 BUF_X4 _15002_ (.A(_05357_),
    .Z(_05358_));
 INV_X1 _15003_ (.A(_08567_),
    .ZN(_05359_));
 INV_X1 _15004_ (.A(_08577_),
    .ZN(_05360_));
 INV_X1 _15005_ (.A(_08587_),
    .ZN(_05361_));
 INV_X1 _15006_ (.A(_08597_),
    .ZN(_05362_));
 INV_X1 _15007_ (.A(_08607_),
    .ZN(_05363_));
 INV_X1 _15008_ (.A(_08617_),
    .ZN(_05364_));
 INV_X1 _15009_ (.A(_08627_),
    .ZN(_05365_));
 AOI21_X2 _15010_ (.A(_08632_),
    .B1(_08556_),
    .B2(_05316_),
    .ZN(_05366_));
 OAI21_X2 _15011_ (.A(_05365_),
    .B1(_08626_),
    .B2(_05366_),
    .ZN(_05367_));
 AOI21_X2 _15012_ (.A(_08622_),
    .B1(_05367_),
    .B2(_05320_),
    .ZN(_05368_));
 OAI21_X2 _15013_ (.A(_05364_),
    .B1(_08616_),
    .B2(_05368_),
    .ZN(_05369_));
 AOI21_X2 _15014_ (.A(_08612_),
    .B1(_05369_),
    .B2(_05312_),
    .ZN(_05370_));
 OAI21_X2 _15015_ (.A(_05363_),
    .B1(_05311_),
    .B2(_05370_),
    .ZN(_05371_));
 AOI21_X2 _15016_ (.A(_08602_),
    .B1(_05371_),
    .B2(_05309_),
    .ZN(_05372_));
 OAI21_X2 _15017_ (.A(_05362_),
    .B1(_05372_),
    .B2(_08596_),
    .ZN(_05373_));
 AOI21_X2 _15018_ (.A(_08592_),
    .B1(_05373_),
    .B2(_05307_),
    .ZN(_05374_));
 OAI21_X2 _15019_ (.A(_05361_),
    .B1(_05306_),
    .B2(_05374_),
    .ZN(_05375_));
 AOI21_X1 _15020_ (.A(_08582_),
    .B1(_05375_),
    .B2(_05304_),
    .ZN(_05376_));
 OAI21_X2 _15021_ (.A(_05360_),
    .B1(_05376_),
    .B2(_08576_),
    .ZN(_05377_));
 INV_X1 _15022_ (.A(_08571_),
    .ZN(_05378_));
 AOI21_X2 _15023_ (.A(_08572_),
    .B1(_05377_),
    .B2(_05378_),
    .ZN(_05379_));
 OAI21_X2 _15024_ (.A(_05359_),
    .B1(_05379_),
    .B2(_08555_),
    .ZN(_05380_));
 XNOR2_X1 _15025_ (.A(_07347_),
    .B(_08561_),
    .ZN(_05381_));
 XNOR2_X2 _15026_ (.A(_05380_),
    .B(_05381_),
    .ZN(_05382_));
 OAI21_X4 _15027_ (.A(_05365_),
    .B1(_07350_),
    .B2(net495),
    .ZN(_05383_));
 AOI21_X4 _15028_ (.A(_08622_),
    .B1(_05383_),
    .B2(_05320_),
    .ZN(_05384_));
 OAI21_X4 _15029_ (.A(_05364_),
    .B1(_05384_),
    .B2(_08616_),
    .ZN(_05385_));
 AOI21_X4 _15030_ (.A(_08612_),
    .B1(_05385_),
    .B2(_05312_),
    .ZN(_05386_));
 OAI21_X4 _15031_ (.A(_05363_),
    .B1(_05386_),
    .B2(_05311_),
    .ZN(_05387_));
 AOI21_X4 _15032_ (.A(_08602_),
    .B1(_05387_),
    .B2(_05309_),
    .ZN(_05388_));
 OAI21_X4 _15033_ (.A(_05362_),
    .B1(_05388_),
    .B2(_08596_),
    .ZN(_05389_));
 AOI21_X4 _15034_ (.A(_08592_),
    .B1(_05389_),
    .B2(_05307_),
    .ZN(_05390_));
 OAI21_X4 _15035_ (.A(_05361_),
    .B1(_05390_),
    .B2(_05306_),
    .ZN(_05391_));
 AOI21_X4 _15036_ (.A(_08582_),
    .B1(_05391_),
    .B2(_05304_),
    .ZN(_05392_));
 OAI21_X4 _15037_ (.A(_05360_),
    .B1(_05392_),
    .B2(_08576_),
    .ZN(_05393_));
 AOI21_X4 _15038_ (.A(_08572_),
    .B1(_05393_),
    .B2(_05378_),
    .ZN(_05394_));
 XNOR2_X2 _15039_ (.A(_05394_),
    .B(_08555_),
    .ZN(_05395_));
 XNOR2_X2 _15040_ (.A(_05378_),
    .B(net509),
    .ZN(_05396_));
 XNOR2_X2 _15041_ (.A(_05307_),
    .B(net506),
    .ZN(_05397_));
 XNOR2_X2 _15042_ (.A(_05306_),
    .B(net499),
    .ZN(_05398_));
 XNOR2_X1 _15043_ (.A(_05312_),
    .B(_05369_),
    .ZN(_05399_));
 XNOR2_X1 _15044_ (.A(_05311_),
    .B(net507),
    .ZN(_05400_));
 XNOR2_X2 _15045_ (.A(_05320_),
    .B(net489),
    .ZN(_05401_));
 INV_X2 _15046_ (.A(_08558_),
    .ZN(_05402_));
 XOR2_X2 _15047_ (.A(net494),
    .B(net500),
    .Z(_05403_));
 INV_X1 _15048_ (.A(_08616_),
    .ZN(_05404_));
 XNOR2_X2 _15049_ (.A(_05404_),
    .B(net505),
    .ZN(_05405_));
 NOR4_X2 _15050_ (.A1(_05405_),
    .A2(_05402_),
    .A3(_05403_),
    .A4(_07351_),
    .ZN(_05406_));
 NAND4_X1 _15051_ (.A1(_05406_),
    .A2(_05400_),
    .A3(_05401_),
    .A4(_05399_),
    .ZN(_05407_));
 INV_X1 _15052_ (.A(_08596_),
    .ZN(_05408_));
 XNOR2_X2 _15053_ (.A(_05408_),
    .B(net502),
    .ZN(_05409_));
 XNOR2_X2 _15054_ (.A(_08601_),
    .B(net510),
    .ZN(_05410_));
 NOR3_X2 _15055_ (.A1(_05407_),
    .A2(_05409_),
    .A3(_05410_),
    .ZN(_05411_));
 NAND3_X2 _15056_ (.A1(_05398_),
    .A2(_05397_),
    .A3(_05411_),
    .ZN(_05412_));
 INV_X1 _15057_ (.A(_08576_),
    .ZN(_05413_));
 XNOR2_X2 _15058_ (.A(_05413_),
    .B(net504),
    .ZN(_05414_));
 XNOR2_X2 _15059_ (.A(_08581_),
    .B(net503),
    .ZN(_05415_));
 NOR3_X4 _15060_ (.A1(_05414_),
    .A2(_05412_),
    .A3(_05415_),
    .ZN(_05416_));
 NAND3_X2 _15061_ (.A1(_05416_),
    .A2(_05396_),
    .A3(_05395_),
    .ZN(_05417_));
 AND4_X4 _15062_ (.A1(\temp_imag[0] ),
    .A2(_05417_),
    .A3(_05382_),
    .A4(_08563_),
    .ZN(_05418_));
 MUX2_X2 _15063_ (.A(_05358_),
    .B(_05341_),
    .S(_05418_),
    .Z(_05419_));
 BUF_X4 clone125 (.A(_05419_),
    .Z(net125));
 MUX2_X2 _15065_ (.A(_05347_),
    .B(_05356_),
    .S(net138),
    .Z(_05421_));
 MUX2_X2 clone137 (.A(_05347_),
    .B(_05356_),
    .S(net138),
    .Z(net137));
 AOI21_X4 _15067_ (.A(_00843_),
    .B1(_05351_),
    .B2(_05353_),
    .ZN(_05423_));
 AND3_X4 _15068_ (.A1(_05421_),
    .A2(_05343_),
    .A3(_05423_),
    .ZN(_05424_));
 BUF_X8 _15069_ (.A(_05424_),
    .Z(_05425_));
 NAND2_X1 _15070_ (.A1(\samples_imag[0][0] ),
    .A2(net140),
    .ZN(_05426_));
 NOR2_X4 _15071_ (.A1(_05358_),
    .A2(_05418_),
    .ZN(_05427_));
 BUF_X8 _15072_ (.A(_05427_),
    .Z(_05428_));
 BUF_X8 _15073_ (.A(_05419_),
    .Z(_05429_));
 BUF_X16 _15074_ (.A(_05429_),
    .Z(_05430_));
 AOI22_X4 _15075_ (.A1(_05402_),
    .A2(_05428_),
    .B1(net45),
    .B2(_05430_),
    .ZN(_05431_));
 AND3_X1 _15076_ (.A1(_00841_),
    .A2(_05351_),
    .A3(_05353_),
    .ZN(_05432_));
 BUF_X1 _15077_ (.A(_05432_),
    .Z(_05433_));
 CLKBUF_X3 _15078_ (.A(_05433_),
    .Z(_05434_));
 NAND2_X1 _15079_ (.A1(net45),
    .A2(_05434_),
    .ZN(_05435_));
 BUF_X4 _15080_ (.A(_05421_),
    .Z(_05436_));
 MUX2_X1 _15081_ (.A(_05431_),
    .B(_05435_),
    .S(_05436_),
    .Z(_05437_));
 AND2_X2 _15082_ (.A1(_05298_),
    .A2(net153),
    .ZN(_05438_));
 CLKBUF_X3 _15083_ (.A(_05438_),
    .Z(_05439_));
 NAND2_X4 _15084_ (.A1(_05296_),
    .A2(_05297_),
    .ZN(_05440_));
 CLKBUF_X3 _15085_ (.A(_05440_),
    .Z(_05441_));
 NAND2_X4 _15086_ (.A1(_05402_),
    .A2(net520),
    .ZN(_05442_));
 OAI221_X1 _15087_ (.A(_05426_),
    .B1(_05437_),
    .B2(_05439_),
    .C1(_05441_),
    .C2(_05442_),
    .ZN(_00325_));
 NAND2_X1 _15088_ (.A1(\samples_imag[0][10] ),
    .A2(net140),
    .ZN(_05443_));
 NOR3_X2 _15089_ (.A1(_05358_),
    .A2(_05398_),
    .A3(net496),
    .ZN(_05444_));
 AOI21_X4 _15090_ (.A(_05444_),
    .B1(_05430_),
    .B2(net46),
    .ZN(_05445_));
 NAND2_X1 _15091_ (.A1(net46),
    .A2(_05434_),
    .ZN(_05446_));
 MUX2_X1 _15092_ (.A(_05445_),
    .B(_05446_),
    .S(_05436_),
    .Z(_05447_));
 BUF_X4 _15093_ (.A(_05340_),
    .Z(_05448_));
 INV_X1 _15094_ (.A(_05306_),
    .ZN(_05449_));
 INV_X1 _15095_ (.A(_08590_),
    .ZN(_05450_));
 INV_X1 _15096_ (.A(_08600_),
    .ZN(_05451_));
 INV_X1 _15097_ (.A(_05311_),
    .ZN(_05452_));
 INV_X1 _15098_ (.A(_08610_),
    .ZN(_05453_));
 INV_X1 _15099_ (.A(net494),
    .ZN(_05454_));
 NOR2_X2 _15100_ (.A1(_05454_),
    .A2(_07353_),
    .ZN(_05455_));
 OAI21_X1 _15101_ (.A(_08621_),
    .B1(_08625_),
    .B2(_05455_),
    .ZN(_05456_));
 AOI21_X1 _15102_ (.A(_05404_),
    .B1(_05314_),
    .B2(_05456_),
    .ZN(_05457_));
 OAI21_X1 _15103_ (.A(_08611_),
    .B1(_08615_),
    .B2(_05457_),
    .ZN(_05458_));
 AOI21_X2 _15104_ (.A(_05452_),
    .B1(_05453_),
    .B2(_05458_),
    .ZN(_05459_));
 OAI21_X1 _15105_ (.A(_08601_),
    .B1(_08605_),
    .B2(_05459_),
    .ZN(_05460_));
 AOI21_X2 _15106_ (.A(_05408_),
    .B1(_05451_),
    .B2(_05460_),
    .ZN(_05461_));
 OAI21_X1 _15107_ (.A(_08591_),
    .B1(_08595_),
    .B2(_05461_),
    .ZN(_05462_));
 AND3_X1 _15108_ (.A1(_05449_),
    .A2(_05450_),
    .A3(_05462_),
    .ZN(_05463_));
 AOI21_X2 _15109_ (.A(_05449_),
    .B1(_05450_),
    .B2(_05462_),
    .ZN(_05464_));
 OR3_X4 _15110_ (.A1(_05448_),
    .A2(_05463_),
    .A3(_05464_),
    .ZN(_05465_));
 BUF_X16 clone156 (.A(_05695_),
    .Z(net156));
 OAI221_X1 _15112_ (.A(_05443_),
    .B1(_05447_),
    .B2(_05439_),
    .C1(_05441_),
    .C2(_05465_),
    .ZN(_00326_));
 NAND2_X1 _15113_ (.A1(\samples_imag[0][11] ),
    .A2(net140),
    .ZN(_05467_));
 AOI22_X4 _15114_ (.A1(_05415_),
    .A2(_05428_),
    .B1(net47),
    .B2(_05430_),
    .ZN(_05468_));
 NAND2_X1 _15115_ (.A1(net47),
    .A2(_05434_),
    .ZN(_05469_));
 MUX2_X1 _15116_ (.A(_05468_),
    .B(_05469_),
    .S(_05436_),
    .Z(_05470_));
 AND3_X1 _15117_ (.A1(_05304_),
    .A2(_05305_),
    .A3(_05328_),
    .ZN(_05471_));
 OR3_X4 _15118_ (.A1(_05329_),
    .A2(_05448_),
    .A3(_05471_),
    .ZN(_05472_));
 BUF_X4 clone149 (.A(_05622_),
    .Z(net149));
 OAI221_X1 _15120_ (.A(_05467_),
    .B1(_05470_),
    .B2(_05439_),
    .C1(_05441_),
    .C2(_05472_),
    .ZN(_00327_));
 NAND2_X1 _15121_ (.A1(\samples_imag[0][12] ),
    .A2(net140),
    .ZN(_05474_));
 AOI22_X4 _15122_ (.A1(net512),
    .A2(_05428_),
    .B1(net48),
    .B2(_05430_),
    .ZN(_05475_));
 NAND2_X1 _15123_ (.A1(net48),
    .A2(_05434_),
    .ZN(_05476_));
 MUX2_X1 _15124_ (.A(_05475_),
    .B(_05476_),
    .S(_05436_),
    .Z(_05477_));
 INV_X1 _15125_ (.A(_08580_),
    .ZN(_05478_));
 OAI21_X1 _15126_ (.A(_08581_),
    .B1(_08585_),
    .B2(_05464_),
    .ZN(_05479_));
 AND3_X1 _15127_ (.A1(_05413_),
    .A2(_05478_),
    .A3(_05479_),
    .ZN(_05480_));
 AOI21_X2 _15128_ (.A(_05413_),
    .B1(_05478_),
    .B2(_05479_),
    .ZN(_05481_));
 OR3_X4 _15129_ (.A1(_05448_),
    .A2(_05480_),
    .A3(_05481_),
    .ZN(_05482_));
 BUF_X8 clone154 (.A(_05791_),
    .Z(net154));
 OAI221_X1 _15131_ (.A(_05474_),
    .B1(_05477_),
    .B2(_05439_),
    .C1(_05441_),
    .C2(_05482_),
    .ZN(_00328_));
 NAND2_X1 _15132_ (.A1(\samples_imag[0][13] ),
    .A2(_05425_),
    .ZN(_05484_));
 NOR3_X2 _15133_ (.A1(_05358_),
    .A2(_05396_),
    .A3(net496),
    .ZN(_05485_));
 AOI21_X4 _15134_ (.A(_05485_),
    .B1(_05430_),
    .B2(net49),
    .ZN(_05486_));
 NAND2_X1 _15135_ (.A1(net49),
    .A2(_05434_),
    .ZN(_05487_));
 MUX2_X1 _15136_ (.A(_05486_),
    .B(_05487_),
    .S(_05436_),
    .Z(_05488_));
 OR3_X2 _15137_ (.A1(_08571_),
    .A2(_08575_),
    .A3(_05331_),
    .ZN(_05489_));
 NAND3_X4 _15138_ (.A1(_05332_),
    .A2(net520),
    .A3(_05489_),
    .ZN(_05490_));
 OAI221_X1 _15139_ (.A(_05484_),
    .B1(_05488_),
    .B2(_05439_),
    .C1(_05441_),
    .C2(_05490_),
    .ZN(_00329_));
 NAND2_X1 _15140_ (.A1(\samples_imag[0][14] ),
    .A2(_05425_),
    .ZN(_05491_));
 XOR2_X2 _15141_ (.A(_08555_),
    .B(net498),
    .Z(_05492_));
 AOI22_X4 _15142_ (.A1(_05492_),
    .A2(_05428_),
    .B1(_05430_),
    .B2(net50),
    .ZN(_05493_));
 CLKBUF_X3 _15143_ (.A(_05433_),
    .Z(_05494_));
 NAND2_X1 _15144_ (.A1(net50),
    .A2(_05494_),
    .ZN(_05495_));
 MUX2_X1 _15145_ (.A(_05493_),
    .B(_05495_),
    .S(_05421_),
    .Z(_05496_));
 OAI21_X1 _15146_ (.A(_08571_),
    .B1(_08575_),
    .B2(_05481_),
    .ZN(_05497_));
 NAND2_X1 _15147_ (.A1(_05303_),
    .A2(_05497_),
    .ZN(_05498_));
 XOR2_X2 _15148_ (.A(_08566_),
    .B(_05498_),
    .Z(_05499_));
 NAND2_X4 _15149_ (.A1(net520),
    .A2(_05499_),
    .ZN(_05500_));
 OAI221_X1 _15150_ (.A(_05491_),
    .B1(_05496_),
    .B2(_05439_),
    .C1(_05441_),
    .C2(_05500_),
    .ZN(_00330_));
 OR2_X2 _15151_ (.A1(_05358_),
    .A2(_05336_),
    .ZN(_05501_));
 INV_X1 _15152_ (.A(net54),
    .ZN(_05502_));
 AOI22_X4 _15153_ (.A1(net501),
    .A2(_05427_),
    .B1(_05429_),
    .B2(_05502_),
    .ZN(_05503_));
 NOR2_X1 _15154_ (.A1(net139),
    .A2(_05503_),
    .ZN(_05504_));
 AOI22_X1 _15155_ (.A1(net54),
    .A2(_05434_),
    .B1(_05423_),
    .B2(\samples_imag[0][15] ),
    .ZN(_05505_));
 AOI21_X1 _15156_ (.A(_05504_),
    .B1(_05505_),
    .B2(net139),
    .ZN(_05506_));
 MUX2_X1 _15157_ (.A(_05501_),
    .B(_05506_),
    .S(_05343_),
    .Z(_00331_));
 NAND2_X4 _15158_ (.A1(_05425_),
    .A2(\samples_imag[0][1] ),
    .ZN(_05507_));
 AOI22_X4 _15159_ (.A1(_07351_),
    .A2(_05428_),
    .B1(net55),
    .B2(_05430_),
    .ZN(_05508_));
 NAND2_X1 _15160_ (.A1(net55),
    .A2(_05494_),
    .ZN(_05509_));
 MUX2_X1 _15161_ (.A(_05508_),
    .B(_05509_),
    .S(_05421_),
    .Z(_05510_));
 NAND2_X4 _15162_ (.A1(_07354_),
    .A2(net520),
    .ZN(_05511_));
 OAI221_X2 _15163_ (.A(_05507_),
    .B1(_05510_),
    .B2(_05439_),
    .C1(_05441_),
    .C2(_05511_),
    .ZN(_00332_));
 AND2_X1 _15164_ (.A1(_05454_),
    .A2(_07353_),
    .ZN(_05512_));
 NOR3_X4 _15165_ (.A1(_05448_),
    .A2(_05455_),
    .A3(_05512_),
    .ZN(_05513_));
 NAND2_X1 _15166_ (.A1(_05439_),
    .A2(_05513_),
    .ZN(_05514_));
 AOI22_X4 _15167_ (.A1(_05403_),
    .A2(_05428_),
    .B1(net62),
    .B2(_05430_),
    .ZN(_05515_));
 AOI22_X1 _15168_ (.A1(net62),
    .A2(_05434_),
    .B1(_05423_),
    .B2(\samples_imag[0][2] ),
    .ZN(_05516_));
 MUX2_X1 _15169_ (.A(_05515_),
    .B(_05516_),
    .S(net139),
    .Z(_05517_));
 OAI21_X1 _15170_ (.A(_05514_),
    .B1(_05517_),
    .B2(_05439_),
    .ZN(_00333_));
 NAND3_X1 _15171_ (.A1(net63),
    .A2(net139),
    .A3(_05434_),
    .ZN(_05518_));
 NOR3_X2 _15172_ (.A1(_05358_),
    .A2(_05401_),
    .A3(_05418_),
    .ZN(_05519_));
 AOI21_X4 _15173_ (.A(_05519_),
    .B1(net63),
    .B2(_05430_),
    .ZN(_05520_));
 OAI21_X1 _15174_ (.A(_05518_),
    .B1(_05520_),
    .B2(net139),
    .ZN(_05521_));
 NAND2_X1 _15175_ (.A1(_05343_),
    .A2(_05521_),
    .ZN(_05522_));
 XNOR2_X2 _15176_ (.A(_05320_),
    .B(_05319_),
    .ZN(_05523_));
 NOR2_X4 _15177_ (.A1(_05448_),
    .A2(_05523_),
    .ZN(_05524_));
 AOI22_X1 _15178_ (.A1(net140),
    .A2(\samples_imag[0][3] ),
    .B1(_05524_),
    .B2(_05298_),
    .ZN(_05525_));
 NAND2_X1 _15179_ (.A1(_05525_),
    .A2(_05522_),
    .ZN(_00334_));
 NAND2_X1 _15180_ (.A1(\samples_imag[0][4] ),
    .A2(_05425_),
    .ZN(_05526_));
 AOI22_X4 _15181_ (.A1(_05405_),
    .A2(_05427_),
    .B1(net125),
    .B2(net64),
    .ZN(_05527_));
 NAND2_X1 _15182_ (.A1(net64),
    .A2(_05494_),
    .ZN(_05528_));
 MUX2_X1 _15183_ (.A(_05527_),
    .B(_05528_),
    .S(_05421_),
    .Z(_05529_));
 AND3_X1 _15184_ (.A1(_05404_),
    .A2(_05314_),
    .A3(_05456_),
    .ZN(_05530_));
 NOR2_X1 _15185_ (.A1(_05457_),
    .A2(_05530_),
    .ZN(_05531_));
 NAND2_X2 _15186_ (.A1(net520),
    .A2(_05531_),
    .ZN(_05532_));
 OAI221_X1 _15187_ (.A(_05526_),
    .B1(_05529_),
    .B2(_05439_),
    .C1(_05441_),
    .C2(_05532_),
    .ZN(_00335_));
 NAND2_X1 _15188_ (.A1(\samples_imag[0][5] ),
    .A2(_05425_),
    .ZN(_05533_));
 INV_X1 _15189_ (.A(_05399_),
    .ZN(_05534_));
 AOI22_X4 _15190_ (.A1(_05534_),
    .A2(_05428_),
    .B1(net125),
    .B2(net65),
    .ZN(_05535_));
 NAND2_X1 _15191_ (.A1(net65),
    .A2(_05494_),
    .ZN(_05536_));
 MUX2_X1 _15192_ (.A(_05535_),
    .B(_05536_),
    .S(net137),
    .Z(_05537_));
 AND3_X1 _15193_ (.A1(_05312_),
    .A2(_05313_),
    .A3(_05322_),
    .ZN(_05538_));
 OR3_X4 _15194_ (.A1(_05323_),
    .A2(_05448_),
    .A3(_05538_),
    .ZN(_05539_));
 OAI221_X1 _15195_ (.A(_05533_),
    .B1(_05537_),
    .B2(_05438_),
    .C1(_05441_),
    .C2(_05539_),
    .ZN(_00336_));
 NAND2_X1 _15196_ (.A1(_05424_),
    .A2(\samples_imag[0][6] ),
    .ZN(_05540_));
 INV_X1 _15197_ (.A(_05400_),
    .ZN(_05541_));
 AOI22_X4 _15198_ (.A1(_05541_),
    .A2(_05428_),
    .B1(net125),
    .B2(net66),
    .ZN(_05542_));
 NAND2_X1 _15199_ (.A1(net66),
    .A2(_05494_),
    .ZN(_05543_));
 MUX2_X1 _15200_ (.A(_05542_),
    .B(_05543_),
    .S(net137),
    .Z(_05544_));
 AND3_X1 _15201_ (.A1(_05452_),
    .A2(_05453_),
    .A3(_05458_),
    .ZN(_05545_));
 OR3_X4 _15202_ (.A1(_05448_),
    .A2(_05459_),
    .A3(_05545_),
    .ZN(_05546_));
 OAI21_X4 clone153 (.A(_05340_),
    .B1(_05337_),
    .B2(_05341_),
    .ZN(net153));
 OAI221_X1 _15204_ (.A(_05540_),
    .B1(_05544_),
    .B2(_05438_),
    .C1(_05441_),
    .C2(_05546_),
    .ZN(_00337_));
 NAND2_X1 _15205_ (.A1(_05424_),
    .A2(\samples_imag[0][7] ),
    .ZN(_05548_));
 AOI22_X4 _15206_ (.A1(_05410_),
    .A2(_05428_),
    .B1(net125),
    .B2(net67),
    .ZN(_05549_));
 NAND2_X1 _15207_ (.A1(net67),
    .A2(_05494_),
    .ZN(_05550_));
 MUX2_X1 _15208_ (.A(_05549_),
    .B(_05550_),
    .S(net137),
    .Z(_05551_));
 CLKBUF_X3 _15209_ (.A(_05440_),
    .Z(_05552_));
 AND3_X1 _15210_ (.A1(_05309_),
    .A2(_05310_),
    .A3(_05324_),
    .ZN(_05553_));
 OR3_X4 _15211_ (.A1(_05325_),
    .A2(_05448_),
    .A3(_05553_),
    .ZN(_05554_));
 BUF_X8 clone152 (.A(_05798_),
    .Z(net152));
 OAI221_X1 _15213_ (.A(_05548_),
    .B1(_05551_),
    .B2(_05438_),
    .C1(_05552_),
    .C2(_05554_),
    .ZN(_00338_));
 NAND2_X1 _15214_ (.A1(\samples_imag[0][8] ),
    .A2(_05424_),
    .ZN(_05556_));
 AOI22_X4 _15215_ (.A1(_05409_),
    .A2(_05428_),
    .B1(net125),
    .B2(net68),
    .ZN(_05557_));
 NAND2_X1 _15216_ (.A1(net68),
    .A2(_05494_),
    .ZN(_05558_));
 MUX2_X1 _15217_ (.A(_05557_),
    .B(_05558_),
    .S(net137),
    .Z(_05559_));
 AND3_X1 _15218_ (.A1(_05408_),
    .A2(_05451_),
    .A3(_05460_),
    .ZN(_05560_));
 OR3_X4 _15219_ (.A1(_05448_),
    .A2(_05461_),
    .A3(_05560_),
    .ZN(_05561_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 OAI221_X1 _15221_ (.A(_05556_),
    .B1(_05559_),
    .B2(_05438_),
    .C1(_05552_),
    .C2(_05561_),
    .ZN(_00339_));
 NAND2_X1 _15222_ (.A1(\samples_imag[0][9] ),
    .A2(_05424_),
    .ZN(_05563_));
 NOR3_X2 _15223_ (.A1(_05358_),
    .A2(_05397_),
    .A3(net496),
    .ZN(_05564_));
 AOI21_X4 _15224_ (.A(_05564_),
    .B1(_05430_),
    .B2(net69),
    .ZN(_05565_));
 NAND2_X1 _15225_ (.A1(net69),
    .A2(_05494_),
    .ZN(_05566_));
 MUX2_X1 _15226_ (.A(_05565_),
    .B(_05566_),
    .S(net137),
    .Z(_05567_));
 AND3_X1 _15227_ (.A1(_05307_),
    .A2(_05308_),
    .A3(_05326_),
    .ZN(_05568_));
 OR3_X4 _15228_ (.A1(_05327_),
    .A2(_05448_),
    .A3(_05568_),
    .ZN(_05569_));
 BUF_X8 clone158 (.A(_05727_),
    .Z(net158));
 OAI221_X1 _15230_ (.A(_05563_),
    .B1(_05567_),
    .B2(_05438_),
    .C1(_05552_),
    .C2(_05569_),
    .ZN(_00340_));
 BUF_X4 _15231_ (.A(_00842_),
    .Z(_05571_));
 INV_X1 _15232_ (.A(_05344_),
    .ZN(_05572_));
 NAND3_X1 _15233_ (.A1(_05572_),
    .A2(_05345_),
    .A3(_05346_),
    .ZN(_05573_));
 INV_X1 _15234_ (.A(_00027_),
    .ZN(_05574_));
 NOR2_X1 _15235_ (.A1(_05348_),
    .A2(_05574_),
    .ZN(_05575_));
 NAND2_X1 _15236_ (.A1(_05355_),
    .A2(_05575_),
    .ZN(_05576_));
 MUX2_X2 _15237_ (.A(_05573_),
    .B(_05576_),
    .S(_05429_),
    .Z(_05577_));
 NAND3_X4 _15238_ (.A1(_04790_),
    .A2(_05297_),
    .A3(net526),
    .ZN(_05578_));
 AND3_X4 _15239_ (.A1(_05571_),
    .A2(net488),
    .A3(_05578_),
    .ZN(_05579_));
 AND3_X4 clone151 (.A1(_05571_),
    .A2(net488),
    .A3(_05578_),
    .ZN(net151));
 NAND2_X1 _15241_ (.A1(\samples_imag[1][0] ),
    .A2(net151),
    .ZN(_05581_));
 NAND2_X2 _15242_ (.A1(_04790_),
    .A2(_05297_),
    .ZN(_05582_));
 CLKBUF_X3 _15243_ (.A(_05582_),
    .Z(_05583_));
 INV_X4 _15244_ (.A(net513),
    .ZN(_05584_));
 NAND2_X4 _15245_ (.A1(_05584_),
    .A2(_05578_),
    .ZN(_05585_));
 OAI221_X1 _15246_ (.A(_05581_),
    .B1(_05583_),
    .B2(_05442_),
    .C1(net530),
    .C2(_05585_),
    .ZN(_00341_));
 NAND2_X1 _15247_ (.A1(\samples_imag[1][10] ),
    .A2(_05579_),
    .ZN(_05586_));
 OAI221_X1 _15248_ (.A(_05586_),
    .B1(_05583_),
    .B2(_05465_),
    .C1(_05445_),
    .C2(_05585_),
    .ZN(_00342_));
 NAND2_X1 _15249_ (.A1(_05579_),
    .A2(\samples_imag[1][11] ),
    .ZN(_05587_));
 OAI221_X1 _15250_ (.A(_05587_),
    .B1(_05583_),
    .B2(_05472_),
    .C1(net528),
    .C2(_05585_),
    .ZN(_00343_));
 NAND2_X1 _15251_ (.A1(_05579_),
    .A2(\samples_imag[1][12] ),
    .ZN(_05588_));
 OAI221_X1 _15252_ (.A(_05588_),
    .B1(_05583_),
    .B2(_05482_),
    .C1(net529),
    .C2(_05585_),
    .ZN(_00344_));
 NAND2_X1 _15253_ (.A1(_05579_),
    .A2(\samples_imag[1][13] ),
    .ZN(_05589_));
 OAI221_X1 _15254_ (.A(_05589_),
    .B1(_05583_),
    .B2(_05490_),
    .C1(_05486_),
    .C2(_05585_),
    .ZN(_00345_));
 NAND2_X1 _15255_ (.A1(_05579_),
    .A2(\samples_imag[1][14] ),
    .ZN(_05590_));
 OAI221_X1 _15256_ (.A(_05590_),
    .B1(_05583_),
    .B2(_05500_),
    .C1(_05493_),
    .C2(_05585_),
    .ZN(_00346_));
 NAND2_X2 _15257_ (.A1(_05503_),
    .A2(_05584_),
    .ZN(_05591_));
 BUF_X8 _15258_ (.A(_05577_),
    .Z(_05592_));
 NAND3_X1 _15259_ (.A1(_00856_),
    .A2(\samples_imag[1][15] ),
    .A3(_05592_),
    .ZN(_05593_));
 NAND2_X1 _15260_ (.A1(_05591_),
    .A2(_05593_),
    .ZN(_05594_));
 MUX2_X1 _15261_ (.A(_05501_),
    .B(_05594_),
    .S(_05578_),
    .Z(_00347_));
 NAND2_X1 _15262_ (.A1(net151),
    .A2(\samples_imag[1][1] ),
    .ZN(_05595_));
 OAI221_X1 _15263_ (.A(_05595_),
    .B1(_05582_),
    .B2(_05511_),
    .C1(net531),
    .C2(_05585_),
    .ZN(_00348_));
 CLKBUF_X3 _15264_ (.A(_00855_),
    .Z(_05596_));
 NAND3_X1 _15265_ (.A1(_05596_),
    .A2(\samples_imag[1][2] ),
    .A3(_05592_),
    .ZN(_05597_));
 OAI21_X1 _15266_ (.A(_05597_),
    .B1(net144),
    .B2(_05515_),
    .ZN(_05598_));
 MUX2_X1 _15267_ (.A(_05513_),
    .B(_05598_),
    .S(_05578_),
    .Z(_00349_));
 NAND3_X4 _15268_ (.A1(_05596_),
    .A2(\samples_imag[1][3] ),
    .A3(_05592_),
    .ZN(_05599_));
 OAI21_X2 _15269_ (.A(_05599_),
    .B1(net144),
    .B2(_05520_),
    .ZN(_05600_));
 MUX2_X1 _15270_ (.A(_05524_),
    .B(_05600_),
    .S(_05578_),
    .Z(_00350_));
 AND2_X1 _15271_ (.A1(net520),
    .A2(_05531_),
    .ZN(_05601_));
 NAND3_X4 _15272_ (.A1(_05596_),
    .A2(\samples_imag[1][4] ),
    .A3(_05592_),
    .ZN(_05602_));
 OAI21_X2 _15273_ (.A(_05602_),
    .B1(net144),
    .B2(_05527_),
    .ZN(_05603_));
 MUX2_X1 _15274_ (.A(_05601_),
    .B(_05603_),
    .S(_05578_),
    .Z(_00351_));
 INV_X1 _15275_ (.A(_05539_),
    .ZN(_05604_));
 NAND3_X4 _15276_ (.A1(_05596_),
    .A2(\samples_imag[1][5] ),
    .A3(_05592_),
    .ZN(_05605_));
 OAI21_X2 _15277_ (.A(_05605_),
    .B1(net144),
    .B2(_05535_),
    .ZN(_05606_));
 MUX2_X1 _15278_ (.A(_05604_),
    .B(_05606_),
    .S(_05578_),
    .Z(_00352_));
 INV_X1 _15279_ (.A(_05546_),
    .ZN(_05607_));
 NAND3_X1 _15280_ (.A1(_05596_),
    .A2(net534),
    .A3(\samples_imag[1][6] ),
    .ZN(_05608_));
 OAI21_X2 _15281_ (.A(_05608_),
    .B1(net144),
    .B2(_05542_),
    .ZN(_05609_));
 MUX2_X1 _15282_ (.A(_05607_),
    .B(_05609_),
    .S(_05578_),
    .Z(_00353_));
 NAND2_X4 _15283_ (.A1(net151),
    .A2(\samples_imag[1][7] ),
    .ZN(_05610_));
 OAI221_X2 _15284_ (.A(_05610_),
    .B1(_05582_),
    .B2(_05554_),
    .C1(_05549_),
    .C2(_05585_),
    .ZN(_00354_));
 NAND2_X1 _15285_ (.A1(net151),
    .A2(\samples_imag[1][8] ),
    .ZN(_05611_));
 OAI221_X1 _15286_ (.A(_05611_),
    .B1(_05582_),
    .B2(_05561_),
    .C1(_05557_),
    .C2(_05585_),
    .ZN(_00355_));
 NAND2_X1 _15287_ (.A1(net151),
    .A2(\samples_imag[1][9] ),
    .ZN(_05612_));
 OAI221_X1 _15288_ (.A(_05612_),
    .B1(_05582_),
    .B2(_05569_),
    .C1(_05565_),
    .C2(_05585_),
    .ZN(_00356_));
 INV_X1 _15289_ (.A(_05345_),
    .ZN(_05613_));
 NAND3_X1 _15290_ (.A1(_05344_),
    .A2(_05613_),
    .A3(_05346_),
    .ZN(_05614_));
 NAND3_X2 _15291_ (.A1(_05348_),
    .A2(_05574_),
    .A3(_05355_),
    .ZN(_05615_));
 MUX2_X2 _15292_ (.A(_05614_),
    .B(_05615_),
    .S(net138),
    .Z(_05616_));
 MUX2_X2 clone133 (.A(_05614_),
    .B(_05615_),
    .S(net138),
    .Z(net133));
 INV_X1 _15294_ (.A(_04794_),
    .ZN(_05618_));
 NAND2_X2 _15295_ (.A1(_05618_),
    .A2(_04791_),
    .ZN(_05619_));
 NOR2_X2 _15296_ (.A1(_04790_),
    .A2(_05619_),
    .ZN(_05620_));
 NAND2_X2 _15297_ (.A1(net153),
    .A2(_05620_),
    .ZN(_05621_));
 AND3_X2 _15298_ (.A1(_00842_),
    .A2(_05616_),
    .A3(_05621_),
    .ZN(_05622_));
 BUF_X4 _15299_ (.A(_05622_),
    .Z(_05623_));
 NAND2_X1 _15300_ (.A1(\samples_imag[2][0] ),
    .A2(net149),
    .ZN(_05624_));
 OR2_X1 _15301_ (.A1(_04790_),
    .A2(_05619_),
    .ZN(_05625_));
 CLKBUF_X3 _15302_ (.A(_05625_),
    .Z(_05626_));
 CLKBUF_X3 _15303_ (.A(_05626_),
    .Z(_05627_));
 INV_X2 _15304_ (.A(_05616_),
    .ZN(_05628_));
 NAND2_X2 _15305_ (.A1(_05628_),
    .A2(_05621_),
    .ZN(_05629_));
 BUF_X4 _15306_ (.A(_05629_),
    .Z(_05630_));
 OAI221_X1 _15307_ (.A(_05624_),
    .B1(_05627_),
    .B2(_05442_),
    .C1(net530),
    .C2(_05630_),
    .ZN(_00357_));
 NAND2_X1 _15308_ (.A1(\samples_imag[2][10] ),
    .A2(net149),
    .ZN(_05631_));
 OAI221_X1 _15309_ (.A(_05631_),
    .B1(_05627_),
    .B2(_05465_),
    .C1(_05445_),
    .C2(_05630_),
    .ZN(_00358_));
 NAND2_X1 _15310_ (.A1(\samples_imag[2][11] ),
    .A2(_05623_),
    .ZN(_05632_));
 OAI221_X1 _15311_ (.A(_05632_),
    .B1(_05627_),
    .B2(_05472_),
    .C1(net528),
    .C2(_05630_),
    .ZN(_00359_));
 NAND2_X1 _15312_ (.A1(\samples_imag[2][12] ),
    .A2(_05623_),
    .ZN(_05633_));
 OAI221_X1 _15313_ (.A(_05633_),
    .B1(_05627_),
    .B2(_05482_),
    .C1(net529),
    .C2(_05630_),
    .ZN(_00360_));
 NAND2_X1 _15314_ (.A1(\samples_imag[2][13] ),
    .A2(net149),
    .ZN(_05634_));
 OAI221_X1 _15315_ (.A(_05634_),
    .B1(_05627_),
    .B2(_05490_),
    .C1(_05486_),
    .C2(_05630_),
    .ZN(_00361_));
 NAND2_X1 _15316_ (.A1(\samples_imag[2][14] ),
    .A2(net149),
    .ZN(_05635_));
 OAI221_X1 _15317_ (.A(_05635_),
    .B1(_05627_),
    .B2(_05500_),
    .C1(_05493_),
    .C2(_05630_),
    .ZN(_00362_));
 NAND2_X1 _15318_ (.A1(_05503_),
    .A2(_05628_),
    .ZN(_05636_));
 NAND3_X1 _15319_ (.A1(_00856_),
    .A2(\samples_imag[2][15] ),
    .A3(net133),
    .ZN(_05637_));
 NAND2_X1 _15320_ (.A1(_05636_),
    .A2(_05637_),
    .ZN(_05638_));
 MUX2_X1 _15321_ (.A(_05501_),
    .B(_05638_),
    .S(_05621_),
    .Z(_00363_));
 NAND2_X1 _15322_ (.A1(\samples_imag[2][1] ),
    .A2(net149),
    .ZN(_05639_));
 OAI221_X1 _15323_ (.A(_05639_),
    .B1(_05626_),
    .B2(_05511_),
    .C1(net531),
    .C2(_05630_),
    .ZN(_00364_));
 NAND3_X1 _15324_ (.A1(_05596_),
    .A2(\samples_imag[2][2] ),
    .A3(_05616_),
    .ZN(_05640_));
 OAI21_X1 _15325_ (.A(_05640_),
    .B1(_05515_),
    .B2(net133),
    .ZN(_05641_));
 MUX2_X1 _15326_ (.A(_05513_),
    .B(_05641_),
    .S(_05621_),
    .Z(_00365_));
 NAND3_X1 _15327_ (.A1(_05596_),
    .A2(\samples_imag[2][3] ),
    .A3(_05616_),
    .ZN(_05642_));
 OAI21_X1 _15328_ (.A(_05642_),
    .B1(_05520_),
    .B2(net133),
    .ZN(_05643_));
 MUX2_X1 _15329_ (.A(_05524_),
    .B(_05643_),
    .S(_05621_),
    .Z(_00366_));
 NAND3_X1 _15330_ (.A1(_05596_),
    .A2(\samples_imag[2][4] ),
    .A3(_05616_),
    .ZN(_05644_));
 OAI21_X1 _15331_ (.A(_05644_),
    .B1(net133),
    .B2(_05527_),
    .ZN(_05645_));
 MUX2_X1 _15332_ (.A(_05601_),
    .B(_05645_),
    .S(_05621_),
    .Z(_00367_));
 NAND2_X1 _15333_ (.A1(\samples_imag[2][5] ),
    .A2(_05623_),
    .ZN(_05646_));
 OAI221_X1 _15334_ (.A(_05646_),
    .B1(_05626_),
    .B2(_05539_),
    .C1(_05535_),
    .C2(_05630_),
    .ZN(_00368_));
 NAND2_X1 _15335_ (.A1(\samples_imag[2][6] ),
    .A2(_05623_),
    .ZN(_05647_));
 OAI221_X1 _15336_ (.A(_05647_),
    .B1(_05626_),
    .B2(_05546_),
    .C1(_05542_),
    .C2(_05630_),
    .ZN(_00369_));
 NAND2_X1 _15337_ (.A1(_05623_),
    .A2(\samples_imag[2][7] ),
    .ZN(_05648_));
 OAI221_X1 _15338_ (.A(_05648_),
    .B1(_05626_),
    .B2(_05554_),
    .C1(_05549_),
    .C2(_05630_),
    .ZN(_00370_));
 NAND2_X1 _15339_ (.A1(_05622_),
    .A2(\samples_imag[2][8] ),
    .ZN(_05649_));
 OAI221_X1 _15340_ (.A(_05649_),
    .B1(_05626_),
    .B2(_05561_),
    .C1(_05557_),
    .C2(_05629_),
    .ZN(_00371_));
 NAND2_X1 _15341_ (.A1(_05622_),
    .A2(\samples_imag[2][9] ),
    .ZN(_05650_));
 OAI221_X1 _15342_ (.A(_05650_),
    .B1(_05626_),
    .B2(_05569_),
    .C1(_05565_),
    .C2(_05629_),
    .ZN(_00372_));
 NAND3_X1 _15343_ (.A1(_05572_),
    .A2(_05613_),
    .A3(_05346_),
    .ZN(_05651_));
 NOR2_X1 _15344_ (.A1(_05348_),
    .A2(_00027_),
    .ZN(_05652_));
 NAND2_X1 _15345_ (.A1(_05355_),
    .A2(_05652_),
    .ZN(_05653_));
 MUX2_X2 _15346_ (.A(_05651_),
    .B(_05653_),
    .S(_05429_),
    .Z(_05654_));
 NOR2_X2 _15347_ (.A1(_05296_),
    .A2(_05619_),
    .ZN(_05655_));
 NAND2_X2 _15348_ (.A1(net526),
    .A2(_05655_),
    .ZN(_05656_));
 AND3_X4 _15349_ (.A1(_05654_),
    .A2(_05656_),
    .A3(_05571_),
    .ZN(_05657_));
 BUF_X16 _15350_ (.A(_05657_),
    .Z(_05658_));
 NAND2_X4 _15351_ (.A1(\samples_imag[3][0] ),
    .A2(net132),
    .ZN(_05659_));
 OR2_X1 _15352_ (.A1(_05296_),
    .A2(_05619_),
    .ZN(_05660_));
 CLKBUF_X3 _15353_ (.A(_05660_),
    .Z(_05661_));
 CLKBUF_X3 _15354_ (.A(_05661_),
    .Z(_05662_));
 INV_X2 _15355_ (.A(_05654_),
    .ZN(_05663_));
 NAND2_X2 _15356_ (.A1(_05663_),
    .A2(_05656_),
    .ZN(_05664_));
 BUF_X4 _15357_ (.A(_05664_),
    .Z(_05665_));
 OAI221_X2 _15358_ (.A(_05659_),
    .B1(_05662_),
    .B2(_05442_),
    .C1(net530),
    .C2(_05665_),
    .ZN(_00373_));
 NAND2_X4 _15359_ (.A1(\samples_imag[3][10] ),
    .A2(net132),
    .ZN(_05666_));
 OAI221_X2 _15360_ (.A(_05666_),
    .B1(_05662_),
    .B2(_05465_),
    .C1(_05445_),
    .C2(_05665_),
    .ZN(_00374_));
 NAND2_X4 _15361_ (.A1(\samples_imag[3][11] ),
    .A2(_05658_),
    .ZN(_05667_));
 OAI221_X2 _15362_ (.A(_05667_),
    .B1(_05662_),
    .B2(_05472_),
    .C1(net528),
    .C2(_05665_),
    .ZN(_00375_));
 NAND2_X4 _15363_ (.A1(_05658_),
    .A2(\samples_imag[3][12] ),
    .ZN(_05668_));
 OAI221_X2 _15364_ (.A(_05668_),
    .B1(_05662_),
    .B2(_05482_),
    .C1(net529),
    .C2(_05665_),
    .ZN(_00376_));
 NAND2_X4 _15365_ (.A1(_05658_),
    .A2(\samples_imag[3][13] ),
    .ZN(_05669_));
 OAI221_X2 _15366_ (.A(_05669_),
    .B1(_05662_),
    .B2(_05490_),
    .C1(_05486_),
    .C2(_05665_),
    .ZN(_00377_));
 NAND2_X4 _15367_ (.A1(_05658_),
    .A2(\samples_imag[3][14] ),
    .ZN(_05670_));
 OAI221_X2 _15368_ (.A(_05670_),
    .B1(_05662_),
    .B2(_05500_),
    .C1(_05493_),
    .C2(_05665_),
    .ZN(_00378_));
 NAND2_X1 _15369_ (.A1(_05503_),
    .A2(_05663_),
    .ZN(_05671_));
 CLKBUF_X3 _15370_ (.A(_00855_),
    .Z(_05672_));
 NAND3_X1 _15371_ (.A1(_05672_),
    .A2(\samples_imag[3][15] ),
    .A3(_05654_),
    .ZN(_05673_));
 NAND2_X1 _15372_ (.A1(_05671_),
    .A2(_05673_),
    .ZN(_05674_));
 MUX2_X1 _15373_ (.A(_05501_),
    .B(_05674_),
    .S(_05656_),
    .Z(_00379_));
 NAND2_X4 _15374_ (.A1(net132),
    .A2(\samples_imag[3][1] ),
    .ZN(_05675_));
 OAI221_X2 _15375_ (.A(_05675_),
    .B1(_05661_),
    .B2(_05511_),
    .C1(net531),
    .C2(_05665_),
    .ZN(_00380_));
 CLKBUF_X3 _15376_ (.A(_05571_),
    .Z(_05676_));
 NAND3_X1 _15377_ (.A1(_05676_),
    .A2(_05654_),
    .A3(\samples_imag[3][2] ),
    .ZN(_05677_));
 OAI21_X1 _15378_ (.A(_05677_),
    .B1(_05654_),
    .B2(_05515_),
    .ZN(_05678_));
 MUX2_X1 _15379_ (.A(_05513_),
    .B(_05678_),
    .S(_05656_),
    .Z(_00381_));
 AOI22_X1 _15380_ (.A1(_05524_),
    .A2(_05655_),
    .B1(_05657_),
    .B2(\samples_imag[3][3] ),
    .ZN(_05679_));
 OAI21_X1 _15381_ (.A(_05679_),
    .B1(_05665_),
    .B2(_05520_),
    .ZN(_00382_));
 NAND2_X4 _15382_ (.A1(net132),
    .A2(\samples_imag[3][4] ),
    .ZN(_05680_));
 OAI221_X2 _15383_ (.A(_05680_),
    .B1(_05661_),
    .B2(_05532_),
    .C1(_05527_),
    .C2(_05665_),
    .ZN(_00383_));
 NAND2_X4 _15384_ (.A1(net132),
    .A2(\samples_imag[3][5] ),
    .ZN(_05681_));
 OAI221_X2 _15385_ (.A(_05681_),
    .B1(_05661_),
    .B2(_05539_),
    .C1(_05535_),
    .C2(_05665_),
    .ZN(_00384_));
 NAND2_X4 _15386_ (.A1(_05658_),
    .A2(\samples_imag[3][6] ),
    .ZN(_05682_));
 OAI221_X2 _15387_ (.A(_05682_),
    .B1(_05661_),
    .B2(_05546_),
    .C1(_05542_),
    .C2(_05664_),
    .ZN(_00385_));
 NAND2_X1 _15388_ (.A1(_05657_),
    .A2(\samples_imag[3][7] ),
    .ZN(_05683_));
 OAI221_X1 _15389_ (.A(_05683_),
    .B1(_05661_),
    .B2(_05554_),
    .C1(_05549_),
    .C2(_05664_),
    .ZN(_00386_));
 NAND2_X1 _15390_ (.A1(_05657_),
    .A2(\samples_imag[3][8] ),
    .ZN(_05684_));
 OAI221_X1 _15391_ (.A(_05684_),
    .B1(_05661_),
    .B2(_05561_),
    .C1(_05557_),
    .C2(_05664_),
    .ZN(_00387_));
 NAND2_X1 _15392_ (.A1(_05657_),
    .A2(\samples_imag[3][9] ),
    .ZN(_05685_));
 OAI221_X1 _15393_ (.A(_05685_),
    .B1(_05661_),
    .B2(_05569_),
    .C1(_05565_),
    .C2(_05664_),
    .ZN(_00388_));
 INV_X1 _15394_ (.A(_05346_),
    .ZN(_05686_));
 NAND3_X1 _15395_ (.A1(_05344_),
    .A2(_05345_),
    .A3(_05686_),
    .ZN(_05687_));
 NOR3_X2 _15396_ (.A1(_00029_),
    .A2(_05351_),
    .A3(_05354_),
    .ZN(_05688_));
 NAND3_X1 _15397_ (.A1(_05348_),
    .A2(_00027_),
    .A3(_05688_),
    .ZN(_05689_));
 MUX2_X2 _15398_ (.A(_05687_),
    .B(_05689_),
    .S(net497),
    .Z(_05690_));
 OR3_X1 _15399_ (.A1(_05618_),
    .A2(_04791_),
    .A3(\idx2[0] ),
    .ZN(_05691_));
 BUF_X4 _15400_ (.A(_05691_),
    .Z(_05692_));
 INV_X1 _15401_ (.A(_05692_),
    .ZN(_05693_));
 NAND2_X2 _15402_ (.A1(net526),
    .A2(_05693_),
    .ZN(_05694_));
 AND3_X4 _15403_ (.A1(_05571_),
    .A2(_05694_),
    .A3(_05690_),
    .ZN(_05695_));
 BUF_X8 _15404_ (.A(_05695_),
    .Z(_05696_));
 NAND2_X4 _15405_ (.A1(net156),
    .A2(\samples_imag[4][0] ),
    .ZN(_05697_));
 BUF_X4 _15406_ (.A(_05692_),
    .Z(_05698_));
 INV_X2 _15407_ (.A(_05690_),
    .ZN(_05699_));
 NAND2_X2 _15408_ (.A1(_05699_),
    .A2(_05694_),
    .ZN(_05700_));
 BUF_X4 _15409_ (.A(_05700_),
    .Z(_05701_));
 OAI221_X2 _15410_ (.A(_05697_),
    .B1(_05698_),
    .B2(_05442_),
    .C1(net530),
    .C2(_05701_),
    .ZN(_00389_));
 NAND2_X4 _15411_ (.A1(\samples_imag[4][10] ),
    .A2(net156),
    .ZN(_05702_));
 OAI221_X2 _15412_ (.A(_05702_),
    .B1(_05698_),
    .B2(_05465_),
    .C1(_05445_),
    .C2(_05701_),
    .ZN(_00390_));
 NAND2_X4 _15413_ (.A1(\samples_imag[4][11] ),
    .A2(_05696_),
    .ZN(_05703_));
 OAI221_X2 _15414_ (.A(_05703_),
    .B1(_05698_),
    .B2(_05472_),
    .C1(net528),
    .C2(_05701_),
    .ZN(_00391_));
 NAND2_X4 _15415_ (.A1(\samples_imag[4][12] ),
    .A2(_05696_),
    .ZN(_05704_));
 OAI221_X2 _15416_ (.A(_05704_),
    .B1(_05698_),
    .B2(_05482_),
    .C1(net529),
    .C2(_05701_),
    .ZN(_00392_));
 NAND2_X2 _15417_ (.A1(\samples_imag[4][13] ),
    .A2(_05696_),
    .ZN(_05705_));
 OAI221_X1 _15418_ (.A(_05705_),
    .B1(_05698_),
    .B2(_05490_),
    .C1(_05486_),
    .C2(_05701_),
    .ZN(_00393_));
 NAND2_X4 _15419_ (.A1(net156),
    .A2(\samples_imag[4][14] ),
    .ZN(_05706_));
 OAI221_X2 _15420_ (.A(_05706_),
    .B1(_05698_),
    .B2(_05500_),
    .C1(_05493_),
    .C2(_05701_),
    .ZN(_00394_));
 NAND2_X1 _15421_ (.A1(_05503_),
    .A2(_05699_),
    .ZN(_05707_));
 NAND3_X1 _15422_ (.A1(_05672_),
    .A2(\samples_imag[4][15] ),
    .A3(_05690_),
    .ZN(_05708_));
 NAND2_X1 _15423_ (.A1(_05707_),
    .A2(_05708_),
    .ZN(_05709_));
 MUX2_X1 _15424_ (.A(_05501_),
    .B(_05709_),
    .S(_05694_),
    .Z(_00395_));
 NAND2_X4 _15425_ (.A1(net156),
    .A2(\samples_imag[4][1] ),
    .ZN(_05710_));
 OAI221_X2 _15426_ (.A(_05710_),
    .B1(_05692_),
    .B2(_05511_),
    .C1(net531),
    .C2(_05701_),
    .ZN(_00396_));
 NAND3_X1 _15427_ (.A1(_05676_),
    .A2(\samples_imag[4][2] ),
    .A3(_05690_),
    .ZN(_05711_));
 OAI21_X1 _15428_ (.A(_05711_),
    .B1(_05515_),
    .B2(_05690_),
    .ZN(_05712_));
 MUX2_X1 _15429_ (.A(_05513_),
    .B(_05712_),
    .S(_05694_),
    .Z(_00397_));
 NAND3_X1 _15430_ (.A1(_05676_),
    .A2(\samples_imag[4][3] ),
    .A3(_05690_),
    .ZN(_05713_));
 OAI21_X1 _15431_ (.A(_05713_),
    .B1(_05690_),
    .B2(_05520_),
    .ZN(_05714_));
 MUX2_X1 _15432_ (.A(_05524_),
    .B(_05714_),
    .S(_05694_),
    .Z(_00398_));
 NAND2_X4 _15433_ (.A1(_05696_),
    .A2(\samples_imag[4][4] ),
    .ZN(_05715_));
 OAI221_X2 _15434_ (.A(_05715_),
    .B1(_05692_),
    .B2(_05532_),
    .C1(_05527_),
    .C2(_05701_),
    .ZN(_00399_));
 NAND2_X4 _15435_ (.A1(net156),
    .A2(\samples_imag[4][5] ),
    .ZN(_05716_));
 OAI221_X2 _15436_ (.A(_05716_),
    .B1(_05692_),
    .B2(_05539_),
    .C1(_05535_),
    .C2(_05701_),
    .ZN(_00400_));
 NAND2_X4 _15437_ (.A1(_05696_),
    .A2(\samples_imag[4][6] ),
    .ZN(_05717_));
 OAI221_X2 _15438_ (.A(_05717_),
    .B1(_05692_),
    .B2(_05546_),
    .C1(_05542_),
    .C2(_05701_),
    .ZN(_00401_));
 NAND2_X1 _15439_ (.A1(_05695_),
    .A2(\samples_imag[4][7] ),
    .ZN(_05718_));
 OAI221_X1 _15440_ (.A(_05718_),
    .B1(_05692_),
    .B2(_05554_),
    .C1(_05549_),
    .C2(_05700_),
    .ZN(_00402_));
 NAND2_X1 _15441_ (.A1(_05695_),
    .A2(\samples_imag[4][8] ),
    .ZN(_05719_));
 OAI221_X1 _15442_ (.A(_05719_),
    .B1(_05692_),
    .B2(_05561_),
    .C1(_05557_),
    .C2(_05700_),
    .ZN(_00403_));
 NAND2_X1 _15443_ (.A1(_05695_),
    .A2(\samples_imag[4][9] ),
    .ZN(_05720_));
 OAI221_X1 _15444_ (.A(_05720_),
    .B1(_05692_),
    .B2(_05569_),
    .C1(_05565_),
    .C2(_05700_),
    .ZN(_00404_));
 NAND3_X1 _15445_ (.A1(_05572_),
    .A2(_05345_),
    .A3(_05686_),
    .ZN(_05721_));
 NAND2_X1 _15446_ (.A1(_05575_),
    .A2(_05688_),
    .ZN(_05722_));
 MUX2_X2 _15447_ (.A(_05721_),
    .B(_05722_),
    .S(net497),
    .Z(_05723_));
 NAND2_X1 _15448_ (.A1(_04794_),
    .A2(_04790_),
    .ZN(_05724_));
 NOR2_X2 _15449_ (.A1(_04791_),
    .A2(_05724_),
    .ZN(_05725_));
 NAND2_X2 _15450_ (.A1(net526),
    .A2(_05725_),
    .ZN(_05726_));
 AND3_X4 _15451_ (.A1(_05571_),
    .A2(_05726_),
    .A3(_05723_),
    .ZN(_05727_));
 BUF_X8 _15452_ (.A(_05727_),
    .Z(_05728_));
 NAND2_X4 _15453_ (.A1(net158),
    .A2(\samples_imag[5][0] ),
    .ZN(_05729_));
 OR2_X1 _15454_ (.A1(_04791_),
    .A2(_05724_),
    .ZN(_05730_));
 BUF_X4 _15455_ (.A(_05730_),
    .Z(_05731_));
 BUF_X4 _15456_ (.A(_05731_),
    .Z(_05732_));
 INV_X2 _15457_ (.A(_05723_),
    .ZN(_05733_));
 NAND2_X2 _15458_ (.A1(_05733_),
    .A2(_05726_),
    .ZN(_05734_));
 BUF_X4 _15459_ (.A(_05734_),
    .Z(_05735_));
 OAI221_X2 _15460_ (.A(_05729_),
    .B1(_05732_),
    .B2(_05442_),
    .C1(net530),
    .C2(_05735_),
    .ZN(_00405_));
 NAND2_X4 _15461_ (.A1(\samples_imag[5][10] ),
    .A2(net158),
    .ZN(_05736_));
 OAI221_X2 _15462_ (.A(_05736_),
    .B1(_05732_),
    .B2(_05465_),
    .C1(_05445_),
    .C2(_05735_),
    .ZN(_00406_));
 NAND2_X4 _15463_ (.A1(\samples_imag[5][11] ),
    .A2(_05728_),
    .ZN(_05737_));
 OAI221_X2 _15464_ (.A(_05737_),
    .B1(_05732_),
    .B2(_05472_),
    .C1(net528),
    .C2(_05735_),
    .ZN(_00407_));
 NAND2_X4 _15465_ (.A1(\samples_imag[5][12] ),
    .A2(_05728_),
    .ZN(_05738_));
 OAI221_X2 _15466_ (.A(_05738_),
    .B1(_05732_),
    .B2(_05482_),
    .C1(net529),
    .C2(_05735_),
    .ZN(_00408_));
 NAND2_X4 _15467_ (.A1(_05728_),
    .A2(\samples_imag[5][13] ),
    .ZN(_05739_));
 OAI221_X2 _15468_ (.A(_05739_),
    .B1(_05732_),
    .B2(_05490_),
    .C1(_05486_),
    .C2(_05735_),
    .ZN(_00409_));
 NAND2_X2 _15469_ (.A1(\samples_imag[5][14] ),
    .A2(net158),
    .ZN(_05740_));
 OAI221_X1 _15470_ (.A(_05740_),
    .B1(_05732_),
    .B2(_05500_),
    .C1(_05493_),
    .C2(_05735_),
    .ZN(_00410_));
 NAND2_X1 _15471_ (.A1(_05503_),
    .A2(_05733_),
    .ZN(_05741_));
 NAND3_X1 _15472_ (.A1(_05672_),
    .A2(\samples_imag[5][15] ),
    .A3(_05723_),
    .ZN(_05742_));
 NAND2_X1 _15473_ (.A1(_05741_),
    .A2(_05742_),
    .ZN(_05743_));
 MUX2_X1 _15474_ (.A(_05501_),
    .B(_05743_),
    .S(_05726_),
    .Z(_00411_));
 NAND2_X2 _15475_ (.A1(\samples_imag[5][1] ),
    .A2(net158),
    .ZN(_05744_));
 OAI221_X1 _15476_ (.A(_05744_),
    .B1(_05731_),
    .B2(_05511_),
    .C1(net531),
    .C2(_05735_),
    .ZN(_00412_));
 NAND3_X1 _15477_ (.A1(_05676_),
    .A2(\samples_imag[5][2] ),
    .A3(_05723_),
    .ZN(_05745_));
 OAI21_X1 _15478_ (.A(_05745_),
    .B1(_05515_),
    .B2(net527),
    .ZN(_05746_));
 MUX2_X1 _15479_ (.A(_05513_),
    .B(_05746_),
    .S(_05726_),
    .Z(_00413_));
 NAND3_X1 _15480_ (.A1(_05676_),
    .A2(_05723_),
    .A3(\samples_imag[5][3] ),
    .ZN(_05747_));
 OAI21_X1 _15481_ (.A(_05747_),
    .B1(_05723_),
    .B2(_05520_),
    .ZN(_05748_));
 MUX2_X1 _15482_ (.A(_05524_),
    .B(_05748_),
    .S(_05726_),
    .Z(_00414_));
 NAND2_X4 _15483_ (.A1(\samples_imag[5][4] ),
    .A2(_05728_),
    .ZN(_05749_));
 OAI221_X2 _15484_ (.A(_05749_),
    .B1(_05731_),
    .B2(_05532_),
    .C1(_05527_),
    .C2(_05735_),
    .ZN(_00415_));
 NAND2_X4 _15485_ (.A1(net158),
    .A2(\samples_imag[5][5] ),
    .ZN(_05750_));
 OAI221_X2 _15486_ (.A(_05750_),
    .B1(_05731_),
    .B2(_05539_),
    .C1(_05535_),
    .C2(_05735_),
    .ZN(_00416_));
 NAND2_X4 _15487_ (.A1(_05728_),
    .A2(\samples_imag[5][6] ),
    .ZN(_05751_));
 OAI221_X2 _15488_ (.A(_05751_),
    .B1(_05731_),
    .B2(_05546_),
    .C1(_05542_),
    .C2(_05735_),
    .ZN(_00417_));
 NAND2_X1 _15489_ (.A1(_05727_),
    .A2(\samples_imag[5][7] ),
    .ZN(_05752_));
 OAI221_X1 _15490_ (.A(_05752_),
    .B1(_05731_),
    .B2(_05554_),
    .C1(_05549_),
    .C2(_05734_),
    .ZN(_00418_));
 NAND2_X1 _15491_ (.A1(_05727_),
    .A2(\samples_imag[5][8] ),
    .ZN(_05753_));
 OAI221_X1 _15492_ (.A(_05753_),
    .B1(_05731_),
    .B2(_05561_),
    .C1(_05557_),
    .C2(_05734_),
    .ZN(_00419_));
 NAND2_X1 _15493_ (.A1(_05727_),
    .A2(\samples_imag[5][9] ),
    .ZN(_05754_));
 OAI221_X1 _15494_ (.A(_05754_),
    .B1(_05731_),
    .B2(_05569_),
    .C1(_05565_),
    .C2(_05734_),
    .ZN(_00420_));
 NOR2_X1 _15495_ (.A1(_05345_),
    .A2(_05346_),
    .ZN(_05755_));
 NAND2_X1 _15496_ (.A1(_05344_),
    .A2(_05755_),
    .ZN(_05756_));
 NAND3_X1 _15497_ (.A1(_05348_),
    .A2(_05574_),
    .A3(_05688_),
    .ZN(_05757_));
 MUX2_X2 _15498_ (.A(_05756_),
    .B(_05757_),
    .S(_05429_),
    .Z(_05758_));
 AND3_X1 _15499_ (.A1(_04794_),
    .A2(_04791_),
    .A3(_05296_),
    .ZN(_05759_));
 NAND2_X2 _15500_ (.A1(_05759_),
    .A2(net153),
    .ZN(_05760_));
 AND3_X4 _15501_ (.A1(_05758_),
    .A2(_05571_),
    .A3(_05760_),
    .ZN(_05761_));
 BUF_X16 _15502_ (.A(_05761_),
    .Z(_05762_));
 NAND2_X4 _15503_ (.A1(\samples_imag[6][0] ),
    .A2(net131),
    .ZN(_05763_));
 NAND3_X4 _15504_ (.A1(_04794_),
    .A2(_04791_),
    .A3(_05296_),
    .ZN(_05764_));
 BUF_X4 _15505_ (.A(_05764_),
    .Z(_05765_));
 INV_X2 _15506_ (.A(_05758_),
    .ZN(_05766_));
 NAND2_X2 _15507_ (.A1(_05766_),
    .A2(_05760_),
    .ZN(_05767_));
 BUF_X4 _15508_ (.A(_05767_),
    .Z(_05768_));
 OAI221_X2 _15509_ (.A(_05763_),
    .B1(_05765_),
    .B2(_05442_),
    .C1(_05431_),
    .C2(_05768_),
    .ZN(_00421_));
 NAND2_X4 _15510_ (.A1(net131),
    .A2(\samples_imag[6][10] ),
    .ZN(_05769_));
 OAI221_X2 _15511_ (.A(_05769_),
    .B1(_05765_),
    .B2(_05465_),
    .C1(_05445_),
    .C2(_05768_),
    .ZN(_00422_));
 NAND2_X4 _15512_ (.A1(net131),
    .A2(\samples_imag[6][11] ),
    .ZN(_05770_));
 OAI221_X2 _15513_ (.A(_05770_),
    .B1(_05765_),
    .B2(_05472_),
    .C1(net528),
    .C2(_05768_),
    .ZN(_00423_));
 NAND2_X4 _15514_ (.A1(net131),
    .A2(\samples_imag[6][12] ),
    .ZN(_05771_));
 OAI221_X2 _15515_ (.A(_05771_),
    .B1(_05765_),
    .B2(_05482_),
    .C1(_05475_),
    .C2(_05768_),
    .ZN(_00424_));
 NAND2_X4 _15516_ (.A1(net131),
    .A2(\samples_imag[6][13] ),
    .ZN(_05772_));
 OAI221_X2 _15517_ (.A(_05772_),
    .B1(_05765_),
    .B2(_05490_),
    .C1(_05486_),
    .C2(_05768_),
    .ZN(_00425_));
 NAND2_X4 _15518_ (.A1(_05762_),
    .A2(\samples_imag[6][14] ),
    .ZN(_05773_));
 OAI221_X2 _15519_ (.A(_05773_),
    .B1(_05765_),
    .B2(_05500_),
    .C1(_05493_),
    .C2(_05768_),
    .ZN(_00426_));
 NAND2_X1 _15520_ (.A1(_05503_),
    .A2(_05766_),
    .ZN(_05774_));
 NAND3_X1 _15521_ (.A1(_05672_),
    .A2(\samples_imag[6][15] ),
    .A3(_05758_),
    .ZN(_05775_));
 NAND2_X1 _15522_ (.A1(_05774_),
    .A2(_05775_),
    .ZN(_05776_));
 MUX2_X1 _15523_ (.A(_05501_),
    .B(_05776_),
    .S(_05760_),
    .Z(_00427_));
 NAND2_X4 _15524_ (.A1(_05762_),
    .A2(\samples_imag[6][1] ),
    .ZN(_05777_));
 OAI221_X2 _15525_ (.A(_05777_),
    .B1(_05764_),
    .B2(_05511_),
    .C1(net531),
    .C2(_05768_),
    .ZN(_00428_));
 NAND3_X1 _15526_ (.A1(_05676_),
    .A2(_05758_),
    .A3(\samples_imag[6][2] ),
    .ZN(_05778_));
 OAI21_X1 _15527_ (.A(_05778_),
    .B1(_05758_),
    .B2(_05515_),
    .ZN(_05779_));
 MUX2_X1 _15528_ (.A(_05513_),
    .B(_05779_),
    .S(_05760_),
    .Z(_00429_));
 AOI22_X1 _15529_ (.A1(_05524_),
    .A2(_05759_),
    .B1(_05761_),
    .B2(\samples_imag[6][3] ),
    .ZN(_05780_));
 OAI21_X1 _15530_ (.A(_05780_),
    .B1(_05768_),
    .B2(_05520_),
    .ZN(_00430_));
 NAND2_X4 _15531_ (.A1(_05762_),
    .A2(\samples_imag[6][4] ),
    .ZN(_05781_));
 OAI221_X2 _15532_ (.A(_05781_),
    .B1(_05764_),
    .B2(_05532_),
    .C1(_05527_),
    .C2(_05768_),
    .ZN(_00431_));
 NAND2_X4 _15533_ (.A1(_05762_),
    .A2(\samples_imag[6][5] ),
    .ZN(_05782_));
 OAI221_X2 _15534_ (.A(_05782_),
    .B1(_05764_),
    .B2(_05539_),
    .C1(_05535_),
    .C2(_05768_),
    .ZN(_00432_));
 NAND2_X4 _15535_ (.A1(_05762_),
    .A2(\samples_imag[6][6] ),
    .ZN(_05783_));
 OAI221_X2 _15536_ (.A(_05783_),
    .B1(_05764_),
    .B2(_05546_),
    .C1(_05542_),
    .C2(_05767_),
    .ZN(_00433_));
 NAND2_X1 _15537_ (.A1(_05761_),
    .A2(\samples_imag[6][7] ),
    .ZN(_05784_));
 OAI221_X1 _15538_ (.A(_05784_),
    .B1(_05764_),
    .B2(_05554_),
    .C1(_05549_),
    .C2(_05767_),
    .ZN(_00434_));
 NAND2_X1 _15539_ (.A1(_05761_),
    .A2(\samples_imag[6][8] ),
    .ZN(_05785_));
 OAI221_X1 _15540_ (.A(_05785_),
    .B1(_05764_),
    .B2(_05561_),
    .C1(_05557_),
    .C2(_05767_),
    .ZN(_00435_));
 NAND2_X1 _15541_ (.A1(_05761_),
    .A2(\samples_imag[6][9] ),
    .ZN(_05786_));
 OAI221_X1 _15542_ (.A(_05786_),
    .B1(_05764_),
    .B2(_05569_),
    .C1(_05565_),
    .C2(_05767_),
    .ZN(_00436_));
 NAND2_X1 _15543_ (.A1(_05572_),
    .A2(_05755_),
    .ZN(_05787_));
 NAND2_X1 _15544_ (.A1(_05652_),
    .A2(_05688_),
    .ZN(_05788_));
 MUX2_X1 _15545_ (.A(_05787_),
    .B(_05788_),
    .S(net497),
    .Z(_05789_));
 NAND4_X4 _15546_ (.A1(_05342_),
    .A2(_04791_),
    .A3(_04790_),
    .A4(_04794_),
    .ZN(_05790_));
 AND3_X4 _15547_ (.A1(_00842_),
    .A2(_05790_),
    .A3(_05789_),
    .ZN(_05791_));
 BUF_X8 _15548_ (.A(_05791_),
    .Z(_05792_));
 NAND2_X1 _15549_ (.A1(\samples_imag[7][0] ),
    .A2(net154),
    .ZN(_05793_));
 NAND3_X4 _15550_ (.A1(_04794_),
    .A2(_04791_),
    .A3(_04790_),
    .ZN(_05794_));
 BUF_X4 _15551_ (.A(_05794_),
    .Z(_05795_));
 BUF_X8 _15552_ (.A(_05789_),
    .Z(_05796_));
 INV_X8 _15553_ (.A(_05796_),
    .ZN(_05797_));
 NAND2_X4 _15554_ (.A1(_05797_),
    .A2(_05790_),
    .ZN(_05798_));
 BUF_X8 _15555_ (.A(_05798_),
    .Z(_05799_));
 OAI221_X2 _15556_ (.A(_05793_),
    .B1(_05795_),
    .B2(_05442_),
    .C1(net530),
    .C2(net152),
    .ZN(_00437_));
 NAND2_X2 _15557_ (.A1(\samples_imag[7][10] ),
    .A2(net154),
    .ZN(_05800_));
 OAI221_X2 _15558_ (.A(_05800_),
    .B1(_05795_),
    .B2(_05465_),
    .C1(_05445_),
    .C2(_05799_),
    .ZN(_00438_));
 NAND2_X2 _15559_ (.A1(\samples_imag[7][11] ),
    .A2(_05792_),
    .ZN(_05801_));
 OAI221_X2 _15560_ (.A(_05801_),
    .B1(_05795_),
    .B2(_05472_),
    .C1(net528),
    .C2(_05799_),
    .ZN(_00439_));
 NAND2_X2 _15561_ (.A1(\samples_imag[7][12] ),
    .A2(_05792_),
    .ZN(_05802_));
 OAI221_X2 _15562_ (.A(_05802_),
    .B1(_05795_),
    .B2(_05482_),
    .C1(_05475_),
    .C2(_05799_),
    .ZN(_00440_));
 NAND2_X2 _15563_ (.A1(\samples_imag[7][13] ),
    .A2(net154),
    .ZN(_05803_));
 OAI221_X2 _15564_ (.A(_05803_),
    .B1(_05795_),
    .B2(_05490_),
    .C1(_05486_),
    .C2(_05799_),
    .ZN(_00441_));
 NAND2_X2 _15565_ (.A1(\samples_imag[7][14] ),
    .A2(net154),
    .ZN(_05804_));
 OAI221_X2 _15566_ (.A(_05804_),
    .B1(_05795_),
    .B2(_05500_),
    .C1(_05799_),
    .C2(_05493_),
    .ZN(_00442_));
 NAND2_X2 _15567_ (.A1(_05503_),
    .A2(_05797_),
    .ZN(_05805_));
 NAND3_X1 _15568_ (.A1(_05672_),
    .A2(\samples_imag[7][15] ),
    .A3(net143),
    .ZN(_05806_));
 NAND2_X1 _15569_ (.A1(_05805_),
    .A2(_05806_),
    .ZN(_05807_));
 MUX2_X1 _15570_ (.A(_05501_),
    .B(_05807_),
    .S(_05790_),
    .Z(_00443_));
 NAND2_X1 _15571_ (.A1(net154),
    .A2(\samples_imag[7][1] ),
    .ZN(_05808_));
 OAI221_X2 _15572_ (.A(_05808_),
    .B1(_05794_),
    .B2(_05511_),
    .C1(net152),
    .C2(net531),
    .ZN(_00444_));
 NAND3_X4 _15573_ (.A1(_05676_),
    .A2(\samples_imag[7][2] ),
    .A3(_05796_),
    .ZN(_05809_));
 OAI21_X2 _15574_ (.A(_05809_),
    .B1(net143),
    .B2(_05515_),
    .ZN(_05810_));
 MUX2_X1 _15575_ (.A(_05513_),
    .B(_05810_),
    .S(_05790_),
    .Z(_00445_));
 NAND3_X4 _15576_ (.A1(_05676_),
    .A2(\samples_imag[7][3] ),
    .A3(_05796_),
    .ZN(_05811_));
 OAI21_X2 _15577_ (.A(_05811_),
    .B1(net143),
    .B2(_05520_),
    .ZN(_05812_));
 MUX2_X1 _15578_ (.A(_05524_),
    .B(_05812_),
    .S(_05790_),
    .Z(_00446_));
 NAND3_X4 _15579_ (.A1(_05796_),
    .A2(\samples_imag[7][4] ),
    .A3(_05676_),
    .ZN(_05813_));
 OAI21_X2 _15580_ (.A(_05813_),
    .B1(net143),
    .B2(_05527_),
    .ZN(_05814_));
 MUX2_X1 _15581_ (.A(_05601_),
    .B(_05814_),
    .S(_05790_),
    .Z(_00447_));
 NAND3_X4 _15582_ (.A1(_05796_),
    .A2(\samples_imag[7][5] ),
    .A3(_05676_),
    .ZN(_05815_));
 OAI21_X2 _15583_ (.A(_05815_),
    .B1(net143),
    .B2(_05535_),
    .ZN(_05816_));
 MUX2_X1 _15584_ (.A(_05604_),
    .B(_05816_),
    .S(_05790_),
    .Z(_00448_));
 NAND2_X2 _15585_ (.A1(\samples_imag[7][6] ),
    .A2(_05792_),
    .ZN(_05817_));
 OAI221_X2 _15586_ (.A(_05817_),
    .B1(_05794_),
    .B2(_05546_),
    .C1(_05542_),
    .C2(net152),
    .ZN(_00449_));
 NAND2_X2 _15587_ (.A1(\samples_imag[7][7] ),
    .A2(_05792_),
    .ZN(_05818_));
 OAI221_X2 _15588_ (.A(_05818_),
    .B1(_05794_),
    .B2(_05554_),
    .C1(_05549_),
    .C2(net152),
    .ZN(_00450_));
 NAND2_X2 _15589_ (.A1(_05792_),
    .A2(\samples_imag[7][8] ),
    .ZN(_05819_));
 OAI221_X2 _15590_ (.A(_05819_),
    .B1(_05794_),
    .B2(_05561_),
    .C1(_05557_),
    .C2(net152),
    .ZN(_00451_));
 NAND2_X1 _15591_ (.A1(\samples_imag[7][9] ),
    .A2(_05791_),
    .ZN(_05820_));
 OAI221_X1 _15592_ (.A(_05820_),
    .B1(_05794_),
    .B2(_05569_),
    .C1(_05798_),
    .C2(_05565_),
    .ZN(_00452_));
 INV_X1 _15593_ (.A(_08651_),
    .ZN(_05821_));
 BUF_X2 _15594_ (.A(_08652_),
    .Z(_05822_));
 INV_X1 _15595_ (.A(_08662_),
    .ZN(_05823_));
 INV_X1 _15596_ (.A(_08666_),
    .ZN(_05824_));
 INV_X1 _15597_ (.A(_08672_),
    .ZN(_05825_));
 INV_X1 _15598_ (.A(_08676_),
    .ZN(_05826_));
 INV_X1 _15599_ (.A(_08682_),
    .ZN(_05827_));
 INV_X1 _15600_ (.A(_08686_),
    .ZN(_05828_));
 INV_X1 _15601_ (.A(_08692_),
    .ZN(_05829_));
 INV_X1 _15602_ (.A(_08696_),
    .ZN(_05830_));
 INV_X1 _15603_ (.A(_08701_),
    .ZN(_05831_));
 INV_X1 _15604_ (.A(_08711_),
    .ZN(_05832_));
 INV_X2 _15605_ (.A(_08712_),
    .ZN(_05833_));
 OAI21_X2 _15606_ (.A(_05832_),
    .B1(_07360_),
    .B2(_05833_),
    .ZN(_05834_));
 BUF_X4 clone58 (.A(_05929_),
    .Z(net58));
 AOI21_X4 _15608_ (.A(_08706_),
    .B1(net448),
    .B2(_05834_),
    .ZN(_05836_));
 BUF_X2 clone57 (.A(_00001_),
    .Z(net57));
 INV_X2 _15610_ (.A(_08702_),
    .ZN(_05838_));
 OAI21_X1 _15611_ (.A(_05831_),
    .B1(_05836_),
    .B2(_05838_),
    .ZN(_05839_));
 NAND2_X1 _15612_ (.A1(_08697_),
    .A2(_05839_),
    .ZN(_05840_));
 AOI21_X2 _15613_ (.A(_05829_),
    .B1(_05830_),
    .B2(_05840_),
    .ZN(_05841_));
 OAI21_X2 _15614_ (.A(_08687_),
    .B1(_08691_),
    .B2(_05841_),
    .ZN(_05842_));
 AOI21_X2 _15615_ (.A(_05827_),
    .B1(_05828_),
    .B2(_05842_),
    .ZN(_05843_));
 OAI21_X2 _15616_ (.A(_08677_),
    .B1(_08681_),
    .B2(_05843_),
    .ZN(_05844_));
 AOI21_X2 _15617_ (.A(_05825_),
    .B1(_05826_),
    .B2(_05844_),
    .ZN(_05845_));
 OAI21_X2 _15618_ (.A(_08667_),
    .B1(_08671_),
    .B2(_05845_),
    .ZN(_05846_));
 AOI21_X1 _15619_ (.A(_05823_),
    .B1(_05824_),
    .B2(_05846_),
    .ZN(_05847_));
 OAI21_X1 _15620_ (.A(_08657_),
    .B1(_08661_),
    .B2(_05847_),
    .ZN(_05848_));
 INV_X2 _15621_ (.A(_05848_),
    .ZN(_05849_));
 OAI21_X4 _15622_ (.A(_05822_),
    .B1(_08656_),
    .B2(_05849_),
    .ZN(_05850_));
 NAND2_X1 _15623_ (.A1(_05821_),
    .A2(_05850_),
    .ZN(_05851_));
 AOI21_X2 _15624_ (.A(_08635_),
    .B1(_05851_),
    .B2(_08647_),
    .ZN(_05852_));
 XNOR2_X1 _15625_ (.A(\temp_real[0] ),
    .B(_08642_),
    .ZN(_05853_));
 XNOR2_X2 _15626_ (.A(_05853_),
    .B(_05852_),
    .ZN(_05854_));
 NAND3_X2 _15627_ (.A1(\temp_real[0] ),
    .A2(_08645_),
    .A3(_05854_),
    .ZN(_05855_));
 AND2_X4 _15628_ (.A1(_05855_),
    .A2(_05302_),
    .ZN(_05856_));
 BUF_X8 clone98 (.A(_05932_),
    .Z(net98));
 INV_X2 _15630_ (.A(_05856_),
    .ZN(_05858_));
 OAI21_X4 _15631_ (.A(_05858_),
    .B1(_05855_),
    .B2(_05341_),
    .ZN(_05859_));
 AND2_X4 _15632_ (.A1(_05859_),
    .A2(_05298_),
    .ZN(_05860_));
 MUX2_X2 clone94 (.A(_05347_),
    .B(_05356_),
    .S(net453),
    .Z(net94));
 INV_X1 _15634_ (.A(_05860_),
    .ZN(_05862_));
 INV_X1 _15635_ (.A(_08648_),
    .ZN(_05863_));
 INV_X1 _15636_ (.A(_08658_),
    .ZN(_05864_));
 INV_X1 _15637_ (.A(_08668_),
    .ZN(_05865_));
 INV_X1 _15638_ (.A(_08678_),
    .ZN(_05866_));
 INV_X1 _15639_ (.A(_08688_),
    .ZN(_05867_));
 INV_X1 _15640_ (.A(_08698_),
    .ZN(_05868_));
 INV_X1 _15641_ (.A(_08708_),
    .ZN(_05869_));
 AOI21_X4 _15642_ (.A(_08713_),
    .B1(net481),
    .B2(_05833_),
    .ZN(_05870_));
 OAI21_X4 _15643_ (.A(_05869_),
    .B1(_05870_),
    .B2(net474),
    .ZN(_05871_));
 AOI21_X4 _15644_ (.A(_08703_),
    .B1(_05838_),
    .B2(_05871_),
    .ZN(_05872_));
 OAI21_X4 _15645_ (.A(_05868_),
    .B1(_05872_),
    .B2(_08697_),
    .ZN(_05873_));
 AOI21_X4 _15646_ (.A(_08693_),
    .B1(_05873_),
    .B2(_05829_),
    .ZN(_05874_));
 OAI21_X4 _15647_ (.A(_05867_),
    .B1(_08687_),
    .B2(_05874_),
    .ZN(_05875_));
 AOI21_X4 _15648_ (.A(_08683_),
    .B1(_05875_),
    .B2(_05827_),
    .ZN(_05876_));
 OAI21_X4 _15649_ (.A(_05866_),
    .B1(_08677_),
    .B2(_05876_),
    .ZN(_05877_));
 AOI21_X4 _15650_ (.A(_08673_),
    .B1(_05877_),
    .B2(_05825_),
    .ZN(_05878_));
 OAI21_X4 _15651_ (.A(_05865_),
    .B1(_05878_),
    .B2(_08667_),
    .ZN(_05879_));
 AOI21_X4 _15652_ (.A(_08663_),
    .B1(_05879_),
    .B2(_05823_),
    .ZN(_05880_));
 OAI21_X4 _15653_ (.A(_05864_),
    .B1(_05880_),
    .B2(_08657_),
    .ZN(_05881_));
 INV_X1 _15654_ (.A(_05822_),
    .ZN(_05882_));
 AOI21_X1 _15655_ (.A(_08653_),
    .B1(_05881_),
    .B2(_05882_),
    .ZN(_05883_));
 OAI21_X2 _15656_ (.A(_05863_),
    .B1(_05883_),
    .B2(_08636_),
    .ZN(_05884_));
 XNOR2_X1 _15657_ (.A(_07355_),
    .B(_08642_),
    .ZN(_05885_));
 XNOR2_X2 _15658_ (.A(_05885_),
    .B(_05884_),
    .ZN(_05886_));
 AND2_X1 _15659_ (.A1(\temp_real[0] ),
    .A2(_08644_),
    .ZN(_05887_));
 OAI21_X2 _15660_ (.A(_05869_),
    .B1(net474),
    .B2(_07358_),
    .ZN(_05888_));
 AOI21_X2 _15661_ (.A(_08703_),
    .B1(_05888_),
    .B2(_05838_),
    .ZN(_05889_));
 OAI21_X2 _15662_ (.A(_05868_),
    .B1(_05889_),
    .B2(_08697_),
    .ZN(_05890_));
 AOI21_X4 _15663_ (.A(_08693_),
    .B1(_05890_),
    .B2(_05829_),
    .ZN(_05891_));
 OAI21_X4 _15664_ (.A(_05867_),
    .B1(_05891_),
    .B2(_08687_),
    .ZN(_05892_));
 AOI21_X4 _15665_ (.A(_08683_),
    .B1(_05892_),
    .B2(_05827_),
    .ZN(_05893_));
 OAI21_X4 _15666_ (.A(_05866_),
    .B1(_05893_),
    .B2(_08677_),
    .ZN(_05894_));
 AOI21_X4 _15667_ (.A(_08673_),
    .B1(_05894_),
    .B2(_05825_),
    .ZN(_05895_));
 OAI21_X2 _15668_ (.A(_05865_),
    .B1(_05895_),
    .B2(_08667_),
    .ZN(_05896_));
 AOI21_X4 _15669_ (.A(_08663_),
    .B1(_05823_),
    .B2(_05896_),
    .ZN(_05897_));
 OAI21_X2 _15670_ (.A(_05864_),
    .B1(_05897_),
    .B2(_08657_),
    .ZN(_05898_));
 AOI21_X2 _15671_ (.A(_08653_),
    .B1(_05882_),
    .B2(_05898_),
    .ZN(_05899_));
 XOR2_X2 _15672_ (.A(_08636_),
    .B(_05899_),
    .Z(_05900_));
 XNOR2_X2 _15673_ (.A(_05881_),
    .B(_05822_),
    .ZN(_05901_));
 XNOR2_X2 _15674_ (.A(_08662_),
    .B(_05879_),
    .ZN(_05902_));
 INV_X1 _15675_ (.A(_08657_),
    .ZN(_05903_));
 XNOR2_X2 _15676_ (.A(_05903_),
    .B(_05897_),
    .ZN(_05904_));
 INV_X1 _15677_ (.A(_08667_),
    .ZN(_05905_));
 XNOR2_X2 _15678_ (.A(_05895_),
    .B(_05905_),
    .ZN(_05906_));
 XNOR2_X2 _15679_ (.A(_08672_),
    .B(net454),
    .ZN(_05907_));
 INV_X1 _15680_ (.A(_08677_),
    .ZN(_05908_));
 XNOR2_X2 _15681_ (.A(_05908_),
    .B(net449),
    .ZN(_05909_));
 XNOR2_X2 _15682_ (.A(_08692_),
    .B(_05873_),
    .ZN(_05910_));
 INV_X1 _15683_ (.A(_08687_),
    .ZN(_05911_));
 XNOR2_X2 _15684_ (.A(_05911_),
    .B(net450),
    .ZN(_05912_));
 XNOR2_X1 _15685_ (.A(net447),
    .B(net457),
    .ZN(_05913_));
 INV_X2 _15686_ (.A(_08639_),
    .ZN(_05914_));
 NOR2_X1 _15687_ (.A1(_07359_),
    .A2(_05914_),
    .ZN(_05915_));
 INV_X1 _15688_ (.A(_08697_),
    .ZN(_05916_));
 XNOR2_X2 _15689_ (.A(_05916_),
    .B(net451),
    .ZN(_05917_));
 XNOR2_X2 _15690_ (.A(net444),
    .B(net455),
    .ZN(_05918_));
 NOR2_X2 _15691_ (.A1(_05917_),
    .A2(_05918_),
    .ZN(_05919_));
 NAND3_X1 _15692_ (.A1(_05913_),
    .A2(_05915_),
    .A3(_05919_),
    .ZN(_05920_));
 XNOR2_X2 _15693_ (.A(_08682_),
    .B(_05875_),
    .ZN(_05921_));
 OR4_X2 _15694_ (.A1(_05910_),
    .A2(_05912_),
    .A3(_05921_),
    .A4(_05920_),
    .ZN(_05922_));
 OR4_X4 _15695_ (.A1(_05922_),
    .A2(_05907_),
    .A3(_05909_),
    .A4(_05906_),
    .ZN(_05923_));
 OR4_X4 _15696_ (.A1(_05923_),
    .A2(_05902_),
    .A3(_05904_),
    .A4(_05901_),
    .ZN(_05924_));
 OAI211_X4 _15697_ (.A(_05886_),
    .B(_05887_),
    .C1(_05924_),
    .C2(_05900_),
    .ZN(_05925_));
 AND2_X4 _15698_ (.A1(_05302_),
    .A2(_05925_),
    .ZN(_05926_));
 BUF_X8 clone59 (.A(_00873_),
    .Z(net59));
 NOR2_X4 _15700_ (.A1(_05925_),
    .A2(_05341_),
    .ZN(_05928_));
 NOR2_X4 _15701_ (.A1(_05928_),
    .A2(_05926_),
    .ZN(_05929_));
 MUX2_X2 _15702_ (.A(_05347_),
    .B(_05356_),
    .S(net453),
    .Z(_05930_));
 BUF_X8 clone97 (.A(_05930_),
    .Z(net97));
 AND3_X4 _15704_ (.A1(_05423_),
    .A2(_05862_),
    .A3(_05930_),
    .ZN(_05932_));
 BUF_X8 _15705_ (.A(_05932_),
    .Z(_05933_));
 NAND2_X1 _15706_ (.A1(\samples_real[0][0] ),
    .A2(net98),
    .ZN(_05934_));
 BUF_X8 _15707_ (.A(net443),
    .Z(_05935_));
 BUF_X16 _15708_ (.A(_05929_),
    .Z(_05936_));
 BUF_X32 _15709_ (.A(_05936_),
    .Z(_05937_));
 AOI22_X4 _15710_ (.A1(_05914_),
    .A2(_05935_),
    .B1(net491),
    .B2(net70),
    .ZN(_05938_));
 NAND2_X1 _15711_ (.A1(net70),
    .A2(_05494_),
    .ZN(_05939_));
 BUF_X4 _15712_ (.A(_05930_),
    .Z(_05940_));
 MUX2_X1 _15713_ (.A(_05938_),
    .B(_05939_),
    .S(net97),
    .Z(_05941_));
 CLKBUF_X3 _15714_ (.A(_05860_),
    .Z(_05942_));
 NAND2_X4 _15715_ (.A1(_05914_),
    .A2(net478),
    .ZN(_05943_));
 OAI221_X1 _15716_ (.A(_05934_),
    .B1(_05941_),
    .B2(_05942_),
    .C1(_05552_),
    .C2(_05943_),
    .ZN(_00453_));
 NAND2_X1 _15717_ (.A1(\samples_real[0][10] ),
    .A2(net98),
    .ZN(_05944_));
 AOI22_X4 _15718_ (.A1(net456),
    .A2(_05935_),
    .B1(net491),
    .B2(net71),
    .ZN(_05945_));
 NAND2_X1 _15719_ (.A1(net71),
    .A2(_05494_),
    .ZN(_05946_));
 MUX2_X1 _15720_ (.A(_05945_),
    .B(_05946_),
    .S(_05940_),
    .Z(_05947_));
 CLKBUF_X3 _15721_ (.A(_05858_),
    .Z(_05948_));
 INV_X1 _15722_ (.A(_08671_),
    .ZN(_05949_));
 INV_X1 _15723_ (.A(_08681_),
    .ZN(_05950_));
 INV_X1 _15724_ (.A(_08691_),
    .ZN(_05951_));
 INV_X1 _15725_ (.A(net446),
    .ZN(_05952_));
 NOR2_X2 _15726_ (.A1(_05952_),
    .A2(_07361_),
    .ZN(_05953_));
 OAI21_X1 _15727_ (.A(net444),
    .B1(_08706_),
    .B2(_05953_),
    .ZN(_05954_));
 AOI21_X1 _15728_ (.A(_05916_),
    .B1(_05831_),
    .B2(_05954_),
    .ZN(_05955_));
 OAI21_X1 _15729_ (.A(_08692_),
    .B1(_08696_),
    .B2(_05955_),
    .ZN(_05956_));
 AOI21_X1 _15730_ (.A(_05911_),
    .B1(_05951_),
    .B2(_05956_),
    .ZN(_05957_));
 OAI21_X1 _15731_ (.A(_08682_),
    .B1(_08686_),
    .B2(_05957_),
    .ZN(_05958_));
 AOI21_X1 _15732_ (.A(_05908_),
    .B1(_05950_),
    .B2(_05958_),
    .ZN(_05959_));
 OAI21_X1 _15733_ (.A(_08672_),
    .B1(_08676_),
    .B2(_05959_),
    .ZN(_05960_));
 AND3_X1 _15734_ (.A1(_05905_),
    .A2(_05949_),
    .A3(_05960_),
    .ZN(_05961_));
 AOI21_X1 _15735_ (.A(_05905_),
    .B1(_05949_),
    .B2(_05960_),
    .ZN(_05962_));
 OR3_X1 _15736_ (.A1(_05948_),
    .A2(_05961_),
    .A3(_05962_),
    .ZN(_05963_));
 CLKBUF_X3 _15737_ (.A(_05963_),
    .Z(_05964_));
 OAI221_X1 _15738_ (.A(_05944_),
    .B1(_05947_),
    .B2(_05942_),
    .C1(_05552_),
    .C2(_05964_),
    .ZN(_00454_));
 NAND2_X1 _15739_ (.A1(\samples_real[0][11] ),
    .A2(net98),
    .ZN(_05965_));
 AOI22_X4 _15740_ (.A1(_05902_),
    .A2(_05935_),
    .B1(_05937_),
    .B2(net72),
    .ZN(_05966_));
 CLKBUF_X3 _15741_ (.A(_05433_),
    .Z(_05967_));
 NAND2_X1 _15742_ (.A1(net72),
    .A2(_05967_),
    .ZN(_05968_));
 MUX2_X1 _15743_ (.A(_05966_),
    .B(_05968_),
    .S(_05940_),
    .Z(_05969_));
 AND3_X1 _15744_ (.A1(_05823_),
    .A2(_05824_),
    .A3(_05846_),
    .ZN(_05970_));
 OR3_X1 _15745_ (.A1(_05847_),
    .A2(_05948_),
    .A3(_05970_),
    .ZN(_05971_));
 BUF_X4 _15746_ (.A(_05971_),
    .Z(_05972_));
 OAI221_X1 _15747_ (.A(_05965_),
    .B1(_05942_),
    .B2(_05969_),
    .C1(_05552_),
    .C2(_05972_),
    .ZN(_00455_));
 NAND2_X1 _15748_ (.A1(\samples_real[0][12] ),
    .A2(_05933_),
    .ZN(_05973_));
 AOI22_X4 _15749_ (.A1(_05904_),
    .A2(_05935_),
    .B1(_05937_),
    .B2(net73),
    .ZN(_05974_));
 NAND2_X1 _15750_ (.A1(net73),
    .A2(_05967_),
    .ZN(_05975_));
 MUX2_X1 _15751_ (.A(_05974_),
    .B(_05975_),
    .S(_05940_),
    .Z(_05976_));
 INV_X1 _15752_ (.A(_08661_),
    .ZN(_05977_));
 OAI21_X1 _15753_ (.A(_08662_),
    .B1(_08666_),
    .B2(_05962_),
    .ZN(_05978_));
 AND3_X1 _15754_ (.A1(_05903_),
    .A2(_05977_),
    .A3(_05978_),
    .ZN(_05979_));
 AOI21_X1 _15755_ (.A(_05903_),
    .B1(_05977_),
    .B2(_05978_),
    .ZN(_05980_));
 OR3_X1 _15756_ (.A1(_05948_),
    .A2(_05979_),
    .A3(_05980_),
    .ZN(_05981_));
 CLKBUF_X3 _15757_ (.A(_05981_),
    .Z(_05982_));
 OAI221_X1 _15758_ (.A(_05973_),
    .B1(_05976_),
    .B2(_05942_),
    .C1(_05552_),
    .C2(_05982_),
    .ZN(_00456_));
 NAND2_X1 _15759_ (.A1(\samples_real[0][13] ),
    .A2(_05933_),
    .ZN(_05983_));
 AOI22_X4 _15760_ (.A1(net464),
    .A2(_05935_),
    .B1(net491),
    .B2(net74),
    .ZN(_05984_));
 NAND2_X1 _15761_ (.A1(net74),
    .A2(_05967_),
    .ZN(_05985_));
 MUX2_X1 _15762_ (.A(_05984_),
    .B(_05985_),
    .S(net97),
    .Z(_05986_));
 OR3_X2 _15763_ (.A1(_05822_),
    .A2(_08656_),
    .A3(_05849_),
    .ZN(_05987_));
 NAND3_X4 _15764_ (.A1(_05850_),
    .A2(net478),
    .A3(_05987_),
    .ZN(_05988_));
 OAI221_X1 _15765_ (.A(_05983_),
    .B1(_05986_),
    .B2(_05942_),
    .C1(_05552_),
    .C2(_05988_),
    .ZN(_00457_));
 NAND2_X1 _15766_ (.A1(\samples_real[0][14] ),
    .A2(_05933_),
    .ZN(_05989_));
 AOI22_X4 _15767_ (.A1(net459),
    .A2(_05935_),
    .B1(net491),
    .B2(net75),
    .ZN(_05990_));
 NAND2_X1 _15768_ (.A1(net75),
    .A2(_05967_),
    .ZN(_05991_));
 MUX2_X1 _15769_ (.A(_05990_),
    .B(_05991_),
    .S(_05940_),
    .Z(_05992_));
 OAI21_X1 _15770_ (.A(_05822_),
    .B1(_08656_),
    .B2(_05980_),
    .ZN(_05993_));
 NAND2_X1 _15771_ (.A1(_05821_),
    .A2(_05993_),
    .ZN(_05994_));
 XOR2_X2 _15772_ (.A(_08647_),
    .B(_05994_),
    .Z(_05995_));
 NAND2_X4 _15773_ (.A1(net478),
    .A2(_05995_),
    .ZN(_05996_));
 OAI221_X1 _15774_ (.A(_05989_),
    .B1(_05992_),
    .B2(_05942_),
    .C1(_05552_),
    .C2(_05996_),
    .ZN(_00458_));
 INV_X1 _15775_ (.A(net76),
    .ZN(_05997_));
 AOI22_X4 _15776_ (.A1(net463),
    .A2(_05926_),
    .B1(_05936_),
    .B2(_05997_),
    .ZN(_05998_));
 NOR2_X4 _15777_ (.A1(net97),
    .A2(_05998_),
    .ZN(_05999_));
 AOI22_X1 _15778_ (.A1(net76),
    .A2(_05434_),
    .B1(_05423_),
    .B2(\samples_real[0][15] ),
    .ZN(_06000_));
 AOI21_X2 _15779_ (.A(_05999_),
    .B1(_06000_),
    .B2(net97),
    .ZN(_06001_));
 OR2_X2 _15780_ (.A1(_05358_),
    .A2(_05854_),
    .ZN(_06002_));
 MUX2_X1 _15781_ (.A(_06001_),
    .B(_06002_),
    .S(_05860_),
    .Z(_00459_));
 NAND2_X1 _15782_ (.A1(\samples_real[0][1] ),
    .A2(_05933_),
    .ZN(_06003_));
 AOI22_X4 _15783_ (.A1(_07359_),
    .A2(_05935_),
    .B1(_05937_),
    .B2(net77),
    .ZN(_06004_));
 NAND2_X1 _15784_ (.A1(net77),
    .A2(_05967_),
    .ZN(_06005_));
 MUX2_X1 _15785_ (.A(_06004_),
    .B(_06005_),
    .S(_05940_),
    .Z(_06006_));
 NAND2_X4 _15786_ (.A1(_07362_),
    .A2(net478),
    .ZN(_06007_));
 OAI221_X1 _15787_ (.A(_06003_),
    .B1(_06006_),
    .B2(_05942_),
    .C1(_05552_),
    .C2(_06007_),
    .ZN(_00460_));
 AND2_X1 _15788_ (.A1(_05952_),
    .A2(_07361_),
    .ZN(_06008_));
 NOR3_X4 _15789_ (.A1(_05948_),
    .A2(_05953_),
    .A3(_06008_),
    .ZN(_06009_));
 NAND2_X1 _15790_ (.A1(_05942_),
    .A2(_06009_),
    .ZN(_06010_));
 INV_X1 _15791_ (.A(_05913_),
    .ZN(_06011_));
 AOI22_X4 _15792_ (.A1(_06011_),
    .A2(_05935_),
    .B1(_05937_),
    .B2(net78),
    .ZN(_06012_));
 AOI22_X1 _15793_ (.A1(net78),
    .A2(_05434_),
    .B1(_05423_),
    .B2(\samples_real[0][2] ),
    .ZN(_06013_));
 MUX2_X1 _15794_ (.A(_06012_),
    .B(_06013_),
    .S(net97),
    .Z(_06014_));
 OAI21_X2 _15795_ (.A(_06010_),
    .B1(_06014_),
    .B2(_05942_),
    .ZN(_00461_));
 NAND2_X4 _15796_ (.A1(_05933_),
    .A2(\samples_real[0][3] ),
    .ZN(_06015_));
 AOI22_X4 _15797_ (.A1(_05918_),
    .A2(_05935_),
    .B1(net491),
    .B2(net79),
    .ZN(_06016_));
 NAND2_X1 _15798_ (.A1(net79),
    .A2(_05967_),
    .ZN(_06017_));
 MUX2_X1 _15799_ (.A(_06016_),
    .B(_06017_),
    .S(_05930_),
    .Z(_06018_));
 XNOR2_X2 _15800_ (.A(net445),
    .B(_05836_),
    .ZN(_06019_));
 NAND2_X4 _15801_ (.A1(net478),
    .A2(_06019_),
    .ZN(_06020_));
 OAI221_X2 _15802_ (.A(_06015_),
    .B1(_06018_),
    .B2(_05942_),
    .C1(_05440_),
    .C2(_06020_),
    .ZN(_00462_));
 NAND2_X4 _15803_ (.A1(net98),
    .A2(\samples_real[0][4] ),
    .ZN(_06021_));
 AOI22_X4 _15804_ (.A1(_05917_),
    .A2(_05935_),
    .B1(_05937_),
    .B2(net80),
    .ZN(_06022_));
 NAND2_X1 _15805_ (.A1(net80),
    .A2(_05967_),
    .ZN(_06023_));
 MUX2_X1 _15806_ (.A(_06022_),
    .B(_06023_),
    .S(net94),
    .Z(_06024_));
 AND3_X1 _15807_ (.A1(_05916_),
    .A2(_05831_),
    .A3(_05954_),
    .ZN(_06025_));
 OR3_X1 _15808_ (.A1(_05948_),
    .A2(_05955_),
    .A3(_06025_),
    .ZN(_06026_));
 CLKBUF_X3 _15809_ (.A(_06026_),
    .Z(_06027_));
 OAI221_X2 _15810_ (.A(_06021_),
    .B1(_06024_),
    .B2(net470),
    .C1(_05440_),
    .C2(_06027_),
    .ZN(_00463_));
 NAND2_X4 _15811_ (.A1(net98),
    .A2(\samples_real[0][5] ),
    .ZN(_06028_));
 AOI22_X4 _15812_ (.A1(_05910_),
    .A2(net443),
    .B1(net58),
    .B2(net81),
    .ZN(_06029_));
 NAND2_X1 _15813_ (.A1(net81),
    .A2(_05967_),
    .ZN(_06030_));
 MUX2_X1 _15814_ (.A(_06029_),
    .B(_06030_),
    .S(net94),
    .Z(_06031_));
 AND3_X1 _15815_ (.A1(_05829_),
    .A2(_05830_),
    .A3(_05840_),
    .ZN(_06032_));
 OR3_X1 _15816_ (.A1(_05841_),
    .A2(_05948_),
    .A3(_06032_),
    .ZN(_06033_));
 BUF_X4 _15817_ (.A(_06033_),
    .Z(_06034_));
 OAI221_X2 _15818_ (.A(_06028_),
    .B1(_06031_),
    .B2(net470),
    .C1(_05440_),
    .C2(_06034_),
    .ZN(_00464_));
 NAND2_X4 _15819_ (.A1(_05932_),
    .A2(\samples_real[0][6] ),
    .ZN(_06035_));
 AOI22_X4 _15820_ (.A1(_05912_),
    .A2(net443),
    .B1(net58),
    .B2(net82),
    .ZN(_06036_));
 NAND2_X1 _15821_ (.A1(net82),
    .A2(_05967_),
    .ZN(_06037_));
 MUX2_X1 _15822_ (.A(_06036_),
    .B(_06037_),
    .S(net94),
    .Z(_06038_));
 AND3_X1 _15823_ (.A1(_05911_),
    .A2(_05951_),
    .A3(_05956_),
    .ZN(_06039_));
 OR3_X1 _15824_ (.A1(_05948_),
    .A2(_05957_),
    .A3(_06039_),
    .ZN(_06040_));
 BUF_X4 _15825_ (.A(_06040_),
    .Z(_06041_));
 OAI221_X2 _15826_ (.A(_06035_),
    .B1(_06038_),
    .B2(_05860_),
    .C1(_05440_),
    .C2(_06041_),
    .ZN(_00465_));
 NAND2_X4 _15827_ (.A1(_05932_),
    .A2(\samples_real[0][7] ),
    .ZN(_06042_));
 AOI22_X4 _15828_ (.A1(net462),
    .A2(net443),
    .B1(net58),
    .B2(net83),
    .ZN(_06043_));
 NAND2_X1 _15829_ (.A1(net83),
    .A2(_05967_),
    .ZN(_06044_));
 MUX2_X1 _15830_ (.A(_06043_),
    .B(_06044_),
    .S(net94),
    .Z(_06045_));
 AND3_X1 _15831_ (.A1(_05827_),
    .A2(_05828_),
    .A3(_05842_),
    .ZN(_06046_));
 OR3_X1 _15832_ (.A1(_05843_),
    .A2(_05948_),
    .A3(_06046_),
    .ZN(_06047_));
 BUF_X4 _15833_ (.A(_06047_),
    .Z(_06048_));
 OAI221_X2 _15834_ (.A(_06042_),
    .B1(_06045_),
    .B2(_05860_),
    .C1(_05440_),
    .C2(_06048_),
    .ZN(_00466_));
 NAND2_X1 _15835_ (.A1(\samples_real[0][8] ),
    .A2(_05932_),
    .ZN(_06049_));
 AOI22_X4 _15836_ (.A1(_05909_),
    .A2(net460),
    .B1(net58),
    .B2(net84),
    .ZN(_06050_));
 NAND2_X1 _15837_ (.A1(net84),
    .A2(_05433_),
    .ZN(_06051_));
 MUX2_X1 _15838_ (.A(_06050_),
    .B(_06051_),
    .S(net461),
    .Z(_06052_));
 AND3_X1 _15839_ (.A1(_05908_),
    .A2(_05950_),
    .A3(_05958_),
    .ZN(_06053_));
 OR3_X1 _15840_ (.A1(_05948_),
    .A2(_05959_),
    .A3(_06053_),
    .ZN(_06054_));
 BUF_X4 _15841_ (.A(_06054_),
    .Z(_06055_));
 OAI221_X1 _15842_ (.A(_06049_),
    .B1(_06052_),
    .B2(net470),
    .C1(_05440_),
    .C2(_06055_),
    .ZN(_00467_));
 NAND2_X1 _15843_ (.A1(\samples_real[0][9] ),
    .A2(_05932_),
    .ZN(_06056_));
 AOI22_X4 _15844_ (.A1(_05907_),
    .A2(_05926_),
    .B1(net58),
    .B2(net85),
    .ZN(_06057_));
 NAND2_X1 _15845_ (.A1(net85),
    .A2(_05433_),
    .ZN(_06058_));
 MUX2_X1 _15846_ (.A(_06057_),
    .B(_06058_),
    .S(net461),
    .Z(_06059_));
 AND3_X1 _15847_ (.A1(_05825_),
    .A2(_05826_),
    .A3(_05844_),
    .ZN(_06060_));
 OR3_X1 _15848_ (.A1(_05845_),
    .A2(_05948_),
    .A3(_06060_),
    .ZN(_06061_));
 BUF_X4 _15849_ (.A(_06061_),
    .Z(_06062_));
 OAI221_X1 _15850_ (.A(_06056_),
    .B1(_06059_),
    .B2(net470),
    .C1(_05440_),
    .C2(_06062_),
    .ZN(_00468_));
 MUX2_X2 _15851_ (.A(_05573_),
    .B(_05576_),
    .S(_05936_),
    .Z(_06063_));
 NAND3_X4 _15852_ (.A1(_04790_),
    .A2(_05297_),
    .A3(_05859_),
    .ZN(_06064_));
 AND3_X4 _15853_ (.A1(_06063_),
    .A2(_05571_),
    .A3(_06064_),
    .ZN(_06065_));
 BUF_X8 _15854_ (.A(_06065_),
    .Z(_06066_));
 NAND2_X4 _15855_ (.A1(\samples_real[1][0] ),
    .A2(net482),
    .ZN(_06067_));
 INV_X4 _15856_ (.A(_06063_),
    .ZN(_06068_));
 NAND2_X4 _15857_ (.A1(_06068_),
    .A2(_06064_),
    .ZN(_06069_));
 BUF_X8 _15858_ (.A(_06069_),
    .Z(_06070_));
 CLKBUF_X3 _15859_ (.A(_05582_),
    .Z(_06071_));
 OAI221_X2 _15860_ (.A(_06067_),
    .B1(_06070_),
    .B2(_05938_),
    .C1(_06071_),
    .C2(_05943_),
    .ZN(_00469_));
 NAND2_X4 _15861_ (.A1(\samples_real[1][10] ),
    .A2(_06066_),
    .ZN(_06072_));
 OAI221_X2 _15862_ (.A(_06072_),
    .B1(_06070_),
    .B2(_05945_),
    .C1(_06071_),
    .C2(_05964_),
    .ZN(_00470_));
 NAND2_X2 _15863_ (.A1(\samples_real[1][11] ),
    .A2(_06066_),
    .ZN(_06073_));
 OAI221_X1 _15864_ (.A(_06073_),
    .B1(_06070_),
    .B2(_05966_),
    .C1(_06071_),
    .C2(_05972_),
    .ZN(_00471_));
 NAND2_X4 _15865_ (.A1(_06066_),
    .A2(\samples_real[1][12] ),
    .ZN(_06074_));
 OAI221_X2 _15866_ (.A(_06074_),
    .B1(_06070_),
    .B2(_05974_),
    .C1(_06071_),
    .C2(_05982_),
    .ZN(_00472_));
 NAND2_X4 _15867_ (.A1(net482),
    .A2(\samples_real[1][13] ),
    .ZN(_06075_));
 OAI221_X2 _15868_ (.A(_06075_),
    .B1(_06070_),
    .B2(_05984_),
    .C1(_06071_),
    .C2(_05988_),
    .ZN(_00473_));
 NAND2_X4 _15869_ (.A1(\samples_real[1][14] ),
    .A2(net482),
    .ZN(_06076_));
 OAI221_X2 _15870_ (.A(_06076_),
    .B1(_06070_),
    .B2(_05990_),
    .C1(_06071_),
    .C2(_05996_),
    .ZN(_00474_));
 NAND2_X4 _15871_ (.A1(_05998_),
    .A2(_06068_),
    .ZN(_06077_));
 NAND3_X2 _15872_ (.A1(_06063_),
    .A2(\samples_real[1][15] ),
    .A3(_05672_),
    .ZN(_06078_));
 NAND2_X2 _15873_ (.A1(_06077_),
    .A2(_06078_),
    .ZN(_06079_));
 MUX2_X1 _15874_ (.A(_06002_),
    .B(_06079_),
    .S(_06064_),
    .Z(_00475_));
 NAND2_X4 _15875_ (.A1(net482),
    .A2(\samples_real[1][1] ),
    .ZN(_06080_));
 OAI221_X2 _15876_ (.A(_06080_),
    .B1(_06070_),
    .B2(_06004_),
    .C1(_06071_),
    .C2(_06007_),
    .ZN(_00476_));
 NAND3_X2 _15877_ (.A1(_06063_),
    .A2(_00855_),
    .A3(\samples_real[1][2] ),
    .ZN(_06081_));
 OAI21_X2 _15878_ (.A(_06081_),
    .B1(_06012_),
    .B2(_06063_),
    .ZN(_06082_));
 MUX2_X1 _15879_ (.A(_06009_),
    .B(_06082_),
    .S(_06064_),
    .Z(_00477_));
 NAND2_X4 _15880_ (.A1(net482),
    .A2(\samples_real[1][3] ),
    .ZN(_06083_));
 OAI221_X2 _15881_ (.A(_06083_),
    .B1(_06070_),
    .B2(_06016_),
    .C1(_06071_),
    .C2(_06020_),
    .ZN(_00478_));
 NAND2_X4 _15882_ (.A1(_06066_),
    .A2(\samples_real[1][4] ),
    .ZN(_06084_));
 OAI221_X2 _15883_ (.A(_06084_),
    .B1(_06070_),
    .B2(_06022_),
    .C1(_06071_),
    .C2(_06027_),
    .ZN(_00479_));
 NAND2_X4 _15884_ (.A1(_06066_),
    .A2(\samples_real[1][5] ),
    .ZN(_06085_));
 OAI221_X2 _15885_ (.A(_06085_),
    .B1(_06070_),
    .B2(_06029_),
    .C1(_06071_),
    .C2(_06034_),
    .ZN(_00480_));
 NAND2_X4 _15886_ (.A1(net486),
    .A2(\samples_real[1][6] ),
    .ZN(_06086_));
 OAI221_X2 _15887_ (.A(_06086_),
    .B1(_06069_),
    .B2(_06036_),
    .C1(_05583_),
    .C2(_06041_),
    .ZN(_00481_));
 NAND2_X2 _15888_ (.A1(_06065_),
    .A2(\samples_real[1][7] ),
    .ZN(_06087_));
 OAI221_X1 _15889_ (.A(_06087_),
    .B1(_06069_),
    .B2(_06043_),
    .C1(_05583_),
    .C2(_06048_),
    .ZN(_00482_));
 NAND2_X4 _15890_ (.A1(net486),
    .A2(\samples_real[1][8] ),
    .ZN(_06088_));
 OAI221_X2 _15891_ (.A(_06088_),
    .B1(_06069_),
    .B2(_06050_),
    .C1(_05583_),
    .C2(_06055_),
    .ZN(_00483_));
 NAND2_X4 _15892_ (.A1(net486),
    .A2(\samples_real[1][9] ),
    .ZN(_06089_));
 OAI221_X2 _15893_ (.A(_06089_),
    .B1(_06069_),
    .B2(_06057_),
    .C1(_05583_),
    .C2(_06062_),
    .ZN(_00484_));
 MUX2_X2 _15894_ (.A(_05614_),
    .B(_05615_),
    .S(_05936_),
    .Z(_06090_));
 NAND2_X2 _15895_ (.A1(_05620_),
    .A2(_05859_),
    .ZN(_06091_));
 AND3_X4 _15896_ (.A1(_06090_),
    .A2(_05571_),
    .A3(_06091_),
    .ZN(_06092_));
 BUF_X8 _15897_ (.A(_06092_),
    .Z(_06093_));
 NAND2_X4 _15898_ (.A1(\samples_real[2][0] ),
    .A2(net483),
    .ZN(_06094_));
 INV_X4 _15899_ (.A(_06090_),
    .ZN(_06095_));
 NAND2_X4 _15900_ (.A1(_06095_),
    .A2(_06091_),
    .ZN(_06096_));
 BUF_X4 _15901_ (.A(_06096_),
    .Z(_06097_));
 BUF_X2 _15902_ (.A(_05626_),
    .Z(_06098_));
 OAI221_X2 _15903_ (.A(_06094_),
    .B1(_06097_),
    .B2(_05938_),
    .C1(_06098_),
    .C2(_05943_),
    .ZN(_00485_));
 NAND2_X4 _15904_ (.A1(\samples_real[2][10] ),
    .A2(net483),
    .ZN(_06099_));
 OAI221_X2 _15905_ (.A(_06099_),
    .B1(_06097_),
    .B2(_05945_),
    .C1(_06098_),
    .C2(_05964_),
    .ZN(_00486_));
 NAND2_X4 _15906_ (.A1(\samples_real[2][11] ),
    .A2(_06093_),
    .ZN(_06100_));
 OAI221_X2 _15907_ (.A(_06100_),
    .B1(_06097_),
    .B2(_05966_),
    .C1(_06098_),
    .C2(_05972_),
    .ZN(_00487_));
 NAND2_X2 _15908_ (.A1(\samples_real[2][12] ),
    .A2(_06093_),
    .ZN(_06101_));
 OAI221_X1 _15909_ (.A(_06101_),
    .B1(_06097_),
    .B2(_05974_),
    .C1(_06098_),
    .C2(_05982_),
    .ZN(_00488_));
 NAND2_X2 _15910_ (.A1(\samples_real[2][13] ),
    .A2(_06093_),
    .ZN(_06102_));
 OAI221_X1 _15911_ (.A(_06102_),
    .B1(_06097_),
    .B2(_05984_),
    .C1(_06098_),
    .C2(_05988_),
    .ZN(_00489_));
 NAND2_X4 _15912_ (.A1(\samples_real[2][14] ),
    .A2(_06093_),
    .ZN(_06103_));
 OAI221_X2 _15913_ (.A(_06103_),
    .B1(_06097_),
    .B2(_05990_),
    .C1(_06098_),
    .C2(_05996_),
    .ZN(_00490_));
 NAND2_X2 _15914_ (.A1(_05998_),
    .A2(_06095_),
    .ZN(_06104_));
 NAND3_X2 _15915_ (.A1(_06090_),
    .A2(\samples_real[2][15] ),
    .A3(_05672_),
    .ZN(_06105_));
 NAND2_X1 _15916_ (.A1(_06104_),
    .A2(_06105_),
    .ZN(_06106_));
 MUX2_X1 _15917_ (.A(_06002_),
    .B(_06106_),
    .S(_06091_),
    .Z(_00491_));
 NAND2_X1 _15918_ (.A1(\samples_real[2][1] ),
    .A2(_06093_),
    .ZN(_06107_));
 OAI221_X1 _15919_ (.A(_06107_),
    .B1(_06097_),
    .B2(_06004_),
    .C1(_06098_),
    .C2(_06007_),
    .ZN(_00492_));
 NAND3_X2 _15920_ (.A1(_06090_),
    .A2(\samples_real[2][2] ),
    .A3(_00855_),
    .ZN(_06108_));
 OAI21_X2 _15921_ (.A(_06108_),
    .B1(_06012_),
    .B2(_06090_),
    .ZN(_06109_));
 MUX2_X1 _15922_ (.A(_06009_),
    .B(_06109_),
    .S(_06091_),
    .Z(_00493_));
 NAND2_X2 _15923_ (.A1(\samples_real[2][3] ),
    .A2(net483),
    .ZN(_06110_));
 OAI221_X1 _15924_ (.A(_06110_),
    .B1(_06097_),
    .B2(_06016_),
    .C1(_06098_),
    .C2(_06020_),
    .ZN(_00494_));
 NAND2_X4 _15925_ (.A1(net483),
    .A2(\samples_real[2][4] ),
    .ZN(_06111_));
 OAI221_X2 _15926_ (.A(_06111_),
    .B1(_06097_),
    .B2(_06022_),
    .C1(_06098_),
    .C2(_06027_),
    .ZN(_00495_));
 NAND2_X4 _15927_ (.A1(\samples_real[2][5] ),
    .A2(net483),
    .ZN(_06112_));
 OAI221_X2 _15928_ (.A(_06112_),
    .B1(_06097_),
    .B2(_06029_),
    .C1(_06098_),
    .C2(_06034_),
    .ZN(_00496_));
 NAND2_X4 _15929_ (.A1(_06092_),
    .A2(\samples_real[2][6] ),
    .ZN(_06113_));
 OAI221_X2 _15930_ (.A(_06113_),
    .B1(_06096_),
    .B2(_06036_),
    .C1(_05627_),
    .C2(_06041_),
    .ZN(_00497_));
 NAND2_X4 _15931_ (.A1(net524),
    .A2(\samples_real[2][7] ),
    .ZN(_06114_));
 OAI221_X2 _15932_ (.A(_06114_),
    .B1(_06096_),
    .B2(_06043_),
    .C1(_05627_),
    .C2(_06048_),
    .ZN(_00498_));
 NAND2_X4 _15933_ (.A1(net524),
    .A2(\samples_real[2][8] ),
    .ZN(_06115_));
 OAI221_X2 _15934_ (.A(_06115_),
    .B1(_06096_),
    .B2(_06050_),
    .C1(_05627_),
    .C2(_06055_),
    .ZN(_00499_));
 NAND2_X2 _15935_ (.A1(_06092_),
    .A2(\samples_real[2][9] ),
    .ZN(_06116_));
 OAI221_X1 _15936_ (.A(_06116_),
    .B1(_06096_),
    .B2(_06057_),
    .C1(_05627_),
    .C2(_06062_),
    .ZN(_00500_));
 MUX2_X2 _15937_ (.A(_05651_),
    .B(_05653_),
    .S(_05936_),
    .Z(_06117_));
 NAND2_X2 _15938_ (.A1(_05655_),
    .A2(_05859_),
    .ZN(_06118_));
 AND3_X4 _15939_ (.A1(_06118_),
    .A2(_05571_),
    .A3(_06117_),
    .ZN(_06119_));
 BUF_X16 _15940_ (.A(_06119_),
    .Z(_06120_));
 NAND2_X4 _15941_ (.A1(\samples_real[3][0] ),
    .A2(net93),
    .ZN(_06121_));
 INV_X4 _15942_ (.A(_06117_),
    .ZN(_06122_));
 NAND2_X2 _15943_ (.A1(_06122_),
    .A2(_06118_),
    .ZN(_06123_));
 BUF_X8 _15944_ (.A(_06123_),
    .Z(_06124_));
 CLKBUF_X3 _15945_ (.A(_05661_),
    .Z(_06125_));
 OAI221_X2 _15946_ (.A(_06121_),
    .B1(_06124_),
    .B2(_05938_),
    .C1(_06125_),
    .C2(_05943_),
    .ZN(_00501_));
 NAND2_X4 _15947_ (.A1(net93),
    .A2(\samples_real[3][10] ),
    .ZN(_06126_));
 OAI221_X2 _15948_ (.A(_06126_),
    .B1(_06124_),
    .B2(_05945_),
    .C1(_06125_),
    .C2(_05964_),
    .ZN(_00502_));
 NAND2_X4 _15949_ (.A1(net93),
    .A2(\samples_real[3][11] ),
    .ZN(_06127_));
 OAI221_X2 _15950_ (.A(_06127_),
    .B1(_06124_),
    .B2(_05966_),
    .C1(_06125_),
    .C2(_05972_),
    .ZN(_00503_));
 NAND2_X4 _15951_ (.A1(net93),
    .A2(\samples_real[3][12] ),
    .ZN(_06128_));
 OAI221_X2 _15952_ (.A(_06128_),
    .B1(_06124_),
    .B2(_05974_),
    .C1(_06125_),
    .C2(_05982_),
    .ZN(_00504_));
 NAND2_X4 _15953_ (.A1(\samples_real[3][13] ),
    .A2(net93),
    .ZN(_06129_));
 OAI221_X2 _15954_ (.A(_06129_),
    .B1(_06124_),
    .B2(_05984_),
    .C1(_06125_),
    .C2(_05988_),
    .ZN(_00505_));
 NAND2_X4 _15955_ (.A1(_06120_),
    .A2(\samples_real[3][14] ),
    .ZN(_06130_));
 OAI221_X2 _15956_ (.A(_06130_),
    .B1(_06124_),
    .B2(_05990_),
    .C1(_06125_),
    .C2(_05996_),
    .ZN(_00506_));
 NAND2_X2 _15957_ (.A1(_05998_),
    .A2(_06122_),
    .ZN(_06131_));
 NAND3_X2 _15958_ (.A1(_06117_),
    .A2(\samples_real[3][15] ),
    .A3(_05672_),
    .ZN(_06132_));
 NAND2_X1 _15959_ (.A1(_06131_),
    .A2(_06132_),
    .ZN(_06133_));
 MUX2_X1 _15960_ (.A(_06002_),
    .B(_06133_),
    .S(_06118_),
    .Z(_00507_));
 NAND2_X4 _15961_ (.A1(_06120_),
    .A2(\samples_real[3][1] ),
    .ZN(_06134_));
 OAI221_X2 _15962_ (.A(_06134_),
    .B1(_06124_),
    .B2(_06004_),
    .C1(_06125_),
    .C2(_06007_),
    .ZN(_00508_));
 NAND3_X2 _15963_ (.A1(_06117_),
    .A2(\samples_real[3][2] ),
    .A3(_00855_),
    .ZN(_06135_));
 OAI21_X2 _15964_ (.A(_06135_),
    .B1(_06012_),
    .B2(_06117_),
    .ZN(_06136_));
 MUX2_X1 _15965_ (.A(_06009_),
    .B(_06136_),
    .S(_06118_),
    .Z(_00509_));
 NAND2_X4 _15966_ (.A1(_06120_),
    .A2(\samples_real[3][3] ),
    .ZN(_06137_));
 OAI221_X2 _15967_ (.A(_06137_),
    .B1(_06124_),
    .B2(_06016_),
    .C1(_06125_),
    .C2(_06020_),
    .ZN(_00510_));
 NAND2_X4 _15968_ (.A1(\samples_real[3][4] ),
    .A2(_06120_),
    .ZN(_06138_));
 OAI221_X2 _15969_ (.A(_06138_),
    .B1(_06124_),
    .B2(_06022_),
    .C1(_06125_),
    .C2(_06027_),
    .ZN(_00511_));
 NAND2_X4 _15970_ (.A1(\samples_real[3][5] ),
    .A2(_06120_),
    .ZN(_06139_));
 OAI221_X2 _15971_ (.A(_06139_),
    .B1(_06124_),
    .B2(_06029_),
    .C1(_06125_),
    .C2(_06034_),
    .ZN(_00512_));
 NAND2_X4 _15972_ (.A1(_06119_),
    .A2(\samples_real[3][6] ),
    .ZN(_06140_));
 OAI221_X2 _15973_ (.A(_06140_),
    .B1(_06123_),
    .B2(_06036_),
    .C1(_05662_),
    .C2(_06041_),
    .ZN(_00513_));
 NAND2_X2 _15974_ (.A1(_06119_),
    .A2(\samples_real[3][7] ),
    .ZN(_06141_));
 OAI221_X1 _15975_ (.A(_06141_),
    .B1(_06123_),
    .B2(_06043_),
    .C1(_05662_),
    .C2(_06048_),
    .ZN(_00514_));
 NAND2_X4 _15976_ (.A1(_06119_),
    .A2(\samples_real[3][8] ),
    .ZN(_06142_));
 OAI221_X2 _15977_ (.A(_06142_),
    .B1(_06123_),
    .B2(_06050_),
    .C1(_05662_),
    .C2(_06055_),
    .ZN(_00515_));
 NAND2_X4 _15978_ (.A1(_06119_),
    .A2(\samples_real[3][9] ),
    .ZN(_06143_));
 OAI221_X2 _15979_ (.A(_06143_),
    .B1(_06123_),
    .B2(_06057_),
    .C1(_05662_),
    .C2(_06062_),
    .ZN(_00516_));
 MUX2_X2 _15980_ (.A(_05687_),
    .B(_05689_),
    .S(net453),
    .Z(_06144_));
 NAND2_X2 _15981_ (.A1(_05693_),
    .A2(_05859_),
    .ZN(_06145_));
 AND3_X4 _15982_ (.A1(_06144_),
    .A2(_06145_),
    .A3(_05571_),
    .ZN(_06146_));
 BUF_X16 _15983_ (.A(_06146_),
    .Z(_06147_));
 NAND2_X4 _15984_ (.A1(net101),
    .A2(\samples_real[4][0] ),
    .ZN(_06148_));
 INV_X4 _15985_ (.A(_06144_),
    .ZN(_06149_));
 NAND2_X4 _15986_ (.A1(_06149_),
    .A2(_06145_),
    .ZN(_06150_));
 BUF_X4 _15987_ (.A(_06150_),
    .Z(_06151_));
 BUF_X2 _15988_ (.A(_05692_),
    .Z(_06152_));
 OAI221_X2 _15989_ (.A(_06148_),
    .B1(_06151_),
    .B2(_05938_),
    .C1(_06152_),
    .C2(_05943_),
    .ZN(_00517_));
 NAND2_X4 _15990_ (.A1(net101),
    .A2(\samples_real[4][10] ),
    .ZN(_06153_));
 OAI221_X2 _15991_ (.A(_06153_),
    .B1(_06151_),
    .B2(_05945_),
    .C1(_06152_),
    .C2(_05964_),
    .ZN(_00518_));
 NAND2_X4 _15992_ (.A1(\samples_real[4][11] ),
    .A2(_06147_),
    .ZN(_06154_));
 OAI221_X2 _15993_ (.A(_06154_),
    .B1(_06151_),
    .B2(_05966_),
    .C1(_06152_),
    .C2(_05972_),
    .ZN(_00519_));
 NAND2_X4 _15994_ (.A1(\samples_real[4][12] ),
    .A2(_06147_),
    .ZN(_06155_));
 OAI221_X2 _15995_ (.A(_06155_),
    .B1(_06151_),
    .B2(_05974_),
    .C1(_06152_),
    .C2(_05982_),
    .ZN(_00520_));
 NAND2_X2 _15996_ (.A1(\samples_real[4][13] ),
    .A2(net101),
    .ZN(_06156_));
 OAI221_X1 _15997_ (.A(_06156_),
    .B1(_06151_),
    .B2(_05984_),
    .C1(_06152_),
    .C2(_05988_),
    .ZN(_00521_));
 NAND2_X4 _15998_ (.A1(_06147_),
    .A2(\samples_real[4][14] ),
    .ZN(_06157_));
 OAI221_X2 _15999_ (.A(_06157_),
    .B1(_06151_),
    .B2(_05990_),
    .C1(_06152_),
    .C2(_05996_),
    .ZN(_00522_));
 NAND2_X2 _16000_ (.A1(_05998_),
    .A2(_06149_),
    .ZN(_06158_));
 NAND3_X1 _16001_ (.A1(_05672_),
    .A2(\samples_real[4][15] ),
    .A3(_06144_),
    .ZN(_06159_));
 NAND2_X1 _16002_ (.A1(_06158_),
    .A2(_06159_),
    .ZN(_06160_));
 MUX2_X1 _16003_ (.A(_06002_),
    .B(_06160_),
    .S(_06145_),
    .Z(_00523_));
 NAND2_X4 _16004_ (.A1(_06147_),
    .A2(\samples_real[4][1] ),
    .ZN(_06161_));
 OAI221_X2 _16005_ (.A(_06161_),
    .B1(_06151_),
    .B2(_06004_),
    .C1(_06152_),
    .C2(_06007_),
    .ZN(_00524_));
 NAND3_X2 _16006_ (.A1(_06144_),
    .A2(\samples_real[4][2] ),
    .A3(_00855_),
    .ZN(_06162_));
 OAI21_X2 _16007_ (.A(_06162_),
    .B1(_06012_),
    .B2(net517),
    .ZN(_06163_));
 MUX2_X1 _16008_ (.A(_06009_),
    .B(_06163_),
    .S(_06145_),
    .Z(_00525_));
 NAND2_X4 _16009_ (.A1(net101),
    .A2(\samples_real[4][3] ),
    .ZN(_06164_));
 OAI221_X2 _16010_ (.A(_06164_),
    .B1(_06151_),
    .B2(_06016_),
    .C1(_06152_),
    .C2(_06020_),
    .ZN(_00526_));
 NAND2_X4 _16011_ (.A1(net101),
    .A2(\samples_real[4][4] ),
    .ZN(_06165_));
 OAI221_X2 _16012_ (.A(_06165_),
    .B1(_06151_),
    .B2(_06022_),
    .C1(_06152_),
    .C2(_06027_),
    .ZN(_00527_));
 NAND2_X4 _16013_ (.A1(_06147_),
    .A2(\samples_real[4][5] ),
    .ZN(_06166_));
 OAI221_X2 _16014_ (.A(_06166_),
    .B1(_06151_),
    .B2(_06029_),
    .C1(_06152_),
    .C2(_06034_),
    .ZN(_00528_));
 NAND2_X2 _16015_ (.A1(_06146_),
    .A2(\samples_real[4][6] ),
    .ZN(_06167_));
 OAI221_X1 _16016_ (.A(_06167_),
    .B1(_06150_),
    .B2(_06036_),
    .C1(_05698_),
    .C2(_06041_),
    .ZN(_00529_));
 NAND2_X2 _16017_ (.A1(_06146_),
    .A2(\samples_real[4][7] ),
    .ZN(_06168_));
 OAI221_X1 _16018_ (.A(_06168_),
    .B1(_06150_),
    .B2(_06043_),
    .C1(_05698_),
    .C2(_06048_),
    .ZN(_00530_));
 NAND2_X2 _16019_ (.A1(_06146_),
    .A2(\samples_real[4][8] ),
    .ZN(_06169_));
 OAI221_X1 _16020_ (.A(_06169_),
    .B1(_06150_),
    .B2(_06050_),
    .C1(_05698_),
    .C2(_06055_),
    .ZN(_00531_));
 NAND2_X4 _16021_ (.A1(_06146_),
    .A2(\samples_real[4][9] ),
    .ZN(_06170_));
 OAI221_X2 _16022_ (.A(_06170_),
    .B1(_06150_),
    .B2(_06057_),
    .C1(_05698_),
    .C2(_06062_),
    .ZN(_00532_));
 MUX2_X2 _16023_ (.A(_05721_),
    .B(_05722_),
    .S(net453),
    .Z(_06171_));
 NAND2_X2 _16024_ (.A1(_05725_),
    .A2(_05859_),
    .ZN(_06172_));
 AND3_X4 _16025_ (.A1(_00842_),
    .A2(_06172_),
    .A3(_06171_),
    .ZN(_06173_));
 BUF_X16 _16026_ (.A(_06173_),
    .Z(_06174_));
 NAND2_X4 _16027_ (.A1(net104),
    .A2(\samples_real[5][0] ),
    .ZN(_06175_));
 INV_X4 _16028_ (.A(_06171_),
    .ZN(_06176_));
 NAND2_X4 _16029_ (.A1(_06176_),
    .A2(_06172_),
    .ZN(_06177_));
 BUF_X8 _16030_ (.A(_06177_),
    .Z(_06178_));
 CLKBUF_X3 _16031_ (.A(_05731_),
    .Z(_06179_));
 OAI221_X2 _16032_ (.A(_06175_),
    .B1(_06178_),
    .B2(_05938_),
    .C1(_06179_),
    .C2(_05943_),
    .ZN(_00533_));
 NAND2_X4 _16033_ (.A1(net104),
    .A2(\samples_real[5][10] ),
    .ZN(_06180_));
 OAI221_X2 _16034_ (.A(_06180_),
    .B1(_06178_),
    .B2(_05945_),
    .C1(_06179_),
    .C2(_05964_),
    .ZN(_00534_));
 NAND2_X4 _16035_ (.A1(\samples_real[5][11] ),
    .A2(_06174_),
    .ZN(_06181_));
 OAI221_X2 _16036_ (.A(_06181_),
    .B1(_06178_),
    .B2(_05966_),
    .C1(_06179_),
    .C2(_05972_),
    .ZN(_00535_));
 NAND2_X4 _16037_ (.A1(\samples_real[5][12] ),
    .A2(_06174_),
    .ZN(_06182_));
 OAI221_X2 _16038_ (.A(_06182_),
    .B1(_06178_),
    .B2(_05974_),
    .C1(_06179_),
    .C2(_05982_),
    .ZN(_00536_));
 NAND2_X4 _16039_ (.A1(net104),
    .A2(\samples_real[5][13] ),
    .ZN(_06183_));
 OAI221_X2 _16040_ (.A(_06183_),
    .B1(_06178_),
    .B2(_05984_),
    .C1(_06179_),
    .C2(_05988_),
    .ZN(_00537_));
 NAND2_X4 _16041_ (.A1(\samples_real[5][14] ),
    .A2(_06174_),
    .ZN(_06184_));
 OAI221_X2 _16042_ (.A(_06184_),
    .B1(_06178_),
    .B2(_05990_),
    .C1(_06179_),
    .C2(_05996_),
    .ZN(_00538_));
 NAND2_X2 _16043_ (.A1(_05998_),
    .A2(_06176_),
    .ZN(_06185_));
 NAND3_X1 _16044_ (.A1(_05672_),
    .A2(\samples_real[5][15] ),
    .A3(_06171_),
    .ZN(_06186_));
 NAND2_X1 _16045_ (.A1(_06185_),
    .A2(_06186_),
    .ZN(_06187_));
 MUX2_X1 _16046_ (.A(_06002_),
    .B(_06187_),
    .S(_06172_),
    .Z(_00539_));
 NAND2_X4 _16047_ (.A1(_06174_),
    .A2(\samples_real[5][1] ),
    .ZN(_06188_));
 OAI221_X2 _16048_ (.A(_06188_),
    .B1(_06178_),
    .B2(_06004_),
    .C1(_06179_),
    .C2(_06007_),
    .ZN(_00540_));
 NAND3_X4 _16049_ (.A1(_00855_),
    .A2(\samples_real[5][2] ),
    .A3(net487),
    .ZN(_06189_));
 OAI21_X2 _16050_ (.A(_06189_),
    .B1(_06012_),
    .B2(net518),
    .ZN(_06190_));
 MUX2_X1 _16051_ (.A(_06009_),
    .B(_06190_),
    .S(_06172_),
    .Z(_00541_));
 NAND2_X4 _16052_ (.A1(net104),
    .A2(\samples_real[5][3] ),
    .ZN(_06191_));
 OAI221_X2 _16053_ (.A(_06191_),
    .B1(_06178_),
    .B2(_06016_),
    .C1(_06179_),
    .C2(_06020_),
    .ZN(_00542_));
 NAND2_X4 _16054_ (.A1(net104),
    .A2(\samples_real[5][4] ),
    .ZN(_06192_));
 OAI221_X2 _16055_ (.A(_06192_),
    .B1(_06178_),
    .B2(_06022_),
    .C1(_06179_),
    .C2(_06027_),
    .ZN(_00543_));
 NAND2_X4 _16056_ (.A1(_06174_),
    .A2(\samples_real[5][5] ),
    .ZN(_06193_));
 OAI221_X2 _16057_ (.A(_06193_),
    .B1(_06178_),
    .B2(_06029_),
    .C1(_06179_),
    .C2(_06034_),
    .ZN(_00544_));
 NAND2_X2 _16058_ (.A1(_06173_),
    .A2(\samples_real[5][6] ),
    .ZN(_06194_));
 OAI221_X1 _16059_ (.A(_06194_),
    .B1(_06177_),
    .B2(_06036_),
    .C1(_05732_),
    .C2(_06041_),
    .ZN(_00545_));
 NAND2_X2 _16060_ (.A1(_06173_),
    .A2(\samples_real[5][7] ),
    .ZN(_06195_));
 OAI221_X1 _16061_ (.A(_06195_),
    .B1(_06177_),
    .B2(_06043_),
    .C1(_05732_),
    .C2(_06048_),
    .ZN(_00546_));
 NAND2_X2 _16062_ (.A1(_06173_),
    .A2(\samples_real[5][8] ),
    .ZN(_06196_));
 OAI221_X1 _16063_ (.A(_06196_),
    .B1(_06177_),
    .B2(_06050_),
    .C1(_05732_),
    .C2(_06055_),
    .ZN(_00547_));
 NAND2_X2 _16064_ (.A1(_06173_),
    .A2(\samples_real[5][9] ),
    .ZN(_06197_));
 OAI221_X1 _16065_ (.A(_06197_),
    .B1(_06177_),
    .B2(_06057_),
    .C1(_05732_),
    .C2(_06062_),
    .ZN(_00548_));
 MUX2_X2 _16066_ (.A(_05756_),
    .B(_05757_),
    .S(net453),
    .Z(_06198_));
 NAND2_X2 _16067_ (.A1(_05759_),
    .A2(_05859_),
    .ZN(_06199_));
 AND3_X4 _16068_ (.A1(_00842_),
    .A2(_06199_),
    .A3(_06198_),
    .ZN(_06200_));
 BUF_X8 _16069_ (.A(_06200_),
    .Z(_06201_));
 NAND2_X4 _16070_ (.A1(net107),
    .A2(\samples_real[6][0] ),
    .ZN(_06202_));
 INV_X4 _16071_ (.A(_06198_),
    .ZN(_06203_));
 NAND2_X4 _16072_ (.A1(_06203_),
    .A2(_06199_),
    .ZN(_06204_));
 BUF_X8 _16073_ (.A(_06204_),
    .Z(_06205_));
 CLKBUF_X3 _16074_ (.A(_05764_),
    .Z(_06206_));
 OAI221_X2 _16075_ (.A(_06202_),
    .B1(_06205_),
    .B2(_05938_),
    .C1(_06206_),
    .C2(_05943_),
    .ZN(_00549_));
 NAND2_X4 _16076_ (.A1(net107),
    .A2(\samples_real[6][10] ),
    .ZN(_06207_));
 OAI221_X2 _16077_ (.A(_06207_),
    .B1(_06205_),
    .B2(_05945_),
    .C1(_06206_),
    .C2(_05964_),
    .ZN(_00550_));
 NAND2_X4 _16078_ (.A1(_06201_),
    .A2(\samples_real[6][11] ),
    .ZN(_06208_));
 OAI221_X2 _16079_ (.A(_06208_),
    .B1(_06205_),
    .B2(_05966_),
    .C1(_06206_),
    .C2(_05972_),
    .ZN(_00551_));
 NAND2_X4 _16080_ (.A1(_06201_),
    .A2(\samples_real[6][12] ),
    .ZN(_06209_));
 OAI221_X2 _16081_ (.A(_06209_),
    .B1(_06205_),
    .B2(_05974_),
    .C1(_06206_),
    .C2(_05982_),
    .ZN(_00552_));
 NAND2_X4 _16082_ (.A1(net107),
    .A2(\samples_real[6][13] ),
    .ZN(_06210_));
 OAI221_X2 _16083_ (.A(_06210_),
    .B1(_06205_),
    .B2(_05984_),
    .C1(_06206_),
    .C2(_05988_),
    .ZN(_00553_));
 NAND2_X4 _16084_ (.A1(_06201_),
    .A2(\samples_real[6][14] ),
    .ZN(_06211_));
 OAI221_X2 _16085_ (.A(_06211_),
    .B1(_06205_),
    .B2(_05990_),
    .C1(_06206_),
    .C2(_05996_),
    .ZN(_00554_));
 NAND2_X2 _16086_ (.A1(_05998_),
    .A2(_06203_),
    .ZN(_06212_));
 NAND3_X1 _16087_ (.A1(_05596_),
    .A2(\samples_real[6][15] ),
    .A3(_06198_),
    .ZN(_06213_));
 NAND2_X1 _16088_ (.A1(_06212_),
    .A2(_06213_),
    .ZN(_06214_));
 MUX2_X1 _16089_ (.A(_06002_),
    .B(_06214_),
    .S(_06199_),
    .Z(_00555_));
 NAND2_X4 _16090_ (.A1(_06201_),
    .A2(\samples_real[6][1] ),
    .ZN(_06215_));
 OAI221_X2 _16091_ (.A(_06215_),
    .B1(_06205_),
    .B2(_06004_),
    .C1(_06206_),
    .C2(_06007_),
    .ZN(_00556_));
 NAND3_X1 _16092_ (.A1(_00855_),
    .A2(\samples_real[6][2] ),
    .A3(_06198_),
    .ZN(_06216_));
 OAI21_X2 _16093_ (.A(_06216_),
    .B1(_06012_),
    .B2(net514),
    .ZN(_06217_));
 MUX2_X1 _16094_ (.A(_06009_),
    .B(_06217_),
    .S(_06199_),
    .Z(_00557_));
 NAND2_X4 _16095_ (.A1(net107),
    .A2(\samples_real[6][3] ),
    .ZN(_06218_));
 OAI221_X2 _16096_ (.A(_06218_),
    .B1(_06205_),
    .B2(_06016_),
    .C1(_06206_),
    .C2(_06020_),
    .ZN(_00558_));
 NAND2_X4 _16097_ (.A1(net107),
    .A2(\samples_real[6][4] ),
    .ZN(_06219_));
 OAI221_X2 _16098_ (.A(_06219_),
    .B1(_06205_),
    .B2(_06022_),
    .C1(_06206_),
    .C2(_06027_),
    .ZN(_00559_));
 NAND2_X4 _16099_ (.A1(_06201_),
    .A2(\samples_real[6][5] ),
    .ZN(_06220_));
 OAI221_X1 _16100_ (.A(_06220_),
    .B1(_06205_),
    .B2(_06029_),
    .C1(_06206_),
    .C2(_06034_),
    .ZN(_00560_));
 NAND2_X4 _16101_ (.A1(_06200_),
    .A2(\samples_real[6][6] ),
    .ZN(_06221_));
 OAI221_X2 _16102_ (.A(_06221_),
    .B1(_06204_),
    .B2(_06036_),
    .C1(_05765_),
    .C2(_06041_),
    .ZN(_00561_));
 NAND2_X4 _16103_ (.A1(_06200_),
    .A2(\samples_real[6][7] ),
    .ZN(_06222_));
 OAI221_X2 _16104_ (.A(_06222_),
    .B1(_06204_),
    .B2(_06043_),
    .C1(_05765_),
    .C2(_06048_),
    .ZN(_00562_));
 NAND2_X2 _16105_ (.A1(_06200_),
    .A2(\samples_real[6][8] ),
    .ZN(_06223_));
 OAI221_X1 _16106_ (.A(_06223_),
    .B1(_06204_),
    .B2(_06050_),
    .C1(_05765_),
    .C2(_06055_),
    .ZN(_00563_));
 NAND2_X2 _16107_ (.A1(_06200_),
    .A2(\samples_real[6][9] ),
    .ZN(_06224_));
 OAI221_X1 _16108_ (.A(_06224_),
    .B1(_06204_),
    .B2(_06057_),
    .C1(_05765_),
    .C2(_06062_),
    .ZN(_00564_));
 MUX2_X2 _16109_ (.A(_05787_),
    .B(_05788_),
    .S(net453),
    .Z(_06225_));
 NAND4_X4 _16110_ (.A1(_04794_),
    .A2(_04791_),
    .A3(_04790_),
    .A4(_05859_),
    .ZN(_06226_));
 AND3_X4 _16111_ (.A1(_00842_),
    .A2(_06226_),
    .A3(_06225_),
    .ZN(_06227_));
 BUF_X16 _16112_ (.A(_06227_),
    .Z(_06228_));
 NAND2_X4 _16113_ (.A1(_06228_),
    .A2(\samples_real[7][0] ),
    .ZN(_06229_));
 INV_X4 _16114_ (.A(_06225_),
    .ZN(_06230_));
 NAND2_X4 _16115_ (.A1(_06230_),
    .A2(_06226_),
    .ZN(_06231_));
 BUF_X8 _16116_ (.A(_06231_),
    .Z(_06232_));
 CLKBUF_X3 _16117_ (.A(_05794_),
    .Z(_06233_));
 OAI221_X2 _16118_ (.A(_06229_),
    .B1(_06232_),
    .B2(_05938_),
    .C1(_06233_),
    .C2(_05943_),
    .ZN(_00565_));
 NAND2_X4 _16119_ (.A1(_06228_),
    .A2(\samples_real[7][10] ),
    .ZN(_06234_));
 OAI221_X2 _16120_ (.A(_06234_),
    .B1(_06232_),
    .B2(_05945_),
    .C1(_06233_),
    .C2(_05964_),
    .ZN(_00566_));
 NAND2_X4 _16121_ (.A1(_06228_),
    .A2(\samples_real[7][11] ),
    .ZN(_06235_));
 OAI221_X2 _16122_ (.A(_06235_),
    .B1(_06232_),
    .B2(_05966_),
    .C1(_06233_),
    .C2(_05972_),
    .ZN(_00567_));
 NAND2_X4 _16123_ (.A1(net516),
    .A2(\samples_real[7][12] ),
    .ZN(_06236_));
 OAI221_X2 _16124_ (.A(_06236_),
    .B1(_06232_),
    .B2(_05974_),
    .C1(_06233_),
    .C2(_05982_),
    .ZN(_00568_));
 NAND2_X4 _16125_ (.A1(_06228_),
    .A2(\samples_real[7][13] ),
    .ZN(_06237_));
 OAI221_X2 _16126_ (.A(_06237_),
    .B1(_06232_),
    .B2(_05984_),
    .C1(_06233_),
    .C2(_05988_),
    .ZN(_00569_));
 NAND2_X4 _16127_ (.A1(net516),
    .A2(\samples_real[7][14] ),
    .ZN(_06238_));
 OAI221_X2 _16128_ (.A(_06238_),
    .B1(_06232_),
    .B2(_05990_),
    .C1(_06233_),
    .C2(_05996_),
    .ZN(_00570_));
 NAND2_X2 _16129_ (.A1(_05998_),
    .A2(_06230_),
    .ZN(_06239_));
 NAND3_X1 _16130_ (.A1(_05596_),
    .A2(\samples_real[7][15] ),
    .A3(_06225_),
    .ZN(_06240_));
 NAND2_X1 _16131_ (.A1(_06239_),
    .A2(_06240_),
    .ZN(_06241_));
 MUX2_X1 _16132_ (.A(_06002_),
    .B(_06241_),
    .S(_06226_),
    .Z(_00571_));
 NAND2_X4 _16133_ (.A1(net516),
    .A2(\samples_real[7][1] ),
    .ZN(_06242_));
 OAI221_X2 _16134_ (.A(_06242_),
    .B1(_06232_),
    .B2(_06004_),
    .C1(_06233_),
    .C2(_06007_),
    .ZN(_00572_));
 NAND3_X2 _16135_ (.A1(_00855_),
    .A2(_06225_),
    .A3(\samples_real[7][2] ),
    .ZN(_06243_));
 OAI21_X2 _16136_ (.A(_06243_),
    .B1(_06012_),
    .B2(net515),
    .ZN(_06244_));
 MUX2_X1 _16137_ (.A(_06009_),
    .B(_06244_),
    .S(_06226_),
    .Z(_00573_));
 NAND2_X4 _16138_ (.A1(\samples_real[7][3] ),
    .A2(net516),
    .ZN(_06245_));
 OAI221_X1 _16139_ (.A(_06245_),
    .B1(_06232_),
    .B2(_06016_),
    .C1(_06233_),
    .C2(_06020_),
    .ZN(_00574_));
 NAND2_X4 _16140_ (.A1(net516),
    .A2(\samples_real[7][4] ),
    .ZN(_06246_));
 OAI221_X2 _16141_ (.A(_06246_),
    .B1(_06232_),
    .B2(_06022_),
    .C1(_06233_),
    .C2(_06027_),
    .ZN(_00575_));
 NAND2_X4 _16142_ (.A1(\samples_real[7][5] ),
    .A2(_06228_),
    .ZN(_06247_));
 OAI221_X2 _16143_ (.A(_06247_),
    .B1(_06232_),
    .B2(_06029_),
    .C1(_06233_),
    .C2(_06034_),
    .ZN(_00576_));
 NAND2_X4 _16144_ (.A1(_06227_),
    .A2(\samples_real[7][6] ),
    .ZN(_06248_));
 OAI221_X2 _16145_ (.A(_06248_),
    .B1(_06231_),
    .B2(_06036_),
    .C1(_05795_),
    .C2(_06041_),
    .ZN(_00577_));
 NAND2_X2 _16146_ (.A1(_06227_),
    .A2(\samples_real[7][7] ),
    .ZN(_06249_));
 OAI221_X1 _16147_ (.A(_06249_),
    .B1(_06231_),
    .B2(_06043_),
    .C1(_05795_),
    .C2(_06048_),
    .ZN(_00578_));
 NAND2_X2 _16148_ (.A1(_06227_),
    .A2(\samples_real[7][8] ),
    .ZN(_06250_));
 OAI221_X1 _16149_ (.A(_06250_),
    .B1(_06231_),
    .B2(_06050_),
    .C1(_05795_),
    .C2(_06055_),
    .ZN(_00579_));
 NAND2_X2 _16150_ (.A1(_06227_),
    .A2(\samples_real[7][9] ),
    .ZN(_06251_));
 OAI221_X1 _16151_ (.A(_06251_),
    .B1(_06231_),
    .B2(_06057_),
    .C1(_05795_),
    .C2(_06062_),
    .ZN(_00580_));
 XNOR2_X1 _16152_ (.A(_04839_),
    .B(_04925_),
    .ZN(_06252_));
 XNOR2_X1 _16153_ (.A(_04990_),
    .B(_06252_),
    .ZN(_06253_));
 NOR2_X1 _16154_ (.A1(_04823_),
    .A2(_06253_),
    .ZN(_06254_));
 XNOR2_X1 _16155_ (.A(_04894_),
    .B(_04944_),
    .ZN(_06255_));
 XNOR2_X1 _16156_ (.A(_04882_),
    .B(_06255_),
    .ZN(_06256_));
 NOR2_X1 _16157_ (.A1(_04808_),
    .A2(_06256_),
    .ZN(_06257_));
 XNOR2_X1 _16158_ (.A(_06254_),
    .B(_06257_),
    .ZN(_06258_));
 MUX2_X1 _16159_ (.A(\samples_imag[0][15] ),
    .B(\samples_imag[2][15] ),
    .S(_04875_),
    .Z(_06259_));
 MUX2_X1 _16160_ (.A(\samples_imag[1][15] ),
    .B(\samples_imag[3][15] ),
    .S(_04875_),
    .Z(_06260_));
 MUX2_X1 _16161_ (.A(_06259_),
    .B(_06260_),
    .S(_04867_),
    .Z(_06261_));
 MUX2_X1 _16162_ (.A(\samples_imag[4][15] ),
    .B(\samples_imag[6][15] ),
    .S(_04875_),
    .Z(_06262_));
 MUX2_X1 _16163_ (.A(\samples_imag[5][15] ),
    .B(\samples_imag[7][15] ),
    .S(_04875_),
    .Z(_06263_));
 MUX2_X1 _16164_ (.A(_06262_),
    .B(_06263_),
    .S(_04867_),
    .Z(_06264_));
 MUX2_X1 _16165_ (.A(_06261_),
    .B(_06264_),
    .S(_04893_),
    .Z(_06265_));
 NAND2_X1 _16166_ (.A1(_00022_),
    .A2(_06265_),
    .ZN(_06266_));
 XOR2_X1 _16167_ (.A(_07702_),
    .B(_06266_),
    .Z(_06267_));
 NAND2_X1 _16168_ (.A1(_04981_),
    .A2(_05117_),
    .ZN(_06268_));
 OR2_X1 _16169_ (.A1(_04865_),
    .A2(_05001_),
    .ZN(_06269_));
 XNOR2_X1 _16170_ (.A(_06268_),
    .B(_06269_),
    .ZN(_06270_));
 XNOR2_X1 _16171_ (.A(_06267_),
    .B(_06270_),
    .ZN(_06271_));
 XNOR2_X1 _16172_ (.A(_07401_),
    .B(_07559_),
    .ZN(_06272_));
 XNOR2_X2 _16173_ (.A(_07377_),
    .B(_07410_),
    .ZN(_06273_));
 XNOR2_X2 _16174_ (.A(_06272_),
    .B(_06273_),
    .ZN(_06274_));
 XNOR2_X2 _16175_ (.A(_06271_),
    .B(_06274_),
    .ZN(_06275_));
 XNOR2_X2 _16176_ (.A(_06258_),
    .B(_06275_),
    .ZN(_06276_));
 NAND4_X1 _16177_ (.A1(_09471_),
    .A2(_09511_),
    .A3(_09540_),
    .A4(_09558_),
    .ZN(_06277_));
 NAND4_X1 _16178_ (.A1(_09528_),
    .A2(_09565_),
    .A3(_09485_),
    .A4(_09499_),
    .ZN(_06278_));
 NOR2_X1 _16179_ (.A1(_06277_),
    .A2(_06278_),
    .ZN(_06279_));
 INV_X1 _16180_ (.A(_09571_),
    .ZN(_06280_));
 INV_X1 _16181_ (.A(_07911_),
    .ZN(_06281_));
 NAND4_X1 _16182_ (.A1(_06281_),
    .A2(_09572_),
    .A3(_09574_),
    .A4(_09576_),
    .ZN(_06282_));
 AOI21_X1 _16183_ (.A(_09582_),
    .B1(_07653_),
    .B2(_09583_),
    .ZN(_06283_));
 OAI21_X2 _16184_ (.A(_06280_),
    .B1(_06282_),
    .B2(_06283_),
    .ZN(_06284_));
 INV_X1 _16185_ (.A(_09484_),
    .ZN(_06285_));
 INV_X1 _16186_ (.A(_09510_),
    .ZN(_06286_));
 INV_X1 _16187_ (.A(_09511_),
    .ZN(_06287_));
 INV_X1 _16188_ (.A(_09539_),
    .ZN(_06288_));
 AOI21_X1 _16189_ (.A(_09557_),
    .B1(_09558_),
    .B2(_09564_),
    .ZN(_06289_));
 INV_X1 _16190_ (.A(_09540_),
    .ZN(_06290_));
 OAI21_X1 _16191_ (.A(_06288_),
    .B1(_06289_),
    .B2(_06290_),
    .ZN(_06291_));
 AOI21_X1 _16192_ (.A(_09527_),
    .B1(_06291_),
    .B2(_09528_),
    .ZN(_06292_));
 OAI21_X1 _16193_ (.A(_06286_),
    .B1(_06287_),
    .B2(_06292_),
    .ZN(_06293_));
 AOI21_X1 _16194_ (.A(_09498_),
    .B1(_06293_),
    .B2(_09499_),
    .ZN(_06294_));
 INV_X1 _16195_ (.A(_09485_),
    .ZN(_06295_));
 OAI21_X1 _16196_ (.A(_06285_),
    .B1(_06294_),
    .B2(_06295_),
    .ZN(_06296_));
 AOI221_X2 _16197_ (.A(_09470_),
    .B1(_06279_),
    .B2(_06284_),
    .C1(_06296_),
    .C2(_09471_),
    .ZN(_06297_));
 NOR2_X1 _16198_ (.A1(_04992_),
    .A2(_05010_),
    .ZN(_06298_));
 INV_X1 _16199_ (.A(_00034_),
    .ZN(_06299_));
 NAND2_X1 _16200_ (.A1(_06299_),
    .A2(_04822_),
    .ZN(_06300_));
 XOR2_X2 _16201_ (.A(_06298_),
    .B(_06300_),
    .Z(_06301_));
 NAND2_X1 _16202_ (.A1(_00046_),
    .A2(_05055_),
    .ZN(_06302_));
 XOR2_X1 _16203_ (.A(_09411_),
    .B(_07479_),
    .Z(_06303_));
 XNOR2_X1 _16204_ (.A(_09409_),
    .B(_09399_),
    .ZN(_06304_));
 XNOR2_X1 _16205_ (.A(_06303_),
    .B(_06304_),
    .ZN(_06305_));
 XNOR2_X1 _16206_ (.A(_07429_),
    .B(_07488_),
    .ZN(_06306_));
 XNOR2_X1 _16207_ (.A(_07402_),
    .B(_09396_),
    .ZN(_06307_));
 XNOR2_X1 _16208_ (.A(_06306_),
    .B(_06307_),
    .ZN(_06308_));
 XNOR2_X1 _16209_ (.A(_06305_),
    .B(_06308_),
    .ZN(_06309_));
 XOR2_X1 _16210_ (.A(_07395_),
    .B(_07375_),
    .Z(_06310_));
 XNOR2_X1 _16211_ (.A(_07469_),
    .B(_07536_),
    .ZN(_06311_));
 XNOR2_X1 _16212_ (.A(_06310_),
    .B(_06311_),
    .ZN(_06312_));
 XNOR2_X1 _16213_ (.A(_07420_),
    .B(_07433_),
    .ZN(_06313_));
 XNOR2_X1 _16214_ (.A(_07384_),
    .B(_07407_),
    .ZN(_06314_));
 XNOR2_X1 _16215_ (.A(_06313_),
    .B(_06314_),
    .ZN(_06315_));
 XNOR2_X1 _16216_ (.A(_06312_),
    .B(_06315_),
    .ZN(_06316_));
 XNOR2_X1 _16217_ (.A(_06309_),
    .B(_06316_),
    .ZN(_06317_));
 XOR2_X1 _16218_ (.A(_07437_),
    .B(_09392_),
    .Z(_06318_));
 XNOR2_X1 _16219_ (.A(_07399_),
    .B(_07389_),
    .ZN(_06319_));
 XNOR2_X1 _16220_ (.A(_06318_),
    .B(_06319_),
    .ZN(_06320_));
 XNOR2_X1 _16221_ (.A(_07460_),
    .B(_09408_),
    .ZN(_06321_));
 XNOR2_X1 _16222_ (.A(_09386_),
    .B(_09389_),
    .ZN(_06322_));
 XNOR2_X1 _16223_ (.A(_06321_),
    .B(_06322_),
    .ZN(_06323_));
 XNOR2_X1 _16224_ (.A(_06320_),
    .B(_06323_),
    .ZN(_06324_));
 XNOR2_X2 _16225_ (.A(_07629_),
    .B(_07586_),
    .ZN(_06325_));
 XNOR2_X1 _16226_ (.A(_07474_),
    .B(_07483_),
    .ZN(_06326_));
 XNOR2_X1 _16227_ (.A(_06326_),
    .B(_06325_),
    .ZN(_06327_));
 XNOR2_X1 _16228_ (.A(_06327_),
    .B(_06324_),
    .ZN(_06328_));
 XNOR2_X1 _16229_ (.A(_06328_),
    .B(_06317_),
    .ZN(_06329_));
 XOR2_X2 _16230_ (.A(_00045_),
    .B(_00046_),
    .Z(_06330_));
 XNOR2_X1 _16231_ (.A(_07527_),
    .B(_09446_),
    .ZN(_06331_));
 XNOR2_X1 _16232_ (.A(_07539_),
    .B(_09417_),
    .ZN(_06332_));
 XNOR2_X1 _16233_ (.A(_06331_),
    .B(_06332_),
    .ZN(_06333_));
 XNOR2_X1 _16234_ (.A(_06330_),
    .B(_06333_),
    .ZN(_06334_));
 XNOR2_X1 _16235_ (.A(_06334_),
    .B(_06329_),
    .ZN(_06335_));
 XNOR2_X1 _16236_ (.A(_06335_),
    .B(_06302_),
    .ZN(_06336_));
 XNOR2_X1 _16237_ (.A(_06336_),
    .B(_06301_),
    .ZN(_06337_));
 XNOR2_X1 _16238_ (.A(_06337_),
    .B(_06297_),
    .ZN(_06338_));
 XNOR2_X2 _16239_ (.A(_06338_),
    .B(_06276_),
    .ZN(_06339_));
 MUX2_X1 _16240_ (.A(\temp_imag[0] ),
    .B(_06339_),
    .S(_04778_),
    .Z(_00584_));
 XNOR2_X1 _16241_ (.A(_07984_),
    .B(_07986_),
    .ZN(_06340_));
 XNOR2_X1 _16242_ (.A(_08332_),
    .B(_08256_),
    .ZN(_06341_));
 XNOR2_X1 _16243_ (.A(_06340_),
    .B(_06341_),
    .ZN(_06342_));
 XNOR2_X1 _16244_ (.A(_08135_),
    .B(_07985_),
    .ZN(_06343_));
 XNOR2_X1 _16245_ (.A(_08105_),
    .B(_08004_),
    .ZN(_06344_));
 XNOR2_X1 _16246_ (.A(_06343_),
    .B(_06344_),
    .ZN(_06345_));
 XNOR2_X1 _16247_ (.A(_06342_),
    .B(_06345_),
    .ZN(_06346_));
 MUX2_X1 _16248_ (.A(\samples_real[0][15] ),
    .B(\samples_real[2][15] ),
    .S(net52),
    .Z(_06347_));
 MUX2_X1 _16249_ (.A(\samples_real[1][15] ),
    .B(\samples_real[3][15] ),
    .S(net52),
    .Z(_06348_));
 MUX2_X1 _16250_ (.A(_06347_),
    .B(_06348_),
    .S(_04851_),
    .Z(_06349_));
 MUX2_X1 _16251_ (.A(\samples_real[4][15] ),
    .B(\samples_real[6][15] ),
    .S(net52),
    .Z(_06350_));
 MUX2_X1 _16252_ (.A(\samples_real[5][15] ),
    .B(\samples_real[7][15] ),
    .S(net52),
    .Z(_06351_));
 MUX2_X1 _16253_ (.A(_06350_),
    .B(_06351_),
    .S(_04830_),
    .Z(_06352_));
 MUX2_X1 _16254_ (.A(_06349_),
    .B(_06352_),
    .S(_04847_),
    .Z(_06353_));
 NAND2_X1 _16255_ (.A1(_00022_),
    .A2(_06353_),
    .ZN(_06354_));
 XOR2_X1 _16256_ (.A(_08019_),
    .B(_06354_),
    .Z(_06355_));
 NAND2_X1 _16257_ (.A1(_05125_),
    .A2(_05117_),
    .ZN(_06356_));
 INV_X1 _16258_ (.A(_00021_),
    .ZN(_06357_));
 OR2_X1 _16259_ (.A1(_06357_),
    .A2(_05010_),
    .ZN(_06358_));
 XNOR2_X1 _16260_ (.A(_06356_),
    .B(_06358_),
    .ZN(_06359_));
 XNOR2_X1 _16261_ (.A(_06355_),
    .B(_06359_),
    .ZN(_06360_));
 NAND2_X1 _16262_ (.A1(_00046_),
    .A2(_04822_),
    .ZN(_06361_));
 NAND2_X1 _16263_ (.A1(_06299_),
    .A2(_05055_),
    .ZN(_06362_));
 XOR2_X1 _16264_ (.A(_06361_),
    .B(_06362_),
    .Z(_06363_));
 NAND2_X1 _16265_ (.A1(_00024_),
    .A2(_05121_),
    .ZN(_06364_));
 XNOR2_X1 _16266_ (.A(_07994_),
    .B(_06364_),
    .ZN(_06365_));
 XNOR2_X1 _16267_ (.A(_06363_),
    .B(_06365_),
    .ZN(_06366_));
 XNOR2_X1 _16268_ (.A(_06360_),
    .B(_06366_),
    .ZN(_06367_));
 XNOR2_X1 _16269_ (.A(_06346_),
    .B(_06367_),
    .ZN(_06368_));
 XNOR2_X2 _16270_ (.A(_08214_),
    .B(_09597_),
    .ZN(_06369_));
 XNOR2_X1 _16271_ (.A(_07974_),
    .B(_08152_),
    .ZN(_06370_));
 XNOR2_X2 _16272_ (.A(_06369_),
    .B(_06370_),
    .ZN(_06371_));
 XNOR2_X1 _16273_ (.A(_08026_),
    .B(_08088_),
    .ZN(_06372_));
 XNOR2_X1 _16274_ (.A(_07992_),
    .B(_08015_),
    .ZN(_06373_));
 XNOR2_X1 _16275_ (.A(_06372_),
    .B(_06373_),
    .ZN(_06374_));
 XNOR2_X2 _16276_ (.A(_06371_),
    .B(_06374_),
    .ZN(_06375_));
 XOR2_X1 _16277_ (.A(_07942_),
    .B(_07960_),
    .Z(_06376_));
 XNOR2_X1 _16278_ (.A(_08092_),
    .B(_09615_),
    .ZN(_06377_));
 XNOR2_X1 _16279_ (.A(_06376_),
    .B(_06377_),
    .ZN(_06378_));
 XNOR2_X1 _16280_ (.A(_08063_),
    .B(_07934_),
    .ZN(_06379_));
 XNOR2_X1 _16281_ (.A(_06330_),
    .B(_06379_),
    .ZN(_06380_));
 XNOR2_X1 _16282_ (.A(_06378_),
    .B(_06380_),
    .ZN(_06381_));
 XNOR2_X2 _16283_ (.A(_06375_),
    .B(_06381_),
    .ZN(_06382_));
 XNOR2_X2 _16284_ (.A(_06382_),
    .B(_07953_),
    .ZN(_06383_));
 XNOR2_X1 _16285_ (.A(_04839_),
    .B(_05046_),
    .ZN(_06384_));
 NOR2_X1 _16286_ (.A1(_04895_),
    .A2(_06384_),
    .ZN(_06385_));
 XNOR2_X1 _16287_ (.A(_06385_),
    .B(_06383_),
    .ZN(_06386_));
 XNOR2_X1 _16288_ (.A(_08002_),
    .B(_07997_),
    .ZN(_06387_));
 XNOR2_X1 _16289_ (.A(_07946_),
    .B(_09594_),
    .ZN(_06388_));
 XNOR2_X1 _16290_ (.A(_06387_),
    .B(_06388_),
    .ZN(_06389_));
 XNOR2_X1 _16291_ (.A(_09591_),
    .B(_08029_),
    .ZN(_06390_));
 XNOR2_X1 _16292_ (.A(_07937_),
    .B(_08069_),
    .ZN(_06391_));
 XNOR2_X1 _16293_ (.A(_06390_),
    .B(_06391_),
    .ZN(_06392_));
 XNOR2_X1 _16294_ (.A(_06389_),
    .B(_06392_),
    .ZN(_06393_));
 XOR2_X2 _16295_ (.A(_07979_),
    .B(_07982_),
    .Z(_06394_));
 XNOR2_X1 _16296_ (.A(_09584_),
    .B(_07917_),
    .ZN(_06395_));
 XNOR2_X1 _16297_ (.A(_06394_),
    .B(_06395_),
    .ZN(_06396_));
 XNOR2_X1 _16298_ (.A(_07918_),
    .B(_07926_),
    .ZN(_06397_));
 XNOR2_X1 _16299_ (.A(_07922_),
    .B(_09587_),
    .ZN(_06398_));
 XNOR2_X1 _16300_ (.A(_06397_),
    .B(_06398_),
    .ZN(_06399_));
 XNOR2_X1 _16301_ (.A(_06396_),
    .B(_06399_),
    .ZN(_06400_));
 XNOR2_X1 _16302_ (.A(_06393_),
    .B(_06400_),
    .ZN(_06401_));
 XNOR2_X1 _16303_ (.A(_08126_),
    .B(_08127_),
    .ZN(_06402_));
 XNOR2_X1 _16304_ (.A(_06401_),
    .B(_06402_),
    .ZN(_06403_));
 XNOR2_X1 _16305_ (.A(_06386_),
    .B(_06403_),
    .ZN(_06404_));
 XNOR2_X1 _16306_ (.A(_06404_),
    .B(_06368_),
    .ZN(_06405_));
 INV_X1 _16307_ (.A(_09647_),
    .ZN(_06406_));
 INV_X1 _16308_ (.A(_09662_),
    .ZN(_06407_));
 INV_X1 _16309_ (.A(_09689_),
    .ZN(_06408_));
 INV_X1 _16310_ (.A(_09702_),
    .ZN(_06409_));
 INV_X1 _16311_ (.A(_09718_),
    .ZN(_06410_));
 NAND4_X1 _16312_ (.A1(_08547_),
    .A2(_09747_),
    .A3(_09745_),
    .A4(_09750_),
    .ZN(_06411_));
 NOR3_X1 _16313_ (.A1(_06411_),
    .A2(_08424_),
    .A3(_08552_),
    .ZN(_06412_));
 OAI21_X1 _16314_ (.A(_09736_),
    .B1(_09744_),
    .B2(_06412_),
    .ZN(_06413_));
 INV_X1 _16315_ (.A(_06413_),
    .ZN(_06414_));
 OAI21_X1 _16316_ (.A(_09729_),
    .B1(_09735_),
    .B2(_06414_),
    .ZN(_06415_));
 INV_X1 _16317_ (.A(_09728_),
    .ZN(_06416_));
 AOI21_X1 _16318_ (.A(_06410_),
    .B1(_06415_),
    .B2(_06416_),
    .ZN(_06417_));
 OAI21_X1 _16319_ (.A(_09703_),
    .B1(_09717_),
    .B2(_06417_),
    .ZN(_06418_));
 AOI21_X1 _16320_ (.A(_06408_),
    .B1(_06409_),
    .B2(_06418_),
    .ZN(_06419_));
 OAI21_X1 _16321_ (.A(_09673_),
    .B1(_09688_),
    .B2(_06419_),
    .ZN(_06420_));
 INV_X1 _16322_ (.A(_09672_),
    .ZN(_06421_));
 AOI21_X1 _16323_ (.A(_06407_),
    .B1(_06420_),
    .B2(_06421_),
    .ZN(_06422_));
 OAI21_X1 _16324_ (.A(_09648_),
    .B1(_09661_),
    .B2(_06422_),
    .ZN(_06423_));
 NAND2_X1 _16325_ (.A1(_06406_),
    .A2(_06423_),
    .ZN(_06424_));
 AOI21_X2 _16326_ (.A(_09631_),
    .B1(_06424_),
    .B2(_09632_),
    .ZN(_06425_));
 XNOR2_X2 _16327_ (.A(_06405_),
    .B(_06425_),
    .ZN(_06426_));
 MUX2_X1 _16328_ (.A(\temp_real[0] ),
    .B(_06426_),
    .S(_04778_),
    .Z(_00585_));
 NOR2_X1 _16329_ (.A1(_00006_),
    .A2(_00019_),
    .ZN(_00048_));
 INV_X1 _16330_ (.A(_00048_),
    .ZN(_00047_));
 INV_X1 _16331_ (.A(_00006_),
    .ZN(_06427_));
 NAND2_X1 _16332_ (.A1(_06427_),
    .A2(_00019_),
    .ZN(_00049_));
 NOR2_X1 _16333_ (.A1(_06427_),
    .A2(_00008_),
    .ZN(_00050_));
 NAND2_X1 _16334_ (.A1(net86),
    .A2(_00853_),
    .ZN(_06428_));
 MUX2_X1 _16335_ (.A(\sample_count[2] ),
    .B(\bit_rev_idx[0] ),
    .S(_06428_),
    .Z(_06429_));
 AND2_X1 _16336_ (.A1(_00856_),
    .A2(_06429_),
    .ZN(_00051_));
 MUX2_X1 _16337_ (.A(\sample_count[1] ),
    .B(\bit_rev_idx[1] ),
    .S(_06428_),
    .Z(_06430_));
 AND2_X1 _16338_ (.A1(_00856_),
    .A2(_06430_),
    .ZN(_00052_));
 MUX2_X1 _16339_ (.A(\sample_count[0] ),
    .B(\bit_rev_idx[2] ),
    .S(_06428_),
    .Z(_06431_));
 AND2_X1 _16340_ (.A1(_00856_),
    .A2(_06431_),
    .ZN(_00053_));
 OAI21_X1 _16341_ (.A(_04769_),
    .B1(_00858_),
    .B2(_00860_),
    .ZN(_06432_));
 MUX2_X1 _16342_ (.A(net88),
    .B(_00041_),
    .S(_06432_),
    .Z(_06433_));
 AND2_X1 _16343_ (.A1(_00856_),
    .A2(_06433_),
    .ZN(_00054_));
 NAND2_X1 _16344_ (.A1(_05264_),
    .A2(_04776_),
    .ZN(_06434_));
 NOR2_X1 _16345_ (.A1(_00031_),
    .A2(_00851_),
    .ZN(_06435_));
 NOR3_X2 _16346_ (.A1(_04771_),
    .A2(_09382_),
    .A3(_00020_),
    .ZN(_06436_));
 NAND2_X1 _16347_ (.A1(_04771_),
    .A2(_00853_),
    .ZN(_06437_));
 INV_X1 _16348_ (.A(_00031_),
    .ZN(_06438_));
 OAI21_X2 _16349_ (.A(_06437_),
    .B1(_06438_),
    .B2(_00853_),
    .ZN(_06439_));
 NOR3_X4 _16350_ (.A1(_06435_),
    .A2(_06436_),
    .A3(_06439_),
    .ZN(_06440_));
 MUX2_X1 _16351_ (.A(_05264_),
    .B(_06434_),
    .S(_06440_),
    .Z(_06441_));
 NOR2_X1 _16352_ (.A1(_00845_),
    .A2(_06441_),
    .ZN(_00055_));
 NAND3_X1 _16353_ (.A1(_09358_),
    .A2(_04776_),
    .A3(_06440_),
    .ZN(_06442_));
 INV_X1 _16354_ (.A(\butterfly_count[1] ),
    .ZN(_06443_));
 OAI21_X1 _16355_ (.A(_06442_),
    .B1(_06440_),
    .B2(_06443_),
    .ZN(_06444_));
 AND2_X1 _16356_ (.A1(_00856_),
    .A2(_06444_),
    .ZN(_00056_));
 NAND2_X1 _16357_ (.A1(_09359_),
    .A2(_04776_),
    .ZN(_06445_));
 MUX2_X1 _16358_ (.A(_01169_),
    .B(_06445_),
    .S(_06440_),
    .Z(_06446_));
 NOR2_X1 _16359_ (.A1(_00845_),
    .A2(_06446_),
    .ZN(_00057_));
 BUF_X4 _16360_ (.A(_00857_),
    .Z(_06447_));
 CLKBUF_X3 _16361_ (.A(_06447_),
    .Z(_06448_));
 NAND2_X1 _16362_ (.A1(_06448_),
    .A2(\samples_imag[0][0] ),
    .ZN(_06449_));
 NAND2_X1 _16363_ (.A1(_00859_),
    .A2(net89),
    .ZN(_06450_));
 AOI21_X1 _16364_ (.A(_00845_),
    .B1(_06449_),
    .B2(_06450_),
    .ZN(_00061_));
 NAND2_X1 _16365_ (.A1(_06448_),
    .A2(\samples_imag[6][4] ),
    .ZN(_06451_));
 NAND2_X1 _16366_ (.A1(_00859_),
    .A2(net90),
    .ZN(_06452_));
 AOI21_X1 _16367_ (.A(_00845_),
    .B1(_06451_),
    .B2(_06452_),
    .ZN(_00062_));
 NAND2_X1 _16368_ (.A1(_06448_),
    .A2(\samples_imag[6][5] ),
    .ZN(_06453_));
 NAND2_X1 _16369_ (.A1(_00859_),
    .A2(net91),
    .ZN(_06454_));
 AOI21_X1 _16370_ (.A(_00845_),
    .B1(_06453_),
    .B2(_06454_),
    .ZN(_00063_));
 CLKBUF_X3 _16371_ (.A(_00844_),
    .Z(_06455_));
 NAND2_X1 _16372_ (.A1(_06448_),
    .A2(\samples_imag[6][6] ),
    .ZN(_06456_));
 NAND2_X1 _16373_ (.A1(_00859_),
    .A2(net92),
    .ZN(_06457_));
 AOI21_X1 _16374_ (.A(_06455_),
    .B1(_06456_),
    .B2(_06457_),
    .ZN(_00064_));
 NAND2_X1 _16375_ (.A1(_06448_),
    .A2(\samples_imag[6][7] ),
    .ZN(_06458_));
 NAND2_X1 _16376_ (.A1(_00859_),
    .A2(net95),
    .ZN(_06459_));
 AOI21_X1 _16377_ (.A(_06455_),
    .B1(_06458_),
    .B2(_06459_),
    .ZN(_00065_));
 NAND2_X1 _16378_ (.A1(_06448_),
    .A2(\samples_imag[6][8] ),
    .ZN(_06460_));
 NAND2_X1 _16379_ (.A1(_00859_),
    .A2(net96),
    .ZN(_06461_));
 AOI21_X1 _16380_ (.A(_06455_),
    .B1(_06460_),
    .B2(_06461_),
    .ZN(_00066_));
 NAND2_X1 _16381_ (.A1(_06448_),
    .A2(\samples_imag[6][9] ),
    .ZN(_06462_));
 NAND2_X1 _16382_ (.A1(_00859_),
    .A2(net99),
    .ZN(_06463_));
 AOI21_X1 _16383_ (.A(_06455_),
    .B1(_06462_),
    .B2(_06463_),
    .ZN(_00067_));
 NAND2_X1 _16384_ (.A1(_06448_),
    .A2(\samples_imag[6][10] ),
    .ZN(_06464_));
 NAND2_X1 _16385_ (.A1(_00859_),
    .A2(net100),
    .ZN(_06465_));
 AOI21_X1 _16386_ (.A(_06455_),
    .B1(_06464_),
    .B2(_06465_),
    .ZN(_00068_));
 NAND2_X1 _16387_ (.A1(_06448_),
    .A2(\samples_imag[6][11] ),
    .ZN(_06466_));
 NAND2_X1 _16388_ (.A1(_00859_),
    .A2(net102),
    .ZN(_06467_));
 AOI21_X1 _16389_ (.A(_06455_),
    .B1(_06466_),
    .B2(_06467_),
    .ZN(_00069_));
 NAND2_X1 _16390_ (.A1(_06448_),
    .A2(\samples_imag[6][12] ),
    .ZN(_06468_));
 CLKBUF_X3 _16391_ (.A(_00858_),
    .Z(_06469_));
 CLKBUF_X3 _16392_ (.A(_06469_),
    .Z(_06470_));
 NAND2_X1 _16393_ (.A1(_06470_),
    .A2(net103),
    .ZN(_06471_));
 AOI21_X1 _16394_ (.A(_06455_),
    .B1(_06468_),
    .B2(_06471_),
    .ZN(_00070_));
 CLKBUF_X3 _16395_ (.A(_06447_),
    .Z(_06472_));
 NAND2_X1 _16396_ (.A1(_06472_),
    .A2(\samples_imag[6][13] ),
    .ZN(_06473_));
 NAND2_X1 _16397_ (.A1(_06470_),
    .A2(net105),
    .ZN(_06474_));
 AOI21_X1 _16398_ (.A(_06455_),
    .B1(_06473_),
    .B2(_06474_),
    .ZN(_00071_));
 NAND2_X1 _16399_ (.A1(_06472_),
    .A2(\samples_imag[0][10] ),
    .ZN(_06475_));
 NAND2_X1 _16400_ (.A1(_06470_),
    .A2(net106),
    .ZN(_06476_));
 AOI21_X1 _16401_ (.A(_06455_),
    .B1(_06475_),
    .B2(_06476_),
    .ZN(_00072_));
 NAND2_X1 _16402_ (.A1(_06472_),
    .A2(\samples_imag[6][14] ),
    .ZN(_06477_));
 NAND2_X1 _16403_ (.A1(_06470_),
    .A2(net108),
    .ZN(_06478_));
 AOI21_X1 _16404_ (.A(_06455_),
    .B1(_06477_),
    .B2(_06478_),
    .ZN(_00073_));
 CLKBUF_X3 _16405_ (.A(_00844_),
    .Z(_06479_));
 NAND2_X1 _16406_ (.A1(_06472_),
    .A2(\samples_imag[6][15] ),
    .ZN(_06480_));
 NAND2_X1 _16407_ (.A1(_06470_),
    .A2(net109),
    .ZN(_06481_));
 AOI21_X1 _16408_ (.A(_06479_),
    .B1(_06480_),
    .B2(_06481_),
    .ZN(_00074_));
 NAND2_X1 _16409_ (.A1(_06472_),
    .A2(\samples_imag[7][0] ),
    .ZN(_06482_));
 NAND2_X1 _16410_ (.A1(_06470_),
    .A2(net110),
    .ZN(_06483_));
 AOI21_X1 _16411_ (.A(_06479_),
    .B1(_06482_),
    .B2(_06483_),
    .ZN(_00075_));
 NAND2_X1 _16412_ (.A1(_06472_),
    .A2(\samples_imag[7][1] ),
    .ZN(_06484_));
 NAND2_X1 _16413_ (.A1(_06470_),
    .A2(net111),
    .ZN(_06485_));
 AOI21_X1 _16414_ (.A(_06479_),
    .B1(_06484_),
    .B2(_06485_),
    .ZN(_00076_));
 NAND2_X1 _16415_ (.A1(_06472_),
    .A2(\samples_imag[7][2] ),
    .ZN(_06486_));
 NAND2_X1 _16416_ (.A1(_06470_),
    .A2(net112),
    .ZN(_06487_));
 AOI21_X1 _16417_ (.A(_06479_),
    .B1(_06486_),
    .B2(_06487_),
    .ZN(_00077_));
 NAND2_X1 _16418_ (.A1(_06472_),
    .A2(\samples_imag[7][3] ),
    .ZN(_06488_));
 NAND2_X1 _16419_ (.A1(_06470_),
    .A2(net113),
    .ZN(_06489_));
 AOI21_X1 _16420_ (.A(_06479_),
    .B1(_06488_),
    .B2(_06489_),
    .ZN(_00078_));
 NAND2_X1 _16421_ (.A1(_06472_),
    .A2(\samples_imag[7][4] ),
    .ZN(_06490_));
 NAND2_X1 _16422_ (.A1(_06470_),
    .A2(net114),
    .ZN(_06491_));
 AOI21_X1 _16423_ (.A(_06479_),
    .B1(_06490_),
    .B2(_06491_),
    .ZN(_00079_));
 NAND2_X1 _16424_ (.A1(_06472_),
    .A2(\samples_imag[7][5] ),
    .ZN(_06492_));
 CLKBUF_X3 _16425_ (.A(_06469_),
    .Z(_06493_));
 NAND2_X1 _16426_ (.A1(_06493_),
    .A2(net115),
    .ZN(_06494_));
 AOI21_X1 _16427_ (.A(_06479_),
    .B1(_06492_),
    .B2(_06494_),
    .ZN(_00080_));
 CLKBUF_X3 _16428_ (.A(_06447_),
    .Z(_06495_));
 NAND2_X1 _16429_ (.A1(_06495_),
    .A2(\samples_imag[7][6] ),
    .ZN(_06496_));
 NAND2_X1 _16430_ (.A1(_06493_),
    .A2(net116),
    .ZN(_06497_));
 AOI21_X1 _16431_ (.A(_06479_),
    .B1(_06496_),
    .B2(_06497_),
    .ZN(_00081_));
 NAND2_X1 _16432_ (.A1(_06495_),
    .A2(\samples_imag[7][7] ),
    .ZN(_06498_));
 NAND2_X1 _16433_ (.A1(_06493_),
    .A2(net117),
    .ZN(_06499_));
 AOI21_X1 _16434_ (.A(_06479_),
    .B1(_06498_),
    .B2(_06499_),
    .ZN(_00082_));
 NAND2_X1 _16435_ (.A1(_06495_),
    .A2(\samples_imag[0][11] ),
    .ZN(_06500_));
 NAND2_X1 _16436_ (.A1(_06493_),
    .A2(net118),
    .ZN(_06501_));
 AOI21_X1 _16437_ (.A(_06479_),
    .B1(_06500_),
    .B2(_06501_),
    .ZN(_00083_));
 BUF_X4 _16438_ (.A(_00843_),
    .Z(_06502_));
 CLKBUF_X3 _16439_ (.A(_06502_),
    .Z(_06503_));
 NAND2_X1 _16440_ (.A1(_06495_),
    .A2(\samples_imag[7][8] ),
    .ZN(_06504_));
 NAND2_X1 _16441_ (.A1(_06493_),
    .A2(net119),
    .ZN(_06505_));
 AOI21_X1 _16442_ (.A(_06503_),
    .B1(_06504_),
    .B2(_06505_),
    .ZN(_00084_));
 NAND2_X1 _16443_ (.A1(_06495_),
    .A2(\samples_imag[7][9] ),
    .ZN(_06506_));
 NAND2_X1 _16444_ (.A1(_06493_),
    .A2(net120),
    .ZN(_06507_));
 AOI21_X1 _16445_ (.A(_06503_),
    .B1(_06506_),
    .B2(_06507_),
    .ZN(_00085_));
 NAND2_X1 _16446_ (.A1(_06495_),
    .A2(\samples_imag[7][10] ),
    .ZN(_06508_));
 NAND2_X1 _16447_ (.A1(_06493_),
    .A2(net121),
    .ZN(_06509_));
 AOI21_X1 _16448_ (.A(_06503_),
    .B1(_06508_),
    .B2(_06509_),
    .ZN(_00086_));
 NAND2_X1 _16449_ (.A1(_06495_),
    .A2(\samples_imag[7][11] ),
    .ZN(_06510_));
 NAND2_X1 _16450_ (.A1(_06493_),
    .A2(net122),
    .ZN(_06511_));
 AOI21_X1 _16451_ (.A(_06503_),
    .B1(_06510_),
    .B2(_06511_),
    .ZN(_00087_));
 NAND2_X1 _16452_ (.A1(_06495_),
    .A2(\samples_imag[7][12] ),
    .ZN(_06512_));
 NAND2_X1 _16453_ (.A1(_06493_),
    .A2(net123),
    .ZN(_06513_));
 AOI21_X1 _16454_ (.A(_06503_),
    .B1(_06512_),
    .B2(_06513_),
    .ZN(_00088_));
 NAND2_X1 _16455_ (.A1(_06495_),
    .A2(\samples_imag[7][13] ),
    .ZN(_06514_));
 NAND2_X1 _16456_ (.A1(_06493_),
    .A2(net124),
    .ZN(_06515_));
 AOI21_X1 _16457_ (.A(_06503_),
    .B1(_06514_),
    .B2(_06515_),
    .ZN(_00089_));
 NAND2_X1 _16458_ (.A1(_06495_),
    .A2(\samples_imag[7][14] ),
    .ZN(_06516_));
 CLKBUF_X3 _16459_ (.A(_00858_),
    .Z(_06517_));
 CLKBUF_X3 _16460_ (.A(_06517_),
    .Z(_06518_));
 NAND2_X1 _16461_ (.A1(_06518_),
    .A2(net126),
    .ZN(_06519_));
 AOI21_X1 _16462_ (.A(_06503_),
    .B1(_06516_),
    .B2(_06519_),
    .ZN(_00090_));
 BUF_X4 _16463_ (.A(_00857_),
    .Z(_06520_));
 CLKBUF_X3 _16464_ (.A(_06520_),
    .Z(_06521_));
 NAND2_X1 _16465_ (.A1(_06521_),
    .A2(\samples_imag[7][15] ),
    .ZN(_06522_));
 NAND2_X1 _16466_ (.A1(_06518_),
    .A2(net127),
    .ZN(_06523_));
 AOI21_X1 _16467_ (.A(_06503_),
    .B1(_06522_),
    .B2(_06523_),
    .ZN(_00091_));
 NAND2_X1 _16468_ (.A1(_06521_),
    .A2(\samples_imag[0][12] ),
    .ZN(_06524_));
 NAND2_X1 _16469_ (.A1(_06518_),
    .A2(net128),
    .ZN(_06525_));
 AOI21_X1 _16470_ (.A(_06503_),
    .B1(_06524_),
    .B2(_06525_),
    .ZN(_00092_));
 NAND2_X1 _16471_ (.A1(_06521_),
    .A2(\samples_imag[0][13] ),
    .ZN(_06526_));
 NAND2_X1 _16472_ (.A1(_06518_),
    .A2(net134),
    .ZN(_06527_));
 AOI21_X1 _16473_ (.A(_06503_),
    .B1(_06526_),
    .B2(_06527_),
    .ZN(_00093_));
 CLKBUF_X3 _16474_ (.A(_06502_),
    .Z(_06528_));
 NAND2_X1 _16475_ (.A1(_06521_),
    .A2(\samples_imag[0][14] ),
    .ZN(_06529_));
 NAND2_X1 _16476_ (.A1(_06518_),
    .A2(net135),
    .ZN(_06530_));
 AOI21_X1 _16477_ (.A(_06528_),
    .B1(_06529_),
    .B2(_06530_),
    .ZN(_00094_));
 NAND2_X1 _16478_ (.A1(_06521_),
    .A2(\samples_imag[0][15] ),
    .ZN(_06531_));
 NAND2_X1 _16479_ (.A1(_06518_),
    .A2(net136),
    .ZN(_06532_));
 AOI21_X1 _16480_ (.A(_06528_),
    .B1(_06531_),
    .B2(_06532_),
    .ZN(_00095_));
 NAND2_X1 _16481_ (.A1(_06521_),
    .A2(\samples_imag[1][0] ),
    .ZN(_06533_));
 NAND2_X1 _16482_ (.A1(_06518_),
    .A2(net141),
    .ZN(_06534_));
 AOI21_X1 _16483_ (.A(_06528_),
    .B1(_06533_),
    .B2(_06534_),
    .ZN(_00096_));
 NAND2_X1 _16484_ (.A1(_06521_),
    .A2(\samples_imag[1][1] ),
    .ZN(_06535_));
 NAND2_X1 _16485_ (.A1(_06518_),
    .A2(net142),
    .ZN(_06536_));
 AOI21_X1 _16486_ (.A(_06528_),
    .B1(_06535_),
    .B2(_06536_),
    .ZN(_00097_));
 NAND2_X1 _16487_ (.A1(_06521_),
    .A2(\samples_imag[1][2] ),
    .ZN(_06537_));
 NAND2_X1 _16488_ (.A1(_06518_),
    .A2(net145),
    .ZN(_06538_));
 AOI21_X1 _16489_ (.A(_06528_),
    .B1(_06537_),
    .B2(_06538_),
    .ZN(_00098_));
 NAND2_X1 _16490_ (.A1(_06521_),
    .A2(\samples_imag[1][3] ),
    .ZN(_06539_));
 NAND2_X1 _16491_ (.A1(_06518_),
    .A2(net146),
    .ZN(_06540_));
 AOI21_X1 _16492_ (.A(_06528_),
    .B1(_06539_),
    .B2(_06540_),
    .ZN(_00099_));
 NAND2_X1 _16493_ (.A1(_06521_),
    .A2(\samples_imag[0][1] ),
    .ZN(_06541_));
 CLKBUF_X3 _16494_ (.A(_06517_),
    .Z(_06542_));
 NAND2_X1 _16495_ (.A1(_06542_),
    .A2(net147),
    .ZN(_06543_));
 AOI21_X1 _16496_ (.A(_06528_),
    .B1(_06541_),
    .B2(_06543_),
    .ZN(_00100_));
 BUF_X2 _16497_ (.A(_06520_),
    .Z(_06544_));
 NAND2_X1 _16498_ (.A1(_06544_),
    .A2(\samples_imag[1][4] ),
    .ZN(_06545_));
 NAND2_X1 _16499_ (.A1(_06542_),
    .A2(net148),
    .ZN(_06546_));
 AOI21_X1 _16500_ (.A(_06528_),
    .B1(_06545_),
    .B2(_06546_),
    .ZN(_00101_));
 NAND2_X1 _16501_ (.A1(_06544_),
    .A2(\samples_imag[1][5] ),
    .ZN(_06547_));
 NAND2_X1 _16502_ (.A1(_06542_),
    .A2(net150),
    .ZN(_06548_));
 AOI21_X1 _16503_ (.A(_06528_),
    .B1(_06547_),
    .B2(_06548_),
    .ZN(_00102_));
 NAND2_X1 _16504_ (.A1(_06544_),
    .A2(\samples_imag[1][6] ),
    .ZN(_06549_));
 NAND2_X1 _16505_ (.A1(_06542_),
    .A2(net155),
    .ZN(_06550_));
 AOI21_X1 _16506_ (.A(_06528_),
    .B1(_06549_),
    .B2(_06550_),
    .ZN(_00103_));
 CLKBUF_X3 _16507_ (.A(_06502_),
    .Z(_06551_));
 NAND2_X1 _16508_ (.A1(_06544_),
    .A2(\samples_imag[1][7] ),
    .ZN(_06552_));
 NAND2_X1 _16509_ (.A1(_06542_),
    .A2(net157),
    .ZN(_06553_));
 AOI21_X1 _16510_ (.A(_06551_),
    .B1(_06552_),
    .B2(_06553_),
    .ZN(_00104_));
 NAND2_X1 _16511_ (.A1(_06544_),
    .A2(\samples_imag[1][8] ),
    .ZN(_06554_));
 NAND2_X1 _16512_ (.A1(_06542_),
    .A2(net159),
    .ZN(_06555_));
 AOI21_X1 _16513_ (.A(_06551_),
    .B1(_06554_),
    .B2(_06555_),
    .ZN(_00105_));
 NAND2_X1 _16514_ (.A1(_06544_),
    .A2(\samples_imag[1][9] ),
    .ZN(_06556_));
 NAND2_X1 _16515_ (.A1(_06542_),
    .A2(net160),
    .ZN(_06557_));
 AOI21_X1 _16516_ (.A(_06551_),
    .B1(_06556_),
    .B2(_06557_),
    .ZN(_00106_));
 NAND2_X1 _16517_ (.A1(_06544_),
    .A2(\samples_imag[1][10] ),
    .ZN(_06558_));
 NAND2_X1 _16518_ (.A1(_06542_),
    .A2(net161),
    .ZN(_06559_));
 AOI21_X1 _16519_ (.A(_06551_),
    .B1(_06558_),
    .B2(_06559_),
    .ZN(_00107_));
 NAND2_X1 _16520_ (.A1(_06544_),
    .A2(\samples_imag[1][11] ),
    .ZN(_06560_));
 NAND2_X1 _16521_ (.A1(_06542_),
    .A2(net162),
    .ZN(_06561_));
 AOI21_X1 _16522_ (.A(_06551_),
    .B1(_06560_),
    .B2(_06561_),
    .ZN(_00108_));
 NAND2_X1 _16523_ (.A1(_06544_),
    .A2(\samples_imag[1][12] ),
    .ZN(_06562_));
 NAND2_X1 _16524_ (.A1(_06542_),
    .A2(net163),
    .ZN(_06563_));
 AOI21_X1 _16525_ (.A(_06551_),
    .B1(_06562_),
    .B2(_06563_),
    .ZN(_00109_));
 NAND2_X1 _16526_ (.A1(_06544_),
    .A2(\samples_imag[1][13] ),
    .ZN(_06564_));
 CLKBUF_X3 _16527_ (.A(_06517_),
    .Z(_06565_));
 NAND2_X1 _16528_ (.A1(_06565_),
    .A2(net164),
    .ZN(_06566_));
 AOI21_X1 _16529_ (.A(_06551_),
    .B1(_06564_),
    .B2(_06566_),
    .ZN(_00110_));
 CLKBUF_X3 _16530_ (.A(_06520_),
    .Z(_06567_));
 NAND2_X1 _16531_ (.A1(_06567_),
    .A2(\samples_imag[0][2] ),
    .ZN(_06568_));
 NAND2_X1 _16532_ (.A1(_06565_),
    .A2(net165),
    .ZN(_06569_));
 AOI21_X1 _16533_ (.A(_06551_),
    .B1(_06568_),
    .B2(_06569_),
    .ZN(_00111_));
 NAND2_X1 _16534_ (.A1(_06567_),
    .A2(\samples_imag[1][14] ),
    .ZN(_06570_));
 NAND2_X1 _16535_ (.A1(_06565_),
    .A2(net166),
    .ZN(_06571_));
 AOI21_X1 _16536_ (.A(_06551_),
    .B1(_06570_),
    .B2(_06571_),
    .ZN(_00112_));
 NAND2_X1 _16537_ (.A1(_06567_),
    .A2(\samples_imag[1][15] ),
    .ZN(_06572_));
 NAND2_X1 _16538_ (.A1(_06565_),
    .A2(net167),
    .ZN(_06573_));
 AOI21_X1 _16539_ (.A(_06551_),
    .B1(_06572_),
    .B2(_06573_),
    .ZN(_00113_));
 CLKBUF_X3 _16540_ (.A(_06502_),
    .Z(_06574_));
 NAND2_X1 _16541_ (.A1(_06567_),
    .A2(\samples_imag[2][0] ),
    .ZN(_06575_));
 NAND2_X1 _16542_ (.A1(_06565_),
    .A2(net168),
    .ZN(_06576_));
 AOI21_X1 _16543_ (.A(_06574_),
    .B1(_06575_),
    .B2(_06576_),
    .ZN(_00114_));
 NAND2_X1 _16544_ (.A1(_06567_),
    .A2(\samples_imag[2][1] ),
    .ZN(_06577_));
 NAND2_X1 _16545_ (.A1(_06565_),
    .A2(net169),
    .ZN(_06578_));
 AOI21_X1 _16546_ (.A(_06574_),
    .B1(_06577_),
    .B2(_06578_),
    .ZN(_00115_));
 NAND2_X1 _16547_ (.A1(_06567_),
    .A2(\samples_imag[2][2] ),
    .ZN(_06579_));
 NAND2_X1 _16548_ (.A1(_06565_),
    .A2(net170),
    .ZN(_06580_));
 AOI21_X1 _16549_ (.A(_06574_),
    .B1(_06579_),
    .B2(_06580_),
    .ZN(_00116_));
 NAND2_X1 _16550_ (.A1(_06567_),
    .A2(\samples_imag[2][3] ),
    .ZN(_06581_));
 NAND2_X1 _16551_ (.A1(_06565_),
    .A2(net171),
    .ZN(_06582_));
 AOI21_X1 _16552_ (.A(_06574_),
    .B1(_06581_),
    .B2(_06582_),
    .ZN(_00117_));
 NAND2_X1 _16553_ (.A1(_06567_),
    .A2(\samples_imag[2][4] ),
    .ZN(_06583_));
 NAND2_X1 _16554_ (.A1(_06565_),
    .A2(net172),
    .ZN(_06584_));
 AOI21_X1 _16555_ (.A(_06574_),
    .B1(_06583_),
    .B2(_06584_),
    .ZN(_00118_));
 NAND2_X1 _16556_ (.A1(_06567_),
    .A2(\samples_imag[2][5] ),
    .ZN(_06585_));
 NAND2_X1 _16557_ (.A1(_06565_),
    .A2(net173),
    .ZN(_06586_));
 AOI21_X1 _16558_ (.A(_06574_),
    .B1(_06585_),
    .B2(_06586_),
    .ZN(_00119_));
 NAND2_X1 _16559_ (.A1(_06567_),
    .A2(\samples_imag[2][6] ),
    .ZN(_06587_));
 CLKBUF_X3 _16560_ (.A(_06517_),
    .Z(_06588_));
 NAND2_X1 _16561_ (.A1(_06588_),
    .A2(net174),
    .ZN(_06589_));
 AOI21_X1 _16562_ (.A(_06574_),
    .B1(_06587_),
    .B2(_06589_),
    .ZN(_00120_));
 CLKBUF_X3 _16563_ (.A(_06520_),
    .Z(_06590_));
 NAND2_X1 _16564_ (.A1(_06590_),
    .A2(\samples_imag[2][7] ),
    .ZN(_06591_));
 NAND2_X1 _16565_ (.A1(_06588_),
    .A2(net175),
    .ZN(_06592_));
 AOI21_X1 _16566_ (.A(_06574_),
    .B1(_06591_),
    .B2(_06592_),
    .ZN(_00121_));
 NAND2_X1 _16567_ (.A1(_06590_),
    .A2(\samples_imag[0][3] ),
    .ZN(_06593_));
 NAND2_X1 _16568_ (.A1(_06588_),
    .A2(net176),
    .ZN(_06594_));
 AOI21_X1 _16569_ (.A(_06574_),
    .B1(_06593_),
    .B2(_06594_),
    .ZN(_00122_));
 NAND2_X1 _16570_ (.A1(_06590_),
    .A2(\samples_imag[2][8] ),
    .ZN(_06595_));
 NAND2_X1 _16571_ (.A1(_06588_),
    .A2(net177),
    .ZN(_06596_));
 AOI21_X1 _16572_ (.A(_06574_),
    .B1(_06595_),
    .B2(_06596_),
    .ZN(_00123_));
 CLKBUF_X3 _16573_ (.A(_06502_),
    .Z(_06597_));
 NAND2_X1 _16574_ (.A1(_06590_),
    .A2(\samples_imag[2][9] ),
    .ZN(_06598_));
 NAND2_X1 _16575_ (.A1(_06588_),
    .A2(net178),
    .ZN(_06599_));
 AOI21_X1 _16576_ (.A(_06597_),
    .B1(_06598_),
    .B2(_06599_),
    .ZN(_00124_));
 NAND2_X1 _16577_ (.A1(_06590_),
    .A2(\samples_imag[2][10] ),
    .ZN(_06600_));
 NAND2_X1 _16578_ (.A1(_06588_),
    .A2(net179),
    .ZN(_06601_));
 AOI21_X1 _16579_ (.A(_06597_),
    .B1(_06600_),
    .B2(_06601_),
    .ZN(_00125_));
 NAND2_X1 _16580_ (.A1(_06590_),
    .A2(\samples_imag[2][11] ),
    .ZN(_06602_));
 NAND2_X1 _16581_ (.A1(_06588_),
    .A2(net180),
    .ZN(_06603_));
 AOI21_X1 _16582_ (.A(_06597_),
    .B1(_06602_),
    .B2(_06603_),
    .ZN(_00126_));
 NAND2_X1 _16583_ (.A1(_06590_),
    .A2(\samples_imag[2][12] ),
    .ZN(_06604_));
 NAND2_X1 _16584_ (.A1(_06588_),
    .A2(net181),
    .ZN(_06605_));
 AOI21_X1 _16585_ (.A(_06597_),
    .B1(_06604_),
    .B2(_06605_),
    .ZN(_00127_));
 NAND2_X1 _16586_ (.A1(_06590_),
    .A2(\samples_imag[2][13] ),
    .ZN(_06606_));
 NAND2_X1 _16587_ (.A1(_06588_),
    .A2(net182),
    .ZN(_06607_));
 AOI21_X1 _16588_ (.A(_06597_),
    .B1(_06606_),
    .B2(_06607_),
    .ZN(_00128_));
 NAND2_X1 _16589_ (.A1(_06590_),
    .A2(\samples_imag[2][14] ),
    .ZN(_06608_));
 NAND2_X1 _16590_ (.A1(_06588_),
    .A2(net183),
    .ZN(_06609_));
 AOI21_X1 _16591_ (.A(_06597_),
    .B1(_06608_),
    .B2(_06609_),
    .ZN(_00129_));
 NAND2_X1 _16592_ (.A1(_06590_),
    .A2(\samples_imag[2][15] ),
    .ZN(_06610_));
 CLKBUF_X3 _16593_ (.A(_06517_),
    .Z(_06611_));
 NAND2_X1 _16594_ (.A1(_06611_),
    .A2(net184),
    .ZN(_06612_));
 AOI21_X1 _16595_ (.A(_06597_),
    .B1(_06610_),
    .B2(_06612_),
    .ZN(_00130_));
 BUF_X2 _16596_ (.A(_06520_),
    .Z(_06613_));
 NAND2_X1 _16597_ (.A1(_06613_),
    .A2(\samples_imag[3][0] ),
    .ZN(_06614_));
 NAND2_X1 _16598_ (.A1(_06611_),
    .A2(net185),
    .ZN(_06615_));
 AOI21_X1 _16599_ (.A(_06597_),
    .B1(_06614_),
    .B2(_06615_),
    .ZN(_00131_));
 NAND2_X1 _16600_ (.A1(_06613_),
    .A2(\samples_imag[3][1] ),
    .ZN(_06616_));
 NAND2_X1 _16601_ (.A1(_06611_),
    .A2(net186),
    .ZN(_06617_));
 AOI21_X1 _16602_ (.A(_06597_),
    .B1(_06616_),
    .B2(_06617_),
    .ZN(_00132_));
 NAND2_X1 _16603_ (.A1(_06613_),
    .A2(\samples_imag[0][4] ),
    .ZN(_06618_));
 NAND2_X1 _16604_ (.A1(_06611_),
    .A2(net187),
    .ZN(_06619_));
 AOI21_X1 _16605_ (.A(_06597_),
    .B1(_06618_),
    .B2(_06619_),
    .ZN(_00133_));
 CLKBUF_X3 _16606_ (.A(_06502_),
    .Z(_06620_));
 NAND2_X1 _16607_ (.A1(_06613_),
    .A2(\samples_imag[3][2] ),
    .ZN(_06621_));
 NAND2_X1 _16608_ (.A1(_06611_),
    .A2(net188),
    .ZN(_06622_));
 AOI21_X1 _16609_ (.A(_06620_),
    .B1(_06621_),
    .B2(_06622_),
    .ZN(_00134_));
 NAND2_X1 _16610_ (.A1(_06613_),
    .A2(\samples_imag[3][3] ),
    .ZN(_06623_));
 NAND2_X1 _16611_ (.A1(_06611_),
    .A2(net189),
    .ZN(_06624_));
 AOI21_X1 _16612_ (.A(_06620_),
    .B1(_06623_),
    .B2(_06624_),
    .ZN(_00135_));
 NAND2_X1 _16613_ (.A1(_06613_),
    .A2(\samples_imag[3][4] ),
    .ZN(_06625_));
 NAND2_X1 _16614_ (.A1(_06611_),
    .A2(net190),
    .ZN(_06626_));
 AOI21_X1 _16615_ (.A(_06620_),
    .B1(_06625_),
    .B2(_06626_),
    .ZN(_00136_));
 NAND2_X1 _16616_ (.A1(_06613_),
    .A2(\samples_imag[3][5] ),
    .ZN(_06627_));
 NAND2_X1 _16617_ (.A1(_06611_),
    .A2(net191),
    .ZN(_06628_));
 AOI21_X1 _16618_ (.A(_06620_),
    .B1(_06627_),
    .B2(_06628_),
    .ZN(_00137_));
 NAND2_X1 _16619_ (.A1(_06613_),
    .A2(\samples_imag[3][6] ),
    .ZN(_06629_));
 NAND2_X1 _16620_ (.A1(_06611_),
    .A2(net192),
    .ZN(_06630_));
 AOI21_X1 _16621_ (.A(_06620_),
    .B1(_06629_),
    .B2(_06630_),
    .ZN(_00138_));
 NAND2_X1 _16622_ (.A1(_06613_),
    .A2(\samples_imag[3][7] ),
    .ZN(_06631_));
 NAND2_X1 _16623_ (.A1(_06611_),
    .A2(net193),
    .ZN(_06632_));
 AOI21_X1 _16624_ (.A(_06620_),
    .B1(_06631_),
    .B2(_06632_),
    .ZN(_00139_));
 NAND2_X1 _16625_ (.A1(_06613_),
    .A2(\samples_imag[3][8] ),
    .ZN(_06633_));
 CLKBUF_X3 _16626_ (.A(_06517_),
    .Z(_06634_));
 NAND2_X1 _16627_ (.A1(_06634_),
    .A2(net194),
    .ZN(_06635_));
 AOI21_X1 _16628_ (.A(_06620_),
    .B1(_06633_),
    .B2(_06635_),
    .ZN(_00140_));
 BUF_X2 _16629_ (.A(_06520_),
    .Z(_06636_));
 NAND2_X1 _16630_ (.A1(_06636_),
    .A2(\samples_imag[3][9] ),
    .ZN(_06637_));
 NAND2_X1 _16631_ (.A1(_06634_),
    .A2(net195),
    .ZN(_06638_));
 AOI21_X1 _16632_ (.A(_06620_),
    .B1(_06637_),
    .B2(_06638_),
    .ZN(_00141_));
 NAND2_X1 _16633_ (.A1(_06636_),
    .A2(\samples_imag[3][10] ),
    .ZN(_06639_));
 NAND2_X1 _16634_ (.A1(_06634_),
    .A2(net196),
    .ZN(_06640_));
 AOI21_X1 _16635_ (.A(_06620_),
    .B1(_06639_),
    .B2(_06640_),
    .ZN(_00142_));
 NAND2_X1 _16636_ (.A1(_06636_),
    .A2(\samples_imag[3][11] ),
    .ZN(_06641_));
 NAND2_X1 _16637_ (.A1(_06634_),
    .A2(net197),
    .ZN(_06642_));
 AOI21_X1 _16638_ (.A(_06620_),
    .B1(_06641_),
    .B2(_06642_),
    .ZN(_00143_));
 CLKBUF_X3 _16639_ (.A(_06502_),
    .Z(_06643_));
 NAND2_X1 _16640_ (.A1(_06636_),
    .A2(\samples_imag[0][5] ),
    .ZN(_06644_));
 NAND2_X1 _16641_ (.A1(_06634_),
    .A2(net198),
    .ZN(_06645_));
 AOI21_X1 _16642_ (.A(_06643_),
    .B1(_06644_),
    .B2(_06645_),
    .ZN(_00144_));
 NAND2_X1 _16643_ (.A1(_06636_),
    .A2(\samples_imag[3][12] ),
    .ZN(_06646_));
 NAND2_X1 _16644_ (.A1(_06634_),
    .A2(net199),
    .ZN(_06647_));
 AOI21_X1 _16645_ (.A(_06643_),
    .B1(_06646_),
    .B2(_06647_),
    .ZN(_00145_));
 NAND2_X1 _16646_ (.A1(_06636_),
    .A2(\samples_imag[3][13] ),
    .ZN(_06648_));
 NAND2_X1 _16647_ (.A1(_06634_),
    .A2(net200),
    .ZN(_06649_));
 AOI21_X1 _16648_ (.A(_06643_),
    .B1(_06648_),
    .B2(_06649_),
    .ZN(_00146_));
 NAND2_X1 _16649_ (.A1(_06636_),
    .A2(\samples_imag[3][14] ),
    .ZN(_06650_));
 NAND2_X1 _16650_ (.A1(_06634_),
    .A2(net201),
    .ZN(_06651_));
 AOI21_X1 _16651_ (.A(_06643_),
    .B1(_06650_),
    .B2(_06651_),
    .ZN(_00147_));
 NAND2_X1 _16652_ (.A1(_06636_),
    .A2(\samples_imag[3][15] ),
    .ZN(_06652_));
 NAND2_X1 _16653_ (.A1(_06634_),
    .A2(net202),
    .ZN(_06653_));
 AOI21_X1 _16654_ (.A(_06643_),
    .B1(_06652_),
    .B2(_06653_),
    .ZN(_00148_));
 NAND2_X1 _16655_ (.A1(_06636_),
    .A2(\samples_imag[4][0] ),
    .ZN(_06654_));
 NAND2_X1 _16656_ (.A1(_06634_),
    .A2(net203),
    .ZN(_06655_));
 AOI21_X1 _16657_ (.A(_06643_),
    .B1(_06654_),
    .B2(_06655_),
    .ZN(_00149_));
 NAND2_X1 _16658_ (.A1(_06636_),
    .A2(\samples_imag[4][1] ),
    .ZN(_06656_));
 CLKBUF_X3 _16659_ (.A(_06517_),
    .Z(_06657_));
 NAND2_X1 _16660_ (.A1(_06657_),
    .A2(net204),
    .ZN(_06658_));
 AOI21_X1 _16661_ (.A(_06643_),
    .B1(_06656_),
    .B2(_06658_),
    .ZN(_00150_));
 BUF_X2 _16662_ (.A(_06520_),
    .Z(_06659_));
 NAND2_X1 _16663_ (.A1(_06659_),
    .A2(\samples_imag[4][2] ),
    .ZN(_06660_));
 NAND2_X1 _16664_ (.A1(_06657_),
    .A2(net205),
    .ZN(_06661_));
 AOI21_X1 _16665_ (.A(_06643_),
    .B1(_06660_),
    .B2(_06661_),
    .ZN(_00151_));
 NAND2_X1 _16666_ (.A1(_06659_),
    .A2(\samples_imag[4][3] ),
    .ZN(_06662_));
 NAND2_X1 _16667_ (.A1(_06657_),
    .A2(net206),
    .ZN(_06663_));
 AOI21_X1 _16668_ (.A(_06643_),
    .B1(_06662_),
    .B2(_06663_),
    .ZN(_00152_));
 NAND2_X1 _16669_ (.A1(_06659_),
    .A2(\samples_imag[4][4] ),
    .ZN(_06664_));
 NAND2_X1 _16670_ (.A1(_06657_),
    .A2(net207),
    .ZN(_06665_));
 AOI21_X1 _16671_ (.A(_06643_),
    .B1(_06664_),
    .B2(_06665_),
    .ZN(_00153_));
 CLKBUF_X3 _16672_ (.A(_06502_),
    .Z(_06666_));
 NAND2_X1 _16673_ (.A1(_06659_),
    .A2(\samples_imag[4][5] ),
    .ZN(_06667_));
 NAND2_X1 _16674_ (.A1(_06657_),
    .A2(net208),
    .ZN(_06668_));
 AOI21_X1 _16675_ (.A(_06666_),
    .B1(_06667_),
    .B2(_06668_),
    .ZN(_00154_));
 NAND2_X1 _16676_ (.A1(_06659_),
    .A2(\samples_imag[0][6] ),
    .ZN(_06669_));
 NAND2_X1 _16677_ (.A1(_06657_),
    .A2(net209),
    .ZN(_06670_));
 AOI21_X1 _16678_ (.A(_06666_),
    .B1(_06669_),
    .B2(_06670_),
    .ZN(_00155_));
 NAND2_X1 _16679_ (.A1(_06659_),
    .A2(\samples_imag[4][6] ),
    .ZN(_06671_));
 NAND2_X1 _16680_ (.A1(_06657_),
    .A2(net210),
    .ZN(_06672_));
 AOI21_X1 _16681_ (.A(_06666_),
    .B1(_06671_),
    .B2(_06672_),
    .ZN(_00156_));
 NAND2_X1 _16682_ (.A1(_06659_),
    .A2(\samples_imag[4][7] ),
    .ZN(_06673_));
 NAND2_X1 _16683_ (.A1(_06657_),
    .A2(net211),
    .ZN(_06674_));
 AOI21_X1 _16684_ (.A(_06666_),
    .B1(_06673_),
    .B2(_06674_),
    .ZN(_00157_));
 NAND2_X1 _16685_ (.A1(_06659_),
    .A2(\samples_imag[4][8] ),
    .ZN(_06675_));
 NAND2_X1 _16686_ (.A1(_06657_),
    .A2(net212),
    .ZN(_06676_));
 AOI21_X1 _16687_ (.A(_06666_),
    .B1(_06675_),
    .B2(_06676_),
    .ZN(_00158_));
 NAND2_X1 _16688_ (.A1(_06659_),
    .A2(\samples_imag[4][9] ),
    .ZN(_06677_));
 NAND2_X1 _16689_ (.A1(_06657_),
    .A2(net213),
    .ZN(_06678_));
 AOI21_X1 _16690_ (.A(_06666_),
    .B1(_06677_),
    .B2(_06678_),
    .ZN(_00159_));
 NAND2_X1 _16691_ (.A1(_06659_),
    .A2(\samples_imag[4][10] ),
    .ZN(_06679_));
 CLKBUF_X3 _16692_ (.A(_06517_),
    .Z(_06680_));
 NAND2_X1 _16693_ (.A1(_06680_),
    .A2(net214),
    .ZN(_06681_));
 AOI21_X1 _16694_ (.A(_06666_),
    .B1(_06679_),
    .B2(_06681_),
    .ZN(_00160_));
 BUF_X2 _16695_ (.A(_06520_),
    .Z(_06682_));
 NAND2_X1 _16696_ (.A1(_06682_),
    .A2(\samples_imag[4][11] ),
    .ZN(_06683_));
 NAND2_X1 _16697_ (.A1(_06680_),
    .A2(net215),
    .ZN(_06684_));
 AOI21_X1 _16698_ (.A(_06666_),
    .B1(_06683_),
    .B2(_06684_),
    .ZN(_00161_));
 NAND2_X1 _16699_ (.A1(_06682_),
    .A2(\samples_imag[4][12] ),
    .ZN(_06685_));
 NAND2_X1 _16700_ (.A1(_06680_),
    .A2(net216),
    .ZN(_06686_));
 AOI21_X1 _16701_ (.A(_06666_),
    .B1(_06685_),
    .B2(_06686_),
    .ZN(_00162_));
 NAND2_X1 _16702_ (.A1(_06682_),
    .A2(\samples_imag[4][13] ),
    .ZN(_06687_));
 NAND2_X1 _16703_ (.A1(_06680_),
    .A2(net217),
    .ZN(_06688_));
 AOI21_X1 _16704_ (.A(_06666_),
    .B1(_06687_),
    .B2(_06688_),
    .ZN(_00163_));
 CLKBUF_X3 _16705_ (.A(_06502_),
    .Z(_06689_));
 NAND2_X1 _16706_ (.A1(_06682_),
    .A2(\samples_imag[4][14] ),
    .ZN(_06690_));
 NAND2_X1 _16707_ (.A1(_06680_),
    .A2(net218),
    .ZN(_06691_));
 AOI21_X1 _16708_ (.A(_06689_),
    .B1(_06690_),
    .B2(_06691_),
    .ZN(_00164_));
 NAND2_X1 _16709_ (.A1(_06682_),
    .A2(\samples_imag[4][15] ),
    .ZN(_06692_));
 NAND2_X1 _16710_ (.A1(_06680_),
    .A2(net219),
    .ZN(_06693_));
 AOI21_X1 _16711_ (.A(_06689_),
    .B1(_06692_),
    .B2(_06693_),
    .ZN(_00165_));
 NAND2_X1 _16712_ (.A1(_06682_),
    .A2(\samples_imag[0][7] ),
    .ZN(_06694_));
 NAND2_X1 _16713_ (.A1(_06680_),
    .A2(net220),
    .ZN(_06695_));
 AOI21_X1 _16714_ (.A(_06689_),
    .B1(_06694_),
    .B2(_06695_),
    .ZN(_00166_));
 NAND2_X1 _16715_ (.A1(_06682_),
    .A2(\samples_imag[5][0] ),
    .ZN(_06696_));
 NAND2_X1 _16716_ (.A1(_06680_),
    .A2(net221),
    .ZN(_06697_));
 AOI21_X1 _16717_ (.A(_06689_),
    .B1(_06696_),
    .B2(_06697_),
    .ZN(_00167_));
 NAND2_X1 _16718_ (.A1(_06682_),
    .A2(\samples_imag[5][1] ),
    .ZN(_06698_));
 NAND2_X1 _16719_ (.A1(_06680_),
    .A2(net222),
    .ZN(_06699_));
 AOI21_X1 _16720_ (.A(_06689_),
    .B1(_06698_),
    .B2(_06699_),
    .ZN(_00168_));
 NAND2_X1 _16721_ (.A1(_06682_),
    .A2(\samples_imag[5][2] ),
    .ZN(_06700_));
 NAND2_X1 _16722_ (.A1(_06680_),
    .A2(net223),
    .ZN(_06701_));
 AOI21_X1 _16723_ (.A(_06689_),
    .B1(_06700_),
    .B2(_06701_),
    .ZN(_00169_));
 NAND2_X1 _16724_ (.A1(_06682_),
    .A2(\samples_imag[5][3] ),
    .ZN(_06702_));
 BUF_X2 _16725_ (.A(_06517_),
    .Z(_06703_));
 NAND2_X1 _16726_ (.A1(_06703_),
    .A2(net224),
    .ZN(_06704_));
 AOI21_X1 _16727_ (.A(_06689_),
    .B1(_06702_),
    .B2(_06704_),
    .ZN(_00170_));
 BUF_X2 _16728_ (.A(_06520_),
    .Z(_06705_));
 NAND2_X1 _16729_ (.A1(_06705_),
    .A2(\samples_imag[5][4] ),
    .ZN(_06706_));
 NAND2_X1 _16730_ (.A1(_06703_),
    .A2(net225),
    .ZN(_06707_));
 AOI21_X1 _16731_ (.A(_06689_),
    .B1(_06706_),
    .B2(_06707_),
    .ZN(_00171_));
 NAND2_X1 _16732_ (.A1(_06705_),
    .A2(\samples_imag[5][5] ),
    .ZN(_06708_));
 NAND2_X1 _16733_ (.A1(_06703_),
    .A2(net226),
    .ZN(_06709_));
 AOI21_X1 _16734_ (.A(_06689_),
    .B1(_06708_),
    .B2(_06709_),
    .ZN(_00172_));
 NAND2_X1 _16735_ (.A1(_06705_),
    .A2(\samples_imag[5][6] ),
    .ZN(_06710_));
 NAND2_X1 _16736_ (.A1(_06703_),
    .A2(net227),
    .ZN(_06711_));
 AOI21_X1 _16737_ (.A(_06689_),
    .B1(_06710_),
    .B2(_06711_),
    .ZN(_00173_));
 BUF_X2 _16738_ (.A(_06502_),
    .Z(_06712_));
 NAND2_X1 _16739_ (.A1(_06705_),
    .A2(\samples_imag[5][7] ),
    .ZN(_06713_));
 NAND2_X1 _16740_ (.A1(_06703_),
    .A2(net228),
    .ZN(_06714_));
 AOI21_X1 _16741_ (.A(_06712_),
    .B1(_06713_),
    .B2(_06714_),
    .ZN(_00174_));
 NAND2_X1 _16742_ (.A1(_06705_),
    .A2(\samples_imag[5][8] ),
    .ZN(_06715_));
 NAND2_X1 _16743_ (.A1(_06703_),
    .A2(net229),
    .ZN(_06716_));
 AOI21_X1 _16744_ (.A(_06712_),
    .B1(_06715_),
    .B2(_06716_),
    .ZN(_00175_));
 NAND2_X1 _16745_ (.A1(_06705_),
    .A2(\samples_imag[5][9] ),
    .ZN(_06717_));
 NAND2_X1 _16746_ (.A1(_06703_),
    .A2(net230),
    .ZN(_06718_));
 AOI21_X1 _16747_ (.A(_06712_),
    .B1(_06717_),
    .B2(_06718_),
    .ZN(_00176_));
 NAND2_X1 _16748_ (.A1(_06705_),
    .A2(\samples_imag[0][8] ),
    .ZN(_06719_));
 NAND2_X1 _16749_ (.A1(_06703_),
    .A2(net231),
    .ZN(_06720_));
 AOI21_X1 _16750_ (.A(_06712_),
    .B1(_06719_),
    .B2(_06720_),
    .ZN(_00177_));
 NAND2_X1 _16751_ (.A1(_06705_),
    .A2(\samples_imag[5][10] ),
    .ZN(_06721_));
 NAND2_X1 _16752_ (.A1(_06703_),
    .A2(net232),
    .ZN(_06722_));
 AOI21_X1 _16753_ (.A(_06712_),
    .B1(_06721_),
    .B2(_06722_),
    .ZN(_00178_));
 NAND2_X1 _16754_ (.A1(_06705_),
    .A2(\samples_imag[5][11] ),
    .ZN(_06723_));
 NAND2_X1 _16755_ (.A1(_06703_),
    .A2(net233),
    .ZN(_06724_));
 AOI21_X1 _16756_ (.A(_06712_),
    .B1(_06723_),
    .B2(_06724_),
    .ZN(_00179_));
 NAND2_X1 _16757_ (.A1(_06705_),
    .A2(\samples_imag[5][12] ),
    .ZN(_06725_));
 CLKBUF_X3 _16758_ (.A(_06517_),
    .Z(_06726_));
 NAND2_X1 _16759_ (.A1(_06726_),
    .A2(net234),
    .ZN(_06727_));
 AOI21_X1 _16760_ (.A(_06712_),
    .B1(_06725_),
    .B2(_06727_),
    .ZN(_00180_));
 BUF_X4 _16761_ (.A(_06520_),
    .Z(_06728_));
 NAND2_X1 _16762_ (.A1(_06728_),
    .A2(\samples_imag[5][13] ),
    .ZN(_06729_));
 NAND2_X1 _16763_ (.A1(_06726_),
    .A2(net235),
    .ZN(_06730_));
 AOI21_X1 _16764_ (.A(_06712_),
    .B1(_06729_),
    .B2(_06730_),
    .ZN(_00181_));
 NAND2_X1 _16765_ (.A1(_06728_),
    .A2(\samples_imag[5][14] ),
    .ZN(_06731_));
 NAND2_X1 _16766_ (.A1(_06726_),
    .A2(net236),
    .ZN(_06732_));
 AOI21_X1 _16767_ (.A(_06712_),
    .B1(_06731_),
    .B2(_06732_),
    .ZN(_00182_));
 NAND2_X1 _16768_ (.A1(_06728_),
    .A2(\samples_imag[5][15] ),
    .ZN(_06733_));
 NAND2_X1 _16769_ (.A1(_06726_),
    .A2(net237),
    .ZN(_06734_));
 AOI21_X1 _16770_ (.A(_06712_),
    .B1(_06733_),
    .B2(_06734_),
    .ZN(_00183_));
 CLKBUF_X3 _16771_ (.A(_00843_),
    .Z(_06735_));
 BUF_X4 _16772_ (.A(_06735_),
    .Z(_06736_));
 NAND2_X1 _16773_ (.A1(_06728_),
    .A2(\samples_imag[6][0] ),
    .ZN(_06737_));
 NAND2_X1 _16774_ (.A1(_06726_),
    .A2(net238),
    .ZN(_06738_));
 AOI21_X1 _16775_ (.A(_06736_),
    .B1(_06737_),
    .B2(_06738_),
    .ZN(_00184_));
 NAND2_X1 _16776_ (.A1(_06728_),
    .A2(\samples_imag[6][1] ),
    .ZN(_06739_));
 NAND2_X1 _16777_ (.A1(_06726_),
    .A2(net239),
    .ZN(_06740_));
 AOI21_X1 _16778_ (.A(_06736_),
    .B1(_06739_),
    .B2(_06740_),
    .ZN(_00185_));
 NAND2_X1 _16779_ (.A1(_06728_),
    .A2(\samples_imag[6][2] ),
    .ZN(_06741_));
 NAND2_X1 _16780_ (.A1(_06726_),
    .A2(net240),
    .ZN(_06742_));
 AOI21_X1 _16781_ (.A(_06736_),
    .B1(_06741_),
    .B2(_06742_),
    .ZN(_00186_));
 NAND2_X1 _16782_ (.A1(_06728_),
    .A2(\samples_imag[6][3] ),
    .ZN(_06743_));
 NAND2_X1 _16783_ (.A1(_06726_),
    .A2(net241),
    .ZN(_06744_));
 AOI21_X1 _16784_ (.A(_06736_),
    .B1(_06743_),
    .B2(_06744_),
    .ZN(_00187_));
 NAND2_X1 _16785_ (.A1(_06728_),
    .A2(\samples_imag[0][9] ),
    .ZN(_06745_));
 NAND2_X1 _16786_ (.A1(_06726_),
    .A2(net242),
    .ZN(_06746_));
 AOI21_X1 _16787_ (.A(_06736_),
    .B1(_06745_),
    .B2(_06746_),
    .ZN(_00188_));
 NAND2_X1 _16788_ (.A1(_06728_),
    .A2(\samples_real[0][0] ),
    .ZN(_06747_));
 NAND2_X1 _16789_ (.A1(_06726_),
    .A2(net243),
    .ZN(_06748_));
 AOI21_X1 _16790_ (.A(_06736_),
    .B1(_06747_),
    .B2(_06748_),
    .ZN(_00189_));
 NAND2_X1 _16791_ (.A1(_06728_),
    .A2(\samples_real[6][4] ),
    .ZN(_06749_));
 CLKBUF_X3 _16792_ (.A(_00858_),
    .Z(_06750_));
 CLKBUF_X3 _16793_ (.A(_06750_),
    .Z(_06751_));
 NAND2_X1 _16794_ (.A1(_06751_),
    .A2(net244),
    .ZN(_06752_));
 AOI21_X1 _16795_ (.A(_06736_),
    .B1(_06749_),
    .B2(_06752_),
    .ZN(_00190_));
 CLKBUF_X3 _16796_ (.A(_00857_),
    .Z(_06753_));
 BUF_X2 _16797_ (.A(_06753_),
    .Z(_06754_));
 NAND2_X1 _16798_ (.A1(_06754_),
    .A2(\samples_real[6][5] ),
    .ZN(_06755_));
 NAND2_X1 _16799_ (.A1(_06751_),
    .A2(net245),
    .ZN(_06756_));
 AOI21_X1 _16800_ (.A(_06736_),
    .B1(_06755_),
    .B2(_06756_),
    .ZN(_00191_));
 NAND2_X1 _16801_ (.A1(_06754_),
    .A2(\samples_real[6][6] ),
    .ZN(_06757_));
 NAND2_X1 _16802_ (.A1(_06751_),
    .A2(net246),
    .ZN(_06758_));
 AOI21_X1 _16803_ (.A(_06736_),
    .B1(_06757_),
    .B2(_06758_),
    .ZN(_00192_));
 NAND2_X1 _16804_ (.A1(_06754_),
    .A2(\samples_real[6][7] ),
    .ZN(_06759_));
 NAND2_X1 _16805_ (.A1(_06751_),
    .A2(net247),
    .ZN(_06760_));
 AOI21_X1 _16806_ (.A(_06736_),
    .B1(_06759_),
    .B2(_06760_),
    .ZN(_00193_));
 CLKBUF_X3 _16807_ (.A(_06735_),
    .Z(_06761_));
 NAND2_X1 _16808_ (.A1(_06754_),
    .A2(\samples_real[6][8] ),
    .ZN(_06762_));
 NAND2_X1 _16809_ (.A1(_06751_),
    .A2(net248),
    .ZN(_06763_));
 AOI21_X1 _16810_ (.A(_06761_),
    .B1(_06762_),
    .B2(_06763_),
    .ZN(_00194_));
 NAND2_X1 _16811_ (.A1(_06754_),
    .A2(\samples_real[6][9] ),
    .ZN(_06764_));
 NAND2_X1 _16812_ (.A1(_06751_),
    .A2(net249),
    .ZN(_06765_));
 AOI21_X1 _16813_ (.A(_06761_),
    .B1(_06764_),
    .B2(_06765_),
    .ZN(_00195_));
 NAND2_X1 _16814_ (.A1(_06754_),
    .A2(\samples_real[6][10] ),
    .ZN(_06766_));
 NAND2_X1 _16815_ (.A1(_06751_),
    .A2(net250),
    .ZN(_06767_));
 AOI21_X1 _16816_ (.A(_06761_),
    .B1(_06766_),
    .B2(_06767_),
    .ZN(_00196_));
 NAND2_X1 _16817_ (.A1(_06754_),
    .A2(\samples_real[6][11] ),
    .ZN(_06768_));
 NAND2_X1 _16818_ (.A1(_06751_),
    .A2(net251),
    .ZN(_06769_));
 AOI21_X1 _16819_ (.A(_06761_),
    .B1(_06768_),
    .B2(_06769_),
    .ZN(_00197_));
 NAND2_X1 _16820_ (.A1(_06754_),
    .A2(\samples_real[6][12] ),
    .ZN(_06770_));
 NAND2_X1 _16821_ (.A1(_06751_),
    .A2(net252),
    .ZN(_06771_));
 AOI21_X1 _16822_ (.A(_06761_),
    .B1(_06770_),
    .B2(_06771_),
    .ZN(_00198_));
 NAND2_X1 _16823_ (.A1(_06754_),
    .A2(\samples_real[6][13] ),
    .ZN(_06772_));
 NAND2_X1 _16824_ (.A1(_06751_),
    .A2(net253),
    .ZN(_06773_));
 AOI21_X1 _16825_ (.A(_06761_),
    .B1(_06772_),
    .B2(_06773_),
    .ZN(_00199_));
 NAND2_X1 _16826_ (.A1(_06754_),
    .A2(\samples_real[0][10] ),
    .ZN(_06774_));
 CLKBUF_X3 _16827_ (.A(_06750_),
    .Z(_06775_));
 NAND2_X1 _16828_ (.A1(_06775_),
    .A2(net254),
    .ZN(_06776_));
 AOI21_X1 _16829_ (.A(_06761_),
    .B1(_06774_),
    .B2(_06776_),
    .ZN(_00200_));
 BUF_X2 _16830_ (.A(_06753_),
    .Z(_06777_));
 NAND2_X1 _16831_ (.A1(_06777_),
    .A2(\samples_real[6][14] ),
    .ZN(_06778_));
 NAND2_X1 _16832_ (.A1(_06775_),
    .A2(net255),
    .ZN(_06779_));
 AOI21_X1 _16833_ (.A(_06761_),
    .B1(_06778_),
    .B2(_06779_),
    .ZN(_00201_));
 NAND2_X1 _16834_ (.A1(_06777_),
    .A2(\samples_real[6][15] ),
    .ZN(_06780_));
 NAND2_X1 _16835_ (.A1(_06775_),
    .A2(net256),
    .ZN(_06781_));
 AOI21_X1 _16836_ (.A(_06761_),
    .B1(_06780_),
    .B2(_06781_),
    .ZN(_00202_));
 NAND2_X1 _16837_ (.A1(_06777_),
    .A2(\samples_real[7][0] ),
    .ZN(_06782_));
 NAND2_X1 _16838_ (.A1(_06775_),
    .A2(net257),
    .ZN(_06783_));
 AOI21_X1 _16839_ (.A(_06761_),
    .B1(_06782_),
    .B2(_06783_),
    .ZN(_00203_));
 CLKBUF_X3 _16840_ (.A(_06735_),
    .Z(_06784_));
 NAND2_X1 _16841_ (.A1(_06777_),
    .A2(\samples_real[7][1] ),
    .ZN(_06785_));
 NAND2_X1 _16842_ (.A1(_06775_),
    .A2(net258),
    .ZN(_06786_));
 AOI21_X1 _16843_ (.A(_06784_),
    .B1(_06785_),
    .B2(_06786_),
    .ZN(_00204_));
 NAND2_X1 _16844_ (.A1(_06777_),
    .A2(\samples_real[7][2] ),
    .ZN(_06787_));
 NAND2_X1 _16845_ (.A1(_06775_),
    .A2(net259),
    .ZN(_06788_));
 AOI21_X1 _16846_ (.A(_06784_),
    .B1(_06787_),
    .B2(_06788_),
    .ZN(_00205_));
 NAND2_X1 _16847_ (.A1(_06777_),
    .A2(\samples_real[7][3] ),
    .ZN(_06789_));
 NAND2_X1 _16848_ (.A1(_06775_),
    .A2(net260),
    .ZN(_06790_));
 AOI21_X1 _16849_ (.A(_06784_),
    .B1(_06789_),
    .B2(_06790_),
    .ZN(_00206_));
 NAND2_X1 _16850_ (.A1(_06777_),
    .A2(\samples_real[7][4] ),
    .ZN(_06791_));
 NAND2_X1 _16851_ (.A1(_06775_),
    .A2(net261),
    .ZN(_06792_));
 AOI21_X1 _16852_ (.A(_06784_),
    .B1(_06791_),
    .B2(_06792_),
    .ZN(_00207_));
 NAND2_X1 _16853_ (.A1(_06777_),
    .A2(\samples_real[7][5] ),
    .ZN(_06793_));
 NAND2_X1 _16854_ (.A1(_06775_),
    .A2(net262),
    .ZN(_06794_));
 AOI21_X1 _16855_ (.A(_06784_),
    .B1(_06793_),
    .B2(_06794_),
    .ZN(_00208_));
 NAND2_X1 _16856_ (.A1(_06777_),
    .A2(\samples_real[7][6] ),
    .ZN(_06795_));
 NAND2_X1 _16857_ (.A1(_06775_),
    .A2(net263),
    .ZN(_06796_));
 AOI21_X1 _16858_ (.A(_06784_),
    .B1(_06795_),
    .B2(_06796_),
    .ZN(_00209_));
 NAND2_X1 _16859_ (.A1(_06777_),
    .A2(\samples_real[7][7] ),
    .ZN(_06797_));
 CLKBUF_X3 _16860_ (.A(_06750_),
    .Z(_06798_));
 NAND2_X1 _16861_ (.A1(_06798_),
    .A2(net264),
    .ZN(_06799_));
 AOI21_X1 _16862_ (.A(_06784_),
    .B1(_06797_),
    .B2(_06799_),
    .ZN(_00210_));
 BUF_X2 _16863_ (.A(_06753_),
    .Z(_06800_));
 NAND2_X1 _16864_ (.A1(_06800_),
    .A2(\samples_real[0][11] ),
    .ZN(_06801_));
 NAND2_X1 _16865_ (.A1(_06798_),
    .A2(net265),
    .ZN(_06802_));
 AOI21_X1 _16866_ (.A(_06784_),
    .B1(_06801_),
    .B2(_06802_),
    .ZN(_00211_));
 NAND2_X1 _16867_ (.A1(_06800_),
    .A2(\samples_real[7][8] ),
    .ZN(_06803_));
 NAND2_X1 _16868_ (.A1(_06798_),
    .A2(net266),
    .ZN(_06804_));
 AOI21_X1 _16869_ (.A(_06784_),
    .B1(_06803_),
    .B2(_06804_),
    .ZN(_00212_));
 NAND2_X1 _16870_ (.A1(_06800_),
    .A2(\samples_real[7][9] ),
    .ZN(_06805_));
 NAND2_X1 _16871_ (.A1(_06798_),
    .A2(net267),
    .ZN(_06806_));
 AOI21_X1 _16872_ (.A(_06784_),
    .B1(_06805_),
    .B2(_06806_),
    .ZN(_00213_));
 CLKBUF_X3 _16873_ (.A(_06735_),
    .Z(_06807_));
 NAND2_X1 _16874_ (.A1(_06800_),
    .A2(\samples_real[7][10] ),
    .ZN(_06808_));
 NAND2_X1 _16875_ (.A1(_06798_),
    .A2(net268),
    .ZN(_06809_));
 AOI21_X1 _16876_ (.A(_06807_),
    .B1(_06808_),
    .B2(_06809_),
    .ZN(_00214_));
 NAND2_X1 _16877_ (.A1(_06800_),
    .A2(\samples_real[7][11] ),
    .ZN(_06810_));
 NAND2_X1 _16878_ (.A1(_06798_),
    .A2(net269),
    .ZN(_06811_));
 AOI21_X1 _16879_ (.A(_06807_),
    .B1(_06810_),
    .B2(_06811_),
    .ZN(_00215_));
 NAND2_X1 _16880_ (.A1(_06800_),
    .A2(\samples_real[7][12] ),
    .ZN(_06812_));
 NAND2_X1 _16881_ (.A1(_06798_),
    .A2(net270),
    .ZN(_00586_));
 AOI21_X1 _16882_ (.A(_06807_),
    .B1(_06812_),
    .B2(_00586_),
    .ZN(_00216_));
 NAND2_X1 _16883_ (.A1(_06800_),
    .A2(\samples_real[7][13] ),
    .ZN(_00587_));
 NAND2_X1 _16884_ (.A1(_06798_),
    .A2(net271),
    .ZN(_00588_));
 AOI21_X1 _16885_ (.A(_06807_),
    .B1(_00587_),
    .B2(_00588_),
    .ZN(_00217_));
 NAND2_X1 _16886_ (.A1(_06800_),
    .A2(\samples_real[7][14] ),
    .ZN(_00589_));
 NAND2_X1 _16887_ (.A1(_06798_),
    .A2(net272),
    .ZN(_00590_));
 AOI21_X1 _16888_ (.A(_06807_),
    .B1(_00589_),
    .B2(_00590_),
    .ZN(_00218_));
 NAND2_X1 _16889_ (.A1(_06800_),
    .A2(\samples_real[7][15] ),
    .ZN(_00591_));
 NAND2_X1 _16890_ (.A1(_06798_),
    .A2(net273),
    .ZN(_00592_));
 AOI21_X1 _16891_ (.A(_06807_),
    .B1(_00591_),
    .B2(_00592_),
    .ZN(_00219_));
 NAND2_X1 _16892_ (.A1(_06800_),
    .A2(\samples_real[0][12] ),
    .ZN(_00593_));
 CLKBUF_X3 _16893_ (.A(_06750_),
    .Z(_00594_));
 NAND2_X1 _16894_ (.A1(_00594_),
    .A2(net274),
    .ZN(_00595_));
 AOI21_X1 _16895_ (.A(_06807_),
    .B1(_00593_),
    .B2(_00595_),
    .ZN(_00220_));
 BUF_X2 _16896_ (.A(_06753_),
    .Z(_00596_));
 NAND2_X1 _16897_ (.A1(_00596_),
    .A2(\samples_real[0][13] ),
    .ZN(_00597_));
 NAND2_X1 _16898_ (.A1(_00594_),
    .A2(net275),
    .ZN(_00598_));
 AOI21_X1 _16899_ (.A(_06807_),
    .B1(_00597_),
    .B2(_00598_),
    .ZN(_00221_));
 NAND2_X1 _16900_ (.A1(_00596_),
    .A2(\samples_real[0][14] ),
    .ZN(_00599_));
 NAND2_X1 _16901_ (.A1(_00594_),
    .A2(net276),
    .ZN(_00600_));
 AOI21_X1 _16902_ (.A(_06807_),
    .B1(_00599_),
    .B2(_00600_),
    .ZN(_00222_));
 NAND2_X1 _16903_ (.A1(_00596_),
    .A2(\samples_real[0][15] ),
    .ZN(_00601_));
 NAND2_X1 _16904_ (.A1(_00594_),
    .A2(net277),
    .ZN(_00602_));
 AOI21_X1 _16905_ (.A(_06807_),
    .B1(_00601_),
    .B2(_00602_),
    .ZN(_00223_));
 CLKBUF_X3 _16906_ (.A(_06735_),
    .Z(_00603_));
 NAND2_X1 _16907_ (.A1(_00596_),
    .A2(\samples_real[1][0] ),
    .ZN(_00604_));
 NAND2_X1 _16908_ (.A1(_00594_),
    .A2(net278),
    .ZN(_00605_));
 AOI21_X1 _16909_ (.A(_00603_),
    .B1(_00604_),
    .B2(_00605_),
    .ZN(_00224_));
 NAND2_X1 _16910_ (.A1(_00596_),
    .A2(\samples_real[1][1] ),
    .ZN(_00606_));
 NAND2_X1 _16911_ (.A1(_00594_),
    .A2(net279),
    .ZN(_00607_));
 AOI21_X1 _16912_ (.A(_00603_),
    .B1(_00606_),
    .B2(_00607_),
    .ZN(_00225_));
 NAND2_X1 _16913_ (.A1(_00596_),
    .A2(\samples_real[1][2] ),
    .ZN(_00608_));
 NAND2_X1 _16914_ (.A1(_00594_),
    .A2(net280),
    .ZN(_00609_));
 AOI21_X1 _16915_ (.A(_00603_),
    .B1(_00608_),
    .B2(_00609_),
    .ZN(_00226_));
 NAND2_X1 _16916_ (.A1(_00596_),
    .A2(\samples_real[1][3] ),
    .ZN(_00610_));
 NAND2_X1 _16917_ (.A1(_00594_),
    .A2(net281),
    .ZN(_00611_));
 AOI21_X1 _16918_ (.A(_00603_),
    .B1(_00610_),
    .B2(_00611_),
    .ZN(_00227_));
 NAND2_X1 _16919_ (.A1(_00596_),
    .A2(\samples_real[0][1] ),
    .ZN(_00612_));
 NAND2_X1 _16920_ (.A1(_00594_),
    .A2(net282),
    .ZN(_00613_));
 AOI21_X1 _16921_ (.A(_00603_),
    .B1(_00612_),
    .B2(_00613_),
    .ZN(_00228_));
 NAND2_X1 _16922_ (.A1(_00596_),
    .A2(\samples_real[1][4] ),
    .ZN(_00614_));
 NAND2_X1 _16923_ (.A1(_00594_),
    .A2(net283),
    .ZN(_00615_));
 AOI21_X1 _16924_ (.A(_00603_),
    .B1(_00614_),
    .B2(_00615_),
    .ZN(_00229_));
 NAND2_X1 _16925_ (.A1(_00596_),
    .A2(\samples_real[1][5] ),
    .ZN(_00616_));
 CLKBUF_X3 _16926_ (.A(_06750_),
    .Z(_00617_));
 NAND2_X1 _16927_ (.A1(_00617_),
    .A2(net284),
    .ZN(_00618_));
 AOI21_X1 _16928_ (.A(_00603_),
    .B1(_00616_),
    .B2(_00618_),
    .ZN(_00230_));
 CLKBUF_X3 _16929_ (.A(_06753_),
    .Z(_00619_));
 NAND2_X1 _16930_ (.A1(_00619_),
    .A2(\samples_real[1][6] ),
    .ZN(_00620_));
 NAND2_X1 _16931_ (.A1(_00617_),
    .A2(net285),
    .ZN(_00621_));
 AOI21_X1 _16932_ (.A(_00603_),
    .B1(_00620_),
    .B2(_00621_),
    .ZN(_00231_));
 NAND2_X1 _16933_ (.A1(_00619_),
    .A2(\samples_real[1][7] ),
    .ZN(_00622_));
 NAND2_X1 _16934_ (.A1(_00617_),
    .A2(net286),
    .ZN(_00623_));
 AOI21_X1 _16935_ (.A(_00603_),
    .B1(_00622_),
    .B2(_00623_),
    .ZN(_00232_));
 NAND2_X1 _16936_ (.A1(_00619_),
    .A2(\samples_real[1][8] ),
    .ZN(_00624_));
 NAND2_X1 _16937_ (.A1(_00617_),
    .A2(net287),
    .ZN(_00625_));
 AOI21_X1 _16938_ (.A(_00603_),
    .B1(_00624_),
    .B2(_00625_),
    .ZN(_00233_));
 CLKBUF_X3 _16939_ (.A(_06735_),
    .Z(_00626_));
 NAND2_X1 _16940_ (.A1(_00619_),
    .A2(\samples_real[1][9] ),
    .ZN(_00627_));
 NAND2_X1 _16941_ (.A1(_00617_),
    .A2(net288),
    .ZN(_00628_));
 AOI21_X1 _16942_ (.A(_00626_),
    .B1(_00627_),
    .B2(_00628_),
    .ZN(_00234_));
 NAND2_X1 _16943_ (.A1(_00619_),
    .A2(\samples_real[1][10] ),
    .ZN(_00629_));
 NAND2_X1 _16944_ (.A1(_00617_),
    .A2(net289),
    .ZN(_00630_));
 AOI21_X1 _16945_ (.A(_00626_),
    .B1(_00629_),
    .B2(_00630_),
    .ZN(_00235_));
 NAND2_X1 _16946_ (.A1(_00619_),
    .A2(\samples_real[1][11] ),
    .ZN(_00631_));
 NAND2_X1 _16947_ (.A1(_00617_),
    .A2(net290),
    .ZN(_00632_));
 AOI21_X1 _16948_ (.A(_00626_),
    .B1(_00631_),
    .B2(_00632_),
    .ZN(_00236_));
 NAND2_X1 _16949_ (.A1(_00619_),
    .A2(\samples_real[1][12] ),
    .ZN(_00633_));
 NAND2_X1 _16950_ (.A1(_00617_),
    .A2(net291),
    .ZN(_00634_));
 AOI21_X1 _16951_ (.A(_00626_),
    .B1(_00633_),
    .B2(_00634_),
    .ZN(_00237_));
 NAND2_X1 _16952_ (.A1(_00619_),
    .A2(\samples_real[1][13] ),
    .ZN(_00635_));
 NAND2_X1 _16953_ (.A1(_00617_),
    .A2(net292),
    .ZN(_00636_));
 AOI21_X1 _16954_ (.A(_00626_),
    .B1(_00635_),
    .B2(_00636_),
    .ZN(_00238_));
 NAND2_X1 _16955_ (.A1(_00619_),
    .A2(\samples_real[0][2] ),
    .ZN(_00637_));
 NAND2_X1 _16956_ (.A1(_00617_),
    .A2(net293),
    .ZN(_00638_));
 AOI21_X1 _16957_ (.A(_00626_),
    .B1(_00637_),
    .B2(_00638_),
    .ZN(_00239_));
 NAND2_X1 _16958_ (.A1(_00619_),
    .A2(\samples_real[1][14] ),
    .ZN(_00639_));
 CLKBUF_X3 _16959_ (.A(_06750_),
    .Z(_00640_));
 NAND2_X1 _16960_ (.A1(_00640_),
    .A2(net294),
    .ZN(_00641_));
 AOI21_X1 _16961_ (.A(_00626_),
    .B1(_00639_),
    .B2(_00641_),
    .ZN(_00240_));
 CLKBUF_X3 _16962_ (.A(_06753_),
    .Z(_00642_));
 NAND2_X1 _16963_ (.A1(_00642_),
    .A2(\samples_real[1][15] ),
    .ZN(_00643_));
 NAND2_X1 _16964_ (.A1(_00640_),
    .A2(net295),
    .ZN(_00644_));
 AOI21_X1 _16965_ (.A(_00626_),
    .B1(_00643_),
    .B2(_00644_),
    .ZN(_00241_));
 NAND2_X1 _16966_ (.A1(_00642_),
    .A2(\samples_real[2][0] ),
    .ZN(_00645_));
 NAND2_X1 _16967_ (.A1(_00640_),
    .A2(net296),
    .ZN(_00646_));
 AOI21_X1 _16968_ (.A(_00626_),
    .B1(_00645_),
    .B2(_00646_),
    .ZN(_00242_));
 NAND2_X1 _16969_ (.A1(_00642_),
    .A2(\samples_real[2][1] ),
    .ZN(_00647_));
 NAND2_X1 _16970_ (.A1(_00640_),
    .A2(net297),
    .ZN(_00648_));
 AOI21_X1 _16971_ (.A(_00626_),
    .B1(_00647_),
    .B2(_00648_),
    .ZN(_00243_));
 CLKBUF_X3 _16972_ (.A(_06735_),
    .Z(_00649_));
 NAND2_X1 _16973_ (.A1(_00642_),
    .A2(\samples_real[2][2] ),
    .ZN(_00650_));
 NAND2_X1 _16974_ (.A1(_00640_),
    .A2(net298),
    .ZN(_00651_));
 AOI21_X1 _16975_ (.A(_00649_),
    .B1(_00650_),
    .B2(_00651_),
    .ZN(_00244_));
 NAND2_X1 _16976_ (.A1(_00642_),
    .A2(\samples_real[2][3] ),
    .ZN(_00652_));
 NAND2_X1 _16977_ (.A1(_00640_),
    .A2(net299),
    .ZN(_00653_));
 AOI21_X1 _16978_ (.A(_00649_),
    .B1(_00652_),
    .B2(_00653_),
    .ZN(_00245_));
 NAND2_X1 _16979_ (.A1(_00642_),
    .A2(\samples_real[2][4] ),
    .ZN(_00654_));
 NAND2_X1 _16980_ (.A1(_00640_),
    .A2(net300),
    .ZN(_00655_));
 AOI21_X1 _16981_ (.A(_00649_),
    .B1(_00654_),
    .B2(_00655_),
    .ZN(_00246_));
 NAND2_X1 _16982_ (.A1(_00642_),
    .A2(\samples_real[2][5] ),
    .ZN(_00656_));
 NAND2_X1 _16983_ (.A1(_00640_),
    .A2(net301),
    .ZN(_00657_));
 AOI21_X1 _16984_ (.A(_00649_),
    .B1(_00656_),
    .B2(_00657_),
    .ZN(_00247_));
 NAND2_X1 _16985_ (.A1(_00642_),
    .A2(\samples_real[2][6] ),
    .ZN(_00658_));
 NAND2_X1 _16986_ (.A1(_00640_),
    .A2(net302),
    .ZN(_00659_));
 AOI21_X1 _16987_ (.A(_00649_),
    .B1(_00658_),
    .B2(_00659_),
    .ZN(_00248_));
 NAND2_X1 _16988_ (.A1(_00642_),
    .A2(\samples_real[2][7] ),
    .ZN(_00660_));
 NAND2_X1 _16989_ (.A1(_00640_),
    .A2(net303),
    .ZN(_00661_));
 AOI21_X1 _16990_ (.A(_00649_),
    .B1(_00660_),
    .B2(_00661_),
    .ZN(_00249_));
 NAND2_X1 _16991_ (.A1(_00642_),
    .A2(\samples_real[0][3] ),
    .ZN(_00662_));
 CLKBUF_X3 _16992_ (.A(_06750_),
    .Z(_00663_));
 NAND2_X1 _16993_ (.A1(_00663_),
    .A2(net304),
    .ZN(_00664_));
 AOI21_X1 _16994_ (.A(_00649_),
    .B1(_00662_),
    .B2(_00664_),
    .ZN(_00250_));
 CLKBUF_X3 _16995_ (.A(_06753_),
    .Z(_00665_));
 NAND2_X1 _16996_ (.A1(_00665_),
    .A2(\samples_real[2][8] ),
    .ZN(_00666_));
 NAND2_X1 _16997_ (.A1(_00663_),
    .A2(net305),
    .ZN(_00667_));
 AOI21_X1 _16998_ (.A(_00649_),
    .B1(_00666_),
    .B2(_00667_),
    .ZN(_00251_));
 NAND2_X1 _16999_ (.A1(_00665_),
    .A2(\samples_real[2][9] ),
    .ZN(_00668_));
 NAND2_X1 _17000_ (.A1(_00663_),
    .A2(net306),
    .ZN(_00669_));
 AOI21_X1 _17001_ (.A(_00649_),
    .B1(_00668_),
    .B2(_00669_),
    .ZN(_00252_));
 NAND2_X1 _17002_ (.A1(_00665_),
    .A2(\samples_real[2][10] ),
    .ZN(_00670_));
 NAND2_X1 _17003_ (.A1(_00663_),
    .A2(net307),
    .ZN(_00671_));
 AOI21_X1 _17004_ (.A(_00649_),
    .B1(_00670_),
    .B2(_00671_),
    .ZN(_00253_));
 CLKBUF_X3 _17005_ (.A(_06735_),
    .Z(_00672_));
 NAND2_X1 _17006_ (.A1(_00665_),
    .A2(\samples_real[2][11] ),
    .ZN(_00673_));
 NAND2_X1 _17007_ (.A1(_00663_),
    .A2(net308),
    .ZN(_00674_));
 AOI21_X1 _17008_ (.A(_00672_),
    .B1(_00673_),
    .B2(_00674_),
    .ZN(_00254_));
 NAND2_X1 _17009_ (.A1(_00665_),
    .A2(\samples_real[2][12] ),
    .ZN(_00675_));
 NAND2_X1 _17010_ (.A1(_00663_),
    .A2(net309),
    .ZN(_00676_));
 AOI21_X1 _17011_ (.A(_00672_),
    .B1(_00675_),
    .B2(_00676_),
    .ZN(_00255_));
 NAND2_X1 _17012_ (.A1(_00665_),
    .A2(\samples_real[2][13] ),
    .ZN(_00677_));
 NAND2_X1 _17013_ (.A1(_00663_),
    .A2(net310),
    .ZN(_00678_));
 AOI21_X1 _17014_ (.A(_00672_),
    .B1(_00677_),
    .B2(_00678_),
    .ZN(_00256_));
 NAND2_X1 _17015_ (.A1(_00665_),
    .A2(\samples_real[2][14] ),
    .ZN(_00679_));
 NAND2_X1 _17016_ (.A1(_00663_),
    .A2(net311),
    .ZN(_00680_));
 AOI21_X1 _17017_ (.A(_00672_),
    .B1(_00679_),
    .B2(_00680_),
    .ZN(_00257_));
 NAND2_X1 _17018_ (.A1(_00665_),
    .A2(\samples_real[2][15] ),
    .ZN(_00681_));
 NAND2_X1 _17019_ (.A1(_00663_),
    .A2(net312),
    .ZN(_00682_));
 AOI21_X1 _17020_ (.A(_00672_),
    .B1(_00681_),
    .B2(_00682_),
    .ZN(_00258_));
 NAND2_X1 _17021_ (.A1(_00665_),
    .A2(\samples_real[3][0] ),
    .ZN(_00683_));
 NAND2_X1 _17022_ (.A1(_00663_),
    .A2(net313),
    .ZN(_00684_));
 AOI21_X1 _17023_ (.A(_00672_),
    .B1(_00683_),
    .B2(_00684_),
    .ZN(_00259_));
 NAND2_X1 _17024_ (.A1(_00665_),
    .A2(\samples_real[3][1] ),
    .ZN(_00685_));
 CLKBUF_X3 _17025_ (.A(_06750_),
    .Z(_00686_));
 NAND2_X1 _17026_ (.A1(_00686_),
    .A2(net314),
    .ZN(_00687_));
 AOI21_X1 _17027_ (.A(_00672_),
    .B1(_00685_),
    .B2(_00687_),
    .ZN(_00260_));
 BUF_X2 _17028_ (.A(_06753_),
    .Z(_00688_));
 NAND2_X1 _17029_ (.A1(_00688_),
    .A2(\samples_real[0][4] ),
    .ZN(_00689_));
 NAND2_X1 _17030_ (.A1(_00686_),
    .A2(net315),
    .ZN(_00690_));
 AOI21_X1 _17031_ (.A(_00672_),
    .B1(_00689_),
    .B2(_00690_),
    .ZN(_00261_));
 NAND2_X1 _17032_ (.A1(_00688_),
    .A2(\samples_real[3][2] ),
    .ZN(_00691_));
 NAND2_X1 _17033_ (.A1(_00686_),
    .A2(net316),
    .ZN(_00692_));
 AOI21_X1 _17034_ (.A(_00672_),
    .B1(_00691_),
    .B2(_00692_),
    .ZN(_00262_));
 NAND2_X1 _17035_ (.A1(_00688_),
    .A2(\samples_real[3][3] ),
    .ZN(_00693_));
 NAND2_X1 _17036_ (.A1(_00686_),
    .A2(net317),
    .ZN(_00694_));
 AOI21_X1 _17037_ (.A(_00672_),
    .B1(_00693_),
    .B2(_00694_),
    .ZN(_00263_));
 CLKBUF_X3 _17038_ (.A(_06735_),
    .Z(_00695_));
 NAND2_X1 _17039_ (.A1(_00688_),
    .A2(\samples_real[3][4] ),
    .ZN(_00696_));
 NAND2_X1 _17040_ (.A1(_00686_),
    .A2(net318),
    .ZN(_00697_));
 AOI21_X1 _17041_ (.A(_00695_),
    .B1(_00696_),
    .B2(_00697_),
    .ZN(_00264_));
 NAND2_X1 _17042_ (.A1(_00688_),
    .A2(\samples_real[3][5] ),
    .ZN(_00698_));
 NAND2_X1 _17043_ (.A1(_00686_),
    .A2(net319),
    .ZN(_00699_));
 AOI21_X1 _17044_ (.A(_00695_),
    .B1(_00698_),
    .B2(_00699_),
    .ZN(_00265_));
 NAND2_X1 _17045_ (.A1(_00688_),
    .A2(\samples_real[3][6] ),
    .ZN(_00700_));
 NAND2_X1 _17046_ (.A1(_00686_),
    .A2(net320),
    .ZN(_00701_));
 AOI21_X1 _17047_ (.A(_00695_),
    .B1(_00700_),
    .B2(_00701_),
    .ZN(_00266_));
 NAND2_X1 _17048_ (.A1(_00688_),
    .A2(\samples_real[3][7] ),
    .ZN(_00702_));
 NAND2_X1 _17049_ (.A1(_00686_),
    .A2(net321),
    .ZN(_00703_));
 AOI21_X1 _17050_ (.A(_00695_),
    .B1(_00702_),
    .B2(_00703_),
    .ZN(_00267_));
 NAND2_X1 _17051_ (.A1(_00688_),
    .A2(\samples_real[3][8] ),
    .ZN(_00704_));
 NAND2_X1 _17052_ (.A1(_00686_),
    .A2(net322),
    .ZN(_00705_));
 AOI21_X1 _17053_ (.A(_00695_),
    .B1(_00704_),
    .B2(_00705_),
    .ZN(_00268_));
 NAND2_X1 _17054_ (.A1(_00688_),
    .A2(\samples_real[3][9] ),
    .ZN(_00706_));
 NAND2_X1 _17055_ (.A1(_00686_),
    .A2(net323),
    .ZN(_00707_));
 AOI21_X1 _17056_ (.A(_00695_),
    .B1(_00706_),
    .B2(_00707_),
    .ZN(_00269_));
 NAND2_X1 _17057_ (.A1(_00688_),
    .A2(\samples_real[3][10] ),
    .ZN(_00708_));
 CLKBUF_X3 _17058_ (.A(_06750_),
    .Z(_00709_));
 NAND2_X1 _17059_ (.A1(_00709_),
    .A2(net324),
    .ZN(_00710_));
 AOI21_X1 _17060_ (.A(_00695_),
    .B1(_00708_),
    .B2(_00710_),
    .ZN(_00270_));
 BUF_X2 _17061_ (.A(_06753_),
    .Z(_00711_));
 NAND2_X1 _17062_ (.A1(_00711_),
    .A2(\samples_real[3][11] ),
    .ZN(_00712_));
 NAND2_X1 _17063_ (.A1(_00709_),
    .A2(net325),
    .ZN(_00713_));
 AOI21_X1 _17064_ (.A(_00695_),
    .B1(_00712_),
    .B2(_00713_),
    .ZN(_00271_));
 NAND2_X1 _17065_ (.A1(_00711_),
    .A2(\samples_real[0][5] ),
    .ZN(_00714_));
 NAND2_X1 _17066_ (.A1(_00709_),
    .A2(net326),
    .ZN(_00715_));
 AOI21_X1 _17067_ (.A(_00695_),
    .B1(_00714_),
    .B2(_00715_),
    .ZN(_00272_));
 NAND2_X1 _17068_ (.A1(_00711_),
    .A2(\samples_real[3][12] ),
    .ZN(_00716_));
 NAND2_X1 _17069_ (.A1(_00709_),
    .A2(net327),
    .ZN(_00717_));
 AOI21_X1 _17070_ (.A(_00695_),
    .B1(_00716_),
    .B2(_00717_),
    .ZN(_00273_));
 CLKBUF_X3 _17071_ (.A(_06735_),
    .Z(_00718_));
 NAND2_X1 _17072_ (.A1(_00711_),
    .A2(\samples_real[3][13] ),
    .ZN(_00719_));
 NAND2_X1 _17073_ (.A1(_00709_),
    .A2(net328),
    .ZN(_00720_));
 AOI21_X1 _17074_ (.A(_00718_),
    .B1(_00719_),
    .B2(_00720_),
    .ZN(_00274_));
 NAND2_X1 _17075_ (.A1(_00711_),
    .A2(\samples_real[3][14] ),
    .ZN(_00721_));
 NAND2_X1 _17076_ (.A1(_00709_),
    .A2(net329),
    .ZN(_00722_));
 AOI21_X1 _17077_ (.A(_00718_),
    .B1(_00721_),
    .B2(_00722_),
    .ZN(_00275_));
 NAND2_X1 _17078_ (.A1(_00711_),
    .A2(\samples_real[3][15] ),
    .ZN(_00723_));
 NAND2_X1 _17079_ (.A1(_00709_),
    .A2(net330),
    .ZN(_00724_));
 AOI21_X1 _17080_ (.A(_00718_),
    .B1(_00723_),
    .B2(_00724_),
    .ZN(_00276_));
 NAND2_X1 _17081_ (.A1(_00711_),
    .A2(\samples_real[4][0] ),
    .ZN(_00725_));
 NAND2_X1 _17082_ (.A1(_00709_),
    .A2(net331),
    .ZN(_00726_));
 AOI21_X1 _17083_ (.A(_00718_),
    .B1(_00725_),
    .B2(_00726_),
    .ZN(_00277_));
 NAND2_X1 _17084_ (.A1(_00711_),
    .A2(\samples_real[4][1] ),
    .ZN(_00727_));
 NAND2_X1 _17085_ (.A1(_00709_),
    .A2(net332),
    .ZN(_00728_));
 AOI21_X1 _17086_ (.A(_00718_),
    .B1(_00727_),
    .B2(_00728_),
    .ZN(_00278_));
 NAND2_X1 _17087_ (.A1(_00711_),
    .A2(\samples_real[4][2] ),
    .ZN(_00729_));
 NAND2_X1 _17088_ (.A1(_00709_),
    .A2(net333),
    .ZN(_00730_));
 AOI21_X1 _17089_ (.A(_00718_),
    .B1(_00729_),
    .B2(_00730_),
    .ZN(_00279_));
 NAND2_X1 _17090_ (.A1(_00711_),
    .A2(\samples_real[4][3] ),
    .ZN(_00731_));
 CLKBUF_X3 _17091_ (.A(_06750_),
    .Z(_00732_));
 NAND2_X1 _17092_ (.A1(_00732_),
    .A2(net334),
    .ZN(_00733_));
 AOI21_X1 _17093_ (.A(_00718_),
    .B1(_00731_),
    .B2(_00733_),
    .ZN(_00280_));
 BUF_X2 _17094_ (.A(_06753_),
    .Z(_00734_));
 NAND2_X1 _17095_ (.A1(_00734_),
    .A2(\samples_real[4][4] ),
    .ZN(_00735_));
 NAND2_X1 _17096_ (.A1(_00732_),
    .A2(net335),
    .ZN(_00736_));
 AOI21_X1 _17097_ (.A(_00718_),
    .B1(_00735_),
    .B2(_00736_),
    .ZN(_00281_));
 NAND2_X1 _17098_ (.A1(_00734_),
    .A2(\samples_real[4][5] ),
    .ZN(_00737_));
 NAND2_X1 _17099_ (.A1(_00732_),
    .A2(net336),
    .ZN(_00738_));
 AOI21_X1 _17100_ (.A(_00718_),
    .B1(_00737_),
    .B2(_00738_),
    .ZN(_00282_));
 NAND2_X1 _17101_ (.A1(_00734_),
    .A2(\samples_real[0][6] ),
    .ZN(_00739_));
 NAND2_X1 _17102_ (.A1(_00732_),
    .A2(net337),
    .ZN(_00740_));
 AOI21_X1 _17103_ (.A(_00718_),
    .B1(_00739_),
    .B2(_00740_),
    .ZN(_00283_));
 CLKBUF_X3 _17104_ (.A(_00843_),
    .Z(_00741_));
 NAND2_X1 _17105_ (.A1(_00734_),
    .A2(\samples_real[4][6] ),
    .ZN(_00742_));
 NAND2_X1 _17106_ (.A1(_00732_),
    .A2(net338),
    .ZN(_00743_));
 AOI21_X1 _17107_ (.A(_00741_),
    .B1(_00742_),
    .B2(_00743_),
    .ZN(_00284_));
 NAND2_X1 _17108_ (.A1(_00734_),
    .A2(\samples_real[4][7] ),
    .ZN(_00744_));
 NAND2_X1 _17109_ (.A1(_00732_),
    .A2(net339),
    .ZN(_00745_));
 AOI21_X1 _17110_ (.A(_00741_),
    .B1(_00744_),
    .B2(_00745_),
    .ZN(_00285_));
 NAND2_X1 _17111_ (.A1(_00734_),
    .A2(\samples_real[4][8] ),
    .ZN(_00746_));
 NAND2_X1 _17112_ (.A1(_00732_),
    .A2(net340),
    .ZN(_00747_));
 AOI21_X1 _17113_ (.A(_00741_),
    .B1(_00746_),
    .B2(_00747_),
    .ZN(_00286_));
 NAND2_X1 _17114_ (.A1(_00734_),
    .A2(\samples_real[4][9] ),
    .ZN(_00748_));
 NAND2_X1 _17115_ (.A1(_00732_),
    .A2(net341),
    .ZN(_00749_));
 AOI21_X1 _17116_ (.A(_00741_),
    .B1(_00748_),
    .B2(_00749_),
    .ZN(_00287_));
 NAND2_X1 _17117_ (.A1(_00734_),
    .A2(\samples_real[4][10] ),
    .ZN(_00750_));
 NAND2_X1 _17118_ (.A1(_00732_),
    .A2(net342),
    .ZN(_00751_));
 AOI21_X1 _17119_ (.A(_00741_),
    .B1(_00750_),
    .B2(_00751_),
    .ZN(_00288_));
 NAND2_X1 _17120_ (.A1(_00734_),
    .A2(\samples_real[4][11] ),
    .ZN(_00752_));
 NAND2_X1 _17121_ (.A1(_00732_),
    .A2(net343),
    .ZN(_00753_));
 AOI21_X1 _17122_ (.A(_00741_),
    .B1(_00752_),
    .B2(_00753_),
    .ZN(_00289_));
 NAND2_X1 _17123_ (.A1(_00734_),
    .A2(\samples_real[4][12] ),
    .ZN(_00754_));
 CLKBUF_X3 _17124_ (.A(_00858_),
    .Z(_00755_));
 NAND2_X1 _17125_ (.A1(_00755_),
    .A2(net344),
    .ZN(_00756_));
 AOI21_X1 _17126_ (.A(_00741_),
    .B1(_00754_),
    .B2(_00756_),
    .ZN(_00290_));
 CLKBUF_X3 _17127_ (.A(_00857_),
    .Z(_00757_));
 NAND2_X1 _17128_ (.A1(_00757_),
    .A2(\samples_real[4][13] ),
    .ZN(_00758_));
 NAND2_X1 _17129_ (.A1(_00755_),
    .A2(net345),
    .ZN(_00759_));
 AOI21_X1 _17130_ (.A(_00741_),
    .B1(_00758_),
    .B2(_00759_),
    .ZN(_00291_));
 NAND2_X1 _17131_ (.A1(_00757_),
    .A2(\samples_real[4][14] ),
    .ZN(_00760_));
 NAND2_X1 _17132_ (.A1(_00755_),
    .A2(net346),
    .ZN(_00761_));
 AOI21_X1 _17133_ (.A(_00741_),
    .B1(_00760_),
    .B2(_00761_),
    .ZN(_00292_));
 NAND2_X1 _17134_ (.A1(_00757_),
    .A2(\samples_real[4][15] ),
    .ZN(_00762_));
 NAND2_X1 _17135_ (.A1(_00755_),
    .A2(net347),
    .ZN(_00763_));
 AOI21_X1 _17136_ (.A(_00741_),
    .B1(_00762_),
    .B2(_00763_),
    .ZN(_00293_));
 CLKBUF_X3 _17137_ (.A(_00843_),
    .Z(_00764_));
 NAND2_X1 _17138_ (.A1(_00757_),
    .A2(\samples_real[0][7] ),
    .ZN(_00765_));
 NAND2_X1 _17139_ (.A1(_00755_),
    .A2(net348),
    .ZN(_00766_));
 AOI21_X1 _17140_ (.A(_00764_),
    .B1(_00765_),
    .B2(_00766_),
    .ZN(_00294_));
 NAND2_X1 _17141_ (.A1(_00757_),
    .A2(\samples_real[5][0] ),
    .ZN(_00767_));
 NAND2_X1 _17142_ (.A1(_00755_),
    .A2(net349),
    .ZN(_00768_));
 AOI21_X1 _17143_ (.A(_00764_),
    .B1(_00767_),
    .B2(_00768_),
    .ZN(_00295_));
 NAND2_X1 _17144_ (.A1(_00757_),
    .A2(\samples_real[5][1] ),
    .ZN(_00769_));
 NAND2_X1 _17145_ (.A1(_00755_),
    .A2(net350),
    .ZN(_00770_));
 AOI21_X1 _17146_ (.A(_00764_),
    .B1(_00769_),
    .B2(_00770_),
    .ZN(_00296_));
 NAND2_X1 _17147_ (.A1(_00757_),
    .A2(\samples_real[5][2] ),
    .ZN(_00771_));
 NAND2_X1 _17148_ (.A1(_00755_),
    .A2(net351),
    .ZN(_00772_));
 AOI21_X1 _17149_ (.A(_00764_),
    .B1(_00771_),
    .B2(_00772_),
    .ZN(_00297_));
 NAND2_X1 _17150_ (.A1(_00757_),
    .A2(\samples_real[5][3] ),
    .ZN(_00773_));
 NAND2_X1 _17151_ (.A1(_00755_),
    .A2(net352),
    .ZN(_00774_));
 AOI21_X1 _17152_ (.A(_00764_),
    .B1(_00773_),
    .B2(_00774_),
    .ZN(_00298_));
 NAND2_X1 _17153_ (.A1(_00757_),
    .A2(\samples_real[5][4] ),
    .ZN(_00775_));
 NAND2_X1 _17154_ (.A1(_00755_),
    .A2(net353),
    .ZN(_00776_));
 AOI21_X1 _17155_ (.A(_00764_),
    .B1(_00775_),
    .B2(_00776_),
    .ZN(_00299_));
 NAND2_X1 _17156_ (.A1(_00757_),
    .A2(\samples_real[5][5] ),
    .ZN(_00777_));
 CLKBUF_X3 _17157_ (.A(_00858_),
    .Z(_00778_));
 NAND2_X1 _17158_ (.A1(_00778_),
    .A2(net354),
    .ZN(_00779_));
 AOI21_X1 _17159_ (.A(_00764_),
    .B1(_00777_),
    .B2(_00779_),
    .ZN(_00300_));
 CLKBUF_X3 _17160_ (.A(_00857_),
    .Z(_00780_));
 NAND2_X1 _17161_ (.A1(_00780_),
    .A2(\samples_real[5][6] ),
    .ZN(_00781_));
 NAND2_X1 _17162_ (.A1(_00778_),
    .A2(net355),
    .ZN(_00782_));
 AOI21_X1 _17163_ (.A(_00764_),
    .B1(_00781_),
    .B2(_00782_),
    .ZN(_00301_));
 NAND2_X1 _17164_ (.A1(_00780_),
    .A2(\samples_real[5][7] ),
    .ZN(_00783_));
 NAND2_X1 _17165_ (.A1(_00778_),
    .A2(net356),
    .ZN(_00784_));
 AOI21_X1 _17166_ (.A(_00764_),
    .B1(_00783_),
    .B2(_00784_),
    .ZN(_00302_));
 NAND2_X1 _17167_ (.A1(_00780_),
    .A2(\samples_real[5][8] ),
    .ZN(_00785_));
 NAND2_X1 _17168_ (.A1(_00778_),
    .A2(net357),
    .ZN(_00786_));
 AOI21_X1 _17169_ (.A(_00764_),
    .B1(_00785_),
    .B2(_00786_),
    .ZN(_00303_));
 BUF_X4 _17170_ (.A(_00843_),
    .Z(_00787_));
 NAND2_X1 _17171_ (.A1(_00780_),
    .A2(\samples_real[5][9] ),
    .ZN(_00788_));
 NAND2_X1 _17172_ (.A1(_00778_),
    .A2(net358),
    .ZN(_00789_));
 AOI21_X1 _17173_ (.A(_00787_),
    .B1(_00788_),
    .B2(_00789_),
    .ZN(_00304_));
 NAND2_X1 _17174_ (.A1(_00780_),
    .A2(\samples_real[0][8] ),
    .ZN(_00790_));
 NAND2_X1 _17175_ (.A1(_00778_),
    .A2(net359),
    .ZN(_00791_));
 AOI21_X1 _17176_ (.A(_00787_),
    .B1(_00790_),
    .B2(_00791_),
    .ZN(_00305_));
 NAND2_X1 _17177_ (.A1(_00780_),
    .A2(\samples_real[5][10] ),
    .ZN(_00792_));
 NAND2_X1 _17178_ (.A1(_00778_),
    .A2(net360),
    .ZN(_00793_));
 AOI21_X1 _17179_ (.A(_00787_),
    .B1(_00792_),
    .B2(_00793_),
    .ZN(_00306_));
 NAND2_X1 _17180_ (.A1(_00780_),
    .A2(\samples_real[5][11] ),
    .ZN(_00794_));
 NAND2_X1 _17181_ (.A1(_00778_),
    .A2(net361),
    .ZN(_00795_));
 AOI21_X1 _17182_ (.A(_00787_),
    .B1(_00794_),
    .B2(_00795_),
    .ZN(_00307_));
 NAND2_X1 _17183_ (.A1(_00780_),
    .A2(\samples_real[5][12] ),
    .ZN(_00796_));
 NAND2_X1 _17184_ (.A1(_00778_),
    .A2(net362),
    .ZN(_00797_));
 AOI21_X1 _17185_ (.A(_00787_),
    .B1(_00796_),
    .B2(_00797_),
    .ZN(_00308_));
 NAND2_X1 _17186_ (.A1(_00780_),
    .A2(\samples_real[5][13] ),
    .ZN(_00798_));
 NAND2_X1 _17187_ (.A1(_00778_),
    .A2(net363),
    .ZN(_00799_));
 AOI21_X1 _17188_ (.A(_00787_),
    .B1(_00798_),
    .B2(_00799_),
    .ZN(_00309_));
 NAND2_X1 _17189_ (.A1(_00780_),
    .A2(\samples_real[5][14] ),
    .ZN(_00800_));
 NAND2_X1 _17190_ (.A1(_06469_),
    .A2(net364),
    .ZN(_00801_));
 AOI21_X1 _17191_ (.A(_00787_),
    .B1(_00800_),
    .B2(_00801_),
    .ZN(_00310_));
 NAND2_X1 _17192_ (.A1(_06447_),
    .A2(\samples_real[5][15] ),
    .ZN(_00802_));
 NAND2_X1 _17193_ (.A1(_06469_),
    .A2(net365),
    .ZN(_00803_));
 AOI21_X1 _17194_ (.A(_00787_),
    .B1(_00802_),
    .B2(_00803_),
    .ZN(_00311_));
 NAND2_X1 _17195_ (.A1(_06447_),
    .A2(\samples_real[6][0] ),
    .ZN(_00804_));
 NAND2_X1 _17196_ (.A1(_06469_),
    .A2(net366),
    .ZN(_00805_));
 AOI21_X1 _17197_ (.A(_00787_),
    .B1(_00804_),
    .B2(_00805_),
    .ZN(_00312_));
 NAND2_X1 _17198_ (.A1(_06447_),
    .A2(\samples_real[6][1] ),
    .ZN(_00806_));
 NAND2_X1 _17199_ (.A1(_06469_),
    .A2(net367),
    .ZN(_00807_));
 AOI21_X1 _17200_ (.A(_00787_),
    .B1(_00806_),
    .B2(_00807_),
    .ZN(_00313_));
 NAND2_X1 _17201_ (.A1(_06447_),
    .A2(\samples_real[6][2] ),
    .ZN(_00808_));
 NAND2_X1 _17202_ (.A1(_06469_),
    .A2(net368),
    .ZN(_00809_));
 AOI21_X1 _17203_ (.A(_00844_),
    .B1(_00808_),
    .B2(_00809_),
    .ZN(_00314_));
 NAND2_X1 _17204_ (.A1(_06447_),
    .A2(\samples_real[6][3] ),
    .ZN(_00810_));
 NAND2_X1 _17205_ (.A1(_06469_),
    .A2(net369),
    .ZN(_00811_));
 AOI21_X1 _17206_ (.A(_00844_),
    .B1(_00810_),
    .B2(_00811_),
    .ZN(_00315_));
 NAND2_X1 _17207_ (.A1(_06447_),
    .A2(\samples_real[0][9] ),
    .ZN(_00812_));
 NAND2_X1 _17208_ (.A1(_06469_),
    .A2(net370),
    .ZN(_00813_));
 AOI21_X1 _17209_ (.A(_00844_),
    .B1(_00812_),
    .B2(_00813_),
    .ZN(_00316_));
 NAND2_X1 _17210_ (.A1(_00862_),
    .A2(_06437_),
    .ZN(_00814_));
 NOR2_X1 _17211_ (.A1(_05300_),
    .A2(_00814_),
    .ZN(_00815_));
 OAI21_X1 _17212_ (.A(_00815_),
    .B1(_09382_),
    .B2(_04771_),
    .ZN(_00816_));
 NAND2_X1 _17213_ (.A1(net371),
    .A2(_00816_),
    .ZN(_00817_));
 AOI21_X1 _17214_ (.A(_00844_),
    .B1(_00815_),
    .B2(_00020_),
    .ZN(_00818_));
 NAND2_X1 _17215_ (.A1(_00817_),
    .A2(_00818_),
    .ZN(_00317_));
 OAI21_X1 _17216_ (.A(_00856_),
    .B1(_06447_),
    .B2(net372),
    .ZN(_00819_));
 NAND2_X1 _17217_ (.A1(net87),
    .A2(_06469_),
    .ZN(_00820_));
 OAI21_X1 _17218_ (.A(_00820_),
    .B1(net372),
    .B2(net87),
    .ZN(_00821_));
 AOI21_X1 _17219_ (.A(_00819_),
    .B1(_00821_),
    .B2(_00860_),
    .ZN(_00318_));
 AOI21_X1 _17220_ (.A(_00814_),
    .B1(_05352_),
    .B2(_00020_),
    .ZN(_00822_));
 NAND2_X2 _17221_ (.A1(_00852_),
    .A2(_00822_),
    .ZN(_00823_));
 NAND2_X1 _17222_ (.A1(_04770_),
    .A2(_00853_),
    .ZN(_00824_));
 OR3_X1 _17223_ (.A1(\sample_count[0] ),
    .A2(_00823_),
    .A3(_00824_),
    .ZN(_00825_));
 NAND2_X1 _17224_ (.A1(\sample_count[0] ),
    .A2(_00823_),
    .ZN(_00826_));
 AOI21_X1 _17225_ (.A(_00844_),
    .B1(_00825_),
    .B2(_00826_),
    .ZN(_00322_));
 NAND3_X1 _17226_ (.A1(_04770_),
    .A2(_00853_),
    .A3(_09379_),
    .ZN(_00827_));
 NOR2_X1 _17227_ (.A1(_00823_),
    .A2(_00827_),
    .ZN(_00828_));
 AOI21_X1 _17228_ (.A(_00828_),
    .B1(_00823_),
    .B2(\sample_count[1] ),
    .ZN(_00829_));
 NOR2_X1 _17229_ (.A1(_00845_),
    .A2(_00829_),
    .ZN(_00323_));
 NAND2_X1 _17230_ (.A1(_00853_),
    .A2(_09383_),
    .ZN(_00830_));
 MUX2_X1 _17231_ (.A(_00830_),
    .B(_05350_),
    .S(_00823_),
    .Z(_00831_));
 NOR2_X1 _17232_ (.A1(_00845_),
    .A2(_00831_),
    .ZN(_00324_));
 NAND2_X1 _17233_ (.A1(_00851_),
    .A2(_04776_),
    .ZN(_00832_));
 NAND4_X1 _17234_ (.A1(_04798_),
    .A2(_00846_),
    .A3(_06440_),
    .A4(_00832_),
    .ZN(_00833_));
 NAND2_X1 _17235_ (.A1(_06440_),
    .A2(_00832_),
    .ZN(_00834_));
 NAND2_X1 _17236_ (.A1(_00849_),
    .A2(_00834_),
    .ZN(_00835_));
 AOI21_X1 _17237_ (.A(_00844_),
    .B1(_00833_),
    .B2(_00835_),
    .ZN(_00581_));
 NAND2_X1 _17238_ (.A1(_00850_),
    .A2(_00834_),
    .ZN(_00836_));
 NAND2_X1 _17239_ (.A1(_00846_),
    .A2(_09364_),
    .ZN(_00837_));
 OAI21_X1 _17240_ (.A(_00836_),
    .B1(_00837_),
    .B2(_00834_),
    .ZN(_00838_));
 AND2_X1 _17241_ (.A1(_00856_),
    .A2(_00838_),
    .ZN(_00582_));
 NAND2_X1 _17242_ (.A1(_00848_),
    .A2(_00834_),
    .ZN(_00839_));
 OR3_X1 _17243_ (.A1(_04775_),
    .A2(_09343_),
    .A3(_00834_),
    .ZN(_00840_));
 AOI21_X1 _17244_ (.A(_00844_),
    .B1(_00839_),
    .B2(_00840_),
    .ZN(_00583_));
 FA_X1 _17245_ (.A(_07347_),
    .B(_07348_),
    .CI(_07349_),
    .CO(_07350_),
    .S(_07351_));
 FA_X1 _17246_ (.A(\temp_imag[0] ),
    .B(_07348_),
    .CI(_07352_),
    .CO(_07353_),
    .S(_07354_));
 FA_X1 _17247_ (.A(_07355_),
    .B(_07356_),
    .CI(_07357_),
    .CO(_07358_),
    .S(_07359_));
 FA_X1 _17248_ (.A(\temp_real[0] ),
    .B(_07356_),
    .CI(_07360_),
    .CO(_07361_),
    .S(_07362_));
 FA_X1 _17249_ (.A(_07363_),
    .B(_00043_),
    .CI(_07364_),
    .CO(_07365_),
    .S(_07366_));
 FA_X1 _17250_ (.A(_07367_),
    .B(_07368_),
    .CI(_07369_),
    .CO(_07370_),
    .S(_07371_));
 FA_X1 _17251_ (.A(_07372_),
    .B(_07373_),
    .CI(_07374_),
    .CO(_07375_),
    .S(_07376_));
 FA_X1 _17252_ (.A(_07377_),
    .B(_07373_),
    .CI(_07378_),
    .CO(_07379_),
    .S(_07380_));
 FA_X1 _17253_ (.A(_07381_),
    .B(_07383_),
    .CI(_07382_),
    .CO(_07384_),
    .S(_07385_));
 FA_X1 _17254_ (.A(_07386_),
    .B(_07388_),
    .CI(_07387_),
    .CO(_07389_),
    .S(_07390_));
 FA_X1 _17255_ (.A(_07391_),
    .B(_07392_),
    .CI(_07393_),
    .CO(_07394_),
    .S(_07395_));
 FA_X1 _17256_ (.A(_07396_),
    .B(_07397_),
    .CI(_07398_),
    .CO(_07399_),
    .S(_07400_));
 FA_X1 _17257_ (.A(_07392_),
    .B(_07393_),
    .CI(_07401_),
    .CO(_07402_),
    .S(_07403_));
 FA_X1 _17258_ (.A(_07404_),
    .B(_07405_),
    .CI(_07406_),
    .CO(_07407_),
    .S(_07408_));
 FA_X1 _17259_ (.A(_07409_),
    .B(_07410_),
    .CI(_07411_),
    .CO(_07412_),
    .S(_07413_));
 FA_X1 _17260_ (.A(_07414_),
    .B(_07413_),
    .CI(_07415_),
    .CO(_07416_),
    .S(_07417_));
 FA_X1 _17261_ (.A(_07418_),
    .B(_07419_),
    .CI(_07403_),
    .CO(_07420_),
    .S(_07421_));
 FA_X1 _17262_ (.A(_07422_),
    .B(_07423_),
    .CI(_07397_),
    .CO(_07424_),
    .S(_07425_));
 FA_X1 _17263_ (.A(_07426_),
    .B(_07427_),
    .CI(_07428_),
    .CO(_07429_),
    .S(_07430_));
 FA_X1 _17264_ (.A(_07394_),
    .B(_07431_),
    .CI(_07432_),
    .CO(_07433_),
    .S(_07434_));
 FA_X1 _17265_ (.A(_07430_),
    .B(_07436_),
    .CI(_07435_),
    .CO(_07437_),
    .S(_07438_));
 FA_X1 _17266_ (.A(_07439_),
    .B(_07440_),
    .CI(_07417_),
    .CO(_07441_),
    .S(_07442_));
 FA_X1 _17267_ (.A(_07443_),
    .B(_07374_),
    .CI(_07381_),
    .CO(_07415_),
    .S(_07444_));
 FA_X1 _17268_ (.A(_07445_),
    .B(_07446_),
    .CI(_07395_),
    .CO(_07447_),
    .S(_07448_));
 FA_X1 _17269_ (.A(_07382_),
    .B(_07383_),
    .CI(_07449_),
    .CO(_07446_),
    .S(_07450_));
 FA_X1 _17270_ (.A(_07397_),
    .B(_07398_),
    .CI(_07451_),
    .CO(_07452_),
    .S(_07453_));
 FA_X1 _17271_ (.A(_07454_),
    .B(_07448_),
    .CI(_07455_),
    .CO(_07456_),
    .S(_07457_));
 FA_X1 _17272_ (.A(_07434_),
    .B(_07458_),
    .CI(_07459_),
    .CO(_07460_),
    .S(_07461_));
 FA_X1 _17273_ (.A(_07462_),
    .B(_07463_),
    .CI(_07464_),
    .CO(_07458_),
    .S(_07465_));
 FA_X1 _17274_ (.A(_07466_),
    .B(_07467_),
    .CI(_07468_),
    .CO(_07469_),
    .S(_07470_));
 FA_X1 _17275_ (.A(_07471_),
    .B(_07472_),
    .CI(_07473_),
    .CO(_07474_),
    .S(_07475_));
 FA_X1 _17276_ (.A(_07476_),
    .B(_07477_),
    .CI(_07478_),
    .CO(_07479_),
    .S(_07480_));
 FA_X1 _17277_ (.A(_07481_),
    .B(_07475_),
    .CI(_07482_),
    .CO(_07483_),
    .S(_07484_));
 FA_X1 _17278_ (.A(_07472_),
    .B(_07485_),
    .CI(_07473_),
    .CO(_07482_),
    .S(_07486_));
 FA_X1 _17279_ (.A(_07470_),
    .B(_07487_),
    .CI(_07438_),
    .CO(_07488_),
    .S(_07489_));
 FA_X1 _17280_ (.A(_07490_),
    .B(_07491_),
    .CI(_07492_),
    .CO(_07487_),
    .S(_07493_));
 FA_X1 _17281_ (.A(_07494_),
    .B(_07495_),
    .CI(_07496_),
    .CO(_07491_),
    .S(_07497_));
 FA_X1 _17282_ (.A(_07498_),
    .B(_07499_),
    .CI(_07500_),
    .CO(_07501_),
    .S(_07502_));
 FA_X1 _17283_ (.A(_07450_),
    .B(_07503_),
    .CI(_07453_),
    .CO(_07455_),
    .S(_07504_));
 FA_X1 _17284_ (.A(_07409_),
    .B(_07410_),
    .CI(_07383_),
    .CO(_07503_),
    .S(_07505_));
 FA_X1 _17285_ (.A(_07423_),
    .B(_07397_),
    .CI(_07398_),
    .CO(_07506_),
    .S(_07507_));
 FA_X1 _17286_ (.A(_07508_),
    .B(_07504_),
    .CI(_07509_),
    .CO(_07510_),
    .S(_07511_));
 FA_X1 _17287_ (.A(_07465_),
    .B(_07512_),
    .CI(_07513_),
    .CO(_07514_),
    .S(_07515_));
 FA_X1 _17288_ (.A(_07516_),
    .B(_07517_),
    .CI(_07518_),
    .CO(_07512_),
    .S(_07519_));
 FA_X1 _17289_ (.A(_07520_),
    .B(_07521_),
    .CI(_07522_),
    .CO(_07523_),
    .S(_07524_));
 FA_X1 _17290_ (.A(_07480_),
    .B(_07525_),
    .CI(_07526_),
    .CO(_07527_),
    .S(_07528_));
 FA_X1 _17291_ (.A(_07529_),
    .B(_07486_),
    .CI(_07530_),
    .CO(_07531_),
    .S(_07532_));
 FA_X1 _17292_ (.A(_07533_),
    .B(_07485_),
    .CI(_07473_),
    .CO(_07530_),
    .S(_07534_));
 FA_X1 _17293_ (.A(_07523_),
    .B(_07528_),
    .CI(_07535_),
    .CO(_07536_),
    .S(_07537_));
 FA_X1 _17294_ (.A(_07537_),
    .B(_07538_),
    .CI(_07489_),
    .CO(_07539_),
    .S(_07540_));
 FA_X1 _17295_ (.A(_07493_),
    .B(_07541_),
    .CI(_07524_),
    .CO(_07538_),
    .S(_07542_));
 FA_X1 _17296_ (.A(_07543_),
    .B(_07544_),
    .CI(_07511_),
    .CO(_07545_),
    .S(_07546_));
 FA_X1 _17297_ (.A(_07377_),
    .B(_07443_),
    .CI(_07378_),
    .CO(_07547_),
    .S(_07548_));
 FA_X1 _17298_ (.A(_07505_),
    .B(_07549_),
    .CI(_07507_),
    .CO(_07509_),
    .S(_07550_));
 FA_X1 _17299_ (.A(_07374_),
    .B(_07410_),
    .CI(_07381_),
    .CO(_07549_),
    .S(_07551_));
 FA_X1 _17300_ (.A(_07383_),
    .B(_07449_),
    .CI(_07552_),
    .CO(_07553_),
    .S(_07554_));
 FA_X1 _17301_ (.A(_07555_),
    .B(_07550_),
    .CI(_07556_),
    .CO(_07557_),
    .S(_07558_));
 FA_X1 _17302_ (.A(_07559_),
    .B(_07519_),
    .CI(_07560_),
    .CO(_07561_),
    .S(_07562_));
 FA_X1 _17303_ (.A(_07553_),
    .B(_07563_),
    .CI(_07564_),
    .CO(_07560_),
    .S(_07565_));
 FA_X1 _17304_ (.A(_07566_),
    .B(_07567_),
    .CI(_07568_),
    .CO(_07569_),
    .S(_07570_));
 FA_X1 _17305_ (.A(_07571_),
    .B(_07572_),
    .CI(_07573_),
    .CO(_07535_),
    .S(_07574_));
 FA_X1 _17306_ (.A(_07472_),
    .B(_07534_),
    .CI(_07575_),
    .CO(_07576_),
    .S(_07577_));
 FA_X1 _17307_ (.A(_07533_),
    .B(_07485_),
    .CI(_07578_),
    .CO(_07575_),
    .S(_07579_));
 FA_X1 _17308_ (.A(_07569_),
    .B(_07574_),
    .CI(_07580_),
    .CO(_07581_),
    .S(_07582_));
 FA_X1 _17309_ (.A(_07584_),
    .B(_07583_),
    .CI(_07585_),
    .CO(_07586_),
    .S(_07587_));
 FA_X1 _17310_ (.A(_07542_),
    .B(_07589_),
    .CI(_07582_),
    .CO(_07588_),
    .S(_07590_));
 FA_X1 _17311_ (.A(_07591_),
    .B(_07592_),
    .CI(_07570_),
    .CO(_07589_),
    .S(_07593_));
 FA_X1 _17312_ (.A(_07594_),
    .B(_07595_),
    .CI(_07558_),
    .CO(_07596_),
    .S(_07597_));
 FA_X1 _17313_ (.A(_07551_),
    .B(_07598_),
    .CI(_07554_),
    .CO(_07556_),
    .S(_07599_));
 FA_X1 _17314_ (.A(_07373_),
    .B(_07381_),
    .CI(_07411_),
    .CO(_07598_),
    .S(_07600_));
 FA_X1 _17315_ (.A(_07410_),
    .B(_07383_),
    .CI(_07449_),
    .CO(_07601_),
    .S(_07602_));
 FA_X1 _17316_ (.A(_07603_),
    .B(_07565_),
    .CI(_07604_),
    .CO(_07605_),
    .S(_07606_));
 FA_X1 _17317_ (.A(_07601_),
    .B(_07607_),
    .CI(_07608_),
    .CO(_07604_),
    .S(_07609_));
 FA_X1 _17318_ (.A(_07610_),
    .B(_07606_),
    .CI(_07611_),
    .CO(_07612_),
    .S(_07613_));
 FA_X1 _17319_ (.A(_07614_),
    .B(_07615_),
    .CI(_07616_),
    .CO(_07580_),
    .S(_07617_));
 FA_X1 _17320_ (.A(_07473_),
    .B(_07579_),
    .CI(_07618_),
    .CO(_07619_),
    .S(_07620_));
 FA_X1 _17321_ (.A(_07621_),
    .B(_07533_),
    .CI(_07578_),
    .CO(_07618_),
    .S(_07622_));
 FA_X1 _17322_ (.A(_07623_),
    .B(_07617_),
    .CI(_07624_),
    .CO(_07625_),
    .S(_07626_));
 FA_X1 _17323_ (.A(_07628_),
    .B(_07627_),
    .CI(_07587_),
    .CO(_07629_),
    .S(_07630_));
 FA_X1 _17324_ (.A(_07631_),
    .B(_07632_),
    .CI(_07633_),
    .CO(_07627_),
    .S(_07634_));
 FA_X1 _17325_ (.A(_07593_),
    .B(_07636_),
    .CI(_07626_),
    .CO(_07635_),
    .S(_07637_));
 FA_X1 _17326_ (.A(_07638_),
    .B(_07639_),
    .CI(_07640_),
    .CO(_07636_),
    .S(_07641_));
 FA_X1 _17327_ (.A(_07642_),
    .B(_07643_),
    .CI(_07644_),
    .CO(_07645_),
    .S(_07646_));
 FA_X1 _17328_ (.A(_07600_),
    .B(_07647_),
    .CI(_07602_),
    .CO(_07648_),
    .S(_07649_));
 FA_X1 _17329_ (.A(_07377_),
    .B(_07443_),
    .CI(_07411_),
    .CO(_07647_),
    .S(_07650_));
 FA_X1 _17330_ (.A(_07410_),
    .B(_07381_),
    .CI(_07383_),
    .CO(_07651_),
    .S(_07652_));
 FA_X1 _17331_ (.A(_07653_),
    .B(_07609_),
    .CI(_07654_),
    .CO(_07611_),
    .S(_07655_));
 FA_X1 _17332_ (.A(_07651_),
    .B(_07656_),
    .CI(_07657_),
    .CO(_07654_),
    .S(_07658_));
 FA_X1 _17333_ (.A(_07659_),
    .B(_07660_),
    .CI(_07661_),
    .CO(_07662_),
    .S(_07663_));
 FA_X1 _17334_ (.A(_07664_),
    .B(_07665_),
    .CI(_07666_),
    .CO(_07624_),
    .S(_07667_));
 FA_X1 _17335_ (.A(_07485_),
    .B(_07622_),
    .CI(_07668_),
    .CO(_07669_),
    .S(_07670_));
 FA_X1 _17336_ (.A(_07671_),
    .B(_07621_),
    .CI(_07578_),
    .CO(_07668_),
    .S(_07672_));
 FA_X1 _17337_ (.A(_07673_),
    .B(_07674_),
    .CI(_07675_),
    .CO(_07676_),
    .S(_07677_));
 FA_X1 _17338_ (.A(_07634_),
    .B(_07678_),
    .CI(_07679_),
    .CO(_07680_),
    .S(_07681_));
 FA_X1 _17339_ (.A(_07682_),
    .B(_07683_),
    .CI(_07684_),
    .CO(_07678_),
    .S(_07685_));
 FA_X1 _17340_ (.A(_07641_),
    .B(_07687_),
    .CI(_07688_),
    .CO(_07686_),
    .S(_07689_));
 FA_X1 _17341_ (.A(_07690_),
    .B(_07691_),
    .CI(_07663_),
    .CO(_07687_),
    .S(_07692_));
 FA_X1 _17342_ (.A(_07693_),
    .B(_07694_),
    .CI(_07695_),
    .CO(_07691_),
    .S(_07696_));
 FA_X1 _17343_ (.A(_07650_),
    .B(_07697_),
    .CI(_07652_),
    .CO(_07698_),
    .S(_07699_));
 FA_X1 _17344_ (.A(_07701_),
    .B(_07702_),
    .CI(_07498_),
    .CO(_07700_),
    .S(_07703_));
 FA_X1 _17345_ (.A(_07410_),
    .B(_07381_),
    .CI(_07411_),
    .CO(_07704_),
    .S(_07705_));
 FA_X1 _17346_ (.A(_07704_),
    .B(_07706_),
    .CI(_07707_),
    .CO(_07708_),
    .S(_07709_));
 FA_X1 _17347_ (.A(_07710_),
    .B(_07711_),
    .CI(_07712_),
    .CO(_07713_),
    .S(_07714_));
 FA_X1 _17348_ (.A(_07533_),
    .B(_07672_),
    .CI(_07715_),
    .CO(_07716_),
    .S(_07717_));
 FA_X1 _17349_ (.A(_07671_),
    .B(_07718_),
    .CI(_07621_),
    .CO(_07715_),
    .S(_07719_));
 FA_X1 _17350_ (.A(_07720_),
    .B(_07721_),
    .CI(_07722_),
    .CO(_07723_),
    .S(_07724_));
 FA_X1 _17351_ (.A(_07685_),
    .B(_07725_),
    .CI(_07726_),
    .CO(_07727_),
    .S(_07728_));
 FA_X1 _17352_ (.A(_07729_),
    .B(_07730_),
    .CI(_07731_),
    .CO(_07725_),
    .S(_07732_));
 FA_X1 _17353_ (.A(_07692_),
    .B(_07734_),
    .CI(_07735_),
    .CO(_07733_),
    .S(_07736_));
 FA_X1 _17354_ (.A(_07737_),
    .B(_07738_),
    .CI(_07739_),
    .CO(_07740_),
    .S(_07741_));
 FA_X1 _17355_ (.A(_07703_),
    .B(_07742_),
    .CI(_07743_),
    .CO(_07744_),
    .S(_07745_));
 FA_X1 _17356_ (.A(_07443_),
    .B(_07381_),
    .CI(_07411_),
    .CO(_07747_),
    .S(_07748_));
 FA_X1 _17357_ (.A(_07747_),
    .B(_07749_),
    .CI(_07750_),
    .CO(_07751_),
    .S(_07752_));
 FA_X1 _17358_ (.A(_07753_),
    .B(_07754_),
    .CI(_07755_),
    .CO(_07756_),
    .S(_07757_));
 FA_X1 _17359_ (.A(_07578_),
    .B(_07719_),
    .CI(_07758_),
    .CO(_07759_),
    .S(_07760_));
 FA_X1 _17360_ (.A(_07559_),
    .B(_07671_),
    .CI(_07718_),
    .CO(_07758_),
    .S(_07761_));
 FA_X1 _17361_ (.A(_07762_),
    .B(_07763_),
    .CI(_07764_),
    .CO(_07765_),
    .S(_07766_));
 FA_X1 _17362_ (.A(_07732_),
    .B(_07767_),
    .CI(_07768_),
    .CO(_07769_),
    .S(_07770_));
 FA_X1 _17363_ (.A(_07771_),
    .B(_07772_),
    .CI(_07773_),
    .CO(_07767_),
    .S(_07774_));
 FA_X1 _17364_ (.A(_07776_),
    .B(_07777_),
    .CI(_07778_),
    .CO(_07775_),
    .S(_07779_));
 FA_X1 _17365_ (.A(_07780_),
    .B(_07781_),
    .CI(_07782_),
    .CO(_07783_),
    .S(_07784_));
 FA_X1 _17366_ (.A(_07702_),
    .B(_07498_),
    .CI(_07500_),
    .CO(_07785_),
    .S(_07786_));
 FA_X1 _17367_ (.A(_07787_),
    .B(_07788_),
    .CI(_07789_),
    .CO(_07790_),
    .S(_07791_));
 FA_X1 _17368_ (.A(_07792_),
    .B(_07793_),
    .CI(_07794_),
    .CO(_07795_),
    .S(_07796_));
 FA_X1 _17369_ (.A(_07621_),
    .B(_07761_),
    .CI(_07797_),
    .CO(_07798_),
    .S(_07799_));
 FA_X1 _17370_ (.A(_07559_),
    .B(_07603_),
    .CI(_07718_),
    .CO(_07797_),
    .S(_07800_));
 FA_X1 _17371_ (.A(_07801_),
    .B(_07802_),
    .CI(_07803_),
    .CO(_07804_),
    .S(_07805_));
 FA_X1 _17372_ (.A(_07774_),
    .B(_07806_),
    .CI(_07807_),
    .CO(_07808_),
    .S(_07809_));
 FA_X1 _17373_ (.A(_07810_),
    .B(_07811_),
    .CI(_07812_),
    .CO(_07806_),
    .S(_07813_));
 FA_X1 _17374_ (.A(_07815_),
    .B(_07816_),
    .CI(_07817_),
    .CO(_07814_),
    .S(_07818_));
 FA_X1 _17375_ (.A(_07819_),
    .B(_07820_),
    .CI(_07821_),
    .CO(_07822_),
    .S(_07823_));
 FA_X1 _17376_ (.A(_07824_),
    .B(_07825_),
    .CI(_07826_),
    .CO(_07827_),
    .S(_07828_));
 FA_X1 _17377_ (.A(_07671_),
    .B(_07800_),
    .CI(_07829_),
    .CO(_07830_),
    .S(_07831_));
 FA_X1 _17378_ (.A(_07559_),
    .B(_07603_),
    .CI(_07653_),
    .CO(_07829_),
    .S(_07832_));
 FA_X1 _17379_ (.A(_07833_),
    .B(_07834_),
    .CI(_07835_),
    .CO(_07836_),
    .S(_07837_));
 FA_X1 _17380_ (.A(_07813_),
    .B(_07838_),
    .CI(_07839_),
    .CO(_07840_),
    .S(_07841_));
 FA_X1 _17381_ (.A(_07842_),
    .B(_07843_),
    .CI(_07844_),
    .CO(_07838_),
    .S(_07845_));
 FA_X1 _17382_ (.A(_07823_),
    .B(_07846_),
    .CI(_07847_),
    .CO(_07843_),
    .S(_07848_));
 FA_X1 _17383_ (.A(_07849_),
    .B(_07850_),
    .CI(_07851_),
    .CO(_07846_),
    .S(_07852_));
 FA_X1 _17384_ (.A(_07702_),
    .B(_07498_),
    .CI(_07853_),
    .CO(_07854_),
    .S(_07855_));
 FA_X1 _17385_ (.A(_07742_),
    .B(_07856_),
    .CI(_07857_),
    .CO(_07858_),
    .S(_07859_));
 FA_X1 _17386_ (.A(_07845_),
    .B(_07860_),
    .CI(_07861_),
    .CO(_07862_),
    .S(_07863_));
 FA_X1 _17387_ (.A(_07848_),
    .B(_07864_),
    .CI(_07865_),
    .CO(_07860_),
    .S(_07866_));
 FA_X1 _17388_ (.A(_07852_),
    .B(_07867_),
    .CI(_07868_),
    .CO(_07864_),
    .S(_07869_));
 FA_X1 _17389_ (.A(_07870_),
    .B(_07871_),
    .CI(_07872_),
    .CO(_07867_),
    .S(_07873_));
 FA_X1 _17390_ (.A(_07718_),
    .B(_07874_),
    .CI(_07832_),
    .CO(_07875_),
    .S(_07876_));
 FA_X1 _17391_ (.A(_07877_),
    .B(_07878_),
    .CI(_07879_),
    .CO(_07880_),
    .S(_07881_));
 FA_X1 _17392_ (.A(_07866_),
    .B(_07882_),
    .CI(_07883_),
    .CO(_07884_),
    .S(_07885_));
 FA_X1 _17393_ (.A(_07869_),
    .B(_07886_),
    .CI(_07887_),
    .CO(_07882_),
    .S(_07888_));
 FA_X1 _17394_ (.A(_07873_),
    .B(_07889_),
    .CI(_07890_),
    .CO(_07886_),
    .S(_07891_));
 FA_X1 _17395_ (.A(_07892_),
    .B(_07893_),
    .CI(_07894_),
    .CO(_07889_),
    .S(_07895_));
 FA_X1 _17396_ (.A(_07896_),
    .B(_07891_),
    .CI(_07897_),
    .CO(_07898_),
    .S(_07899_));
 FA_X1 _17397_ (.A(_07895_),
    .B(_07900_),
    .CI(_07901_),
    .CO(_07897_),
    .S(_07902_));
 FA_X1 _17398_ (.A(_07904_),
    .B(_07905_),
    .CI(_07906_),
    .CO(_07903_),
    .S(_07907_));
 FA_X1 _17399_ (.A(_07907_),
    .B(_07908_),
    .CI(_07909_),
    .CO(_07910_),
    .S(_07911_));
 FA_X1 _17400_ (.A(_07914_),
    .B(_07915_),
    .CI(_07916_),
    .CO(_07917_),
    .S(_07918_));
 FA_X1 _17401_ (.A(_07919_),
    .B(_07920_),
    .CI(_07921_),
    .CO(_07922_),
    .S(_07923_));
 FA_X1 _17402_ (.A(_07918_),
    .B(_07924_),
    .CI(_07925_),
    .CO(_07926_),
    .S(_07927_));
 FA_X1 _17403_ (.A(_07928_),
    .B(_07929_),
    .CI(_07930_),
    .CO(_07931_),
    .S(_07932_));
 FA_X1 _17404_ (.A(_07934_),
    .B(_07935_),
    .CI(_07936_),
    .CO(_07937_),
    .S(_07938_));
 FA_X1 _17405_ (.A(_07939_),
    .B(_07940_),
    .CI(_07941_),
    .CO(_07942_),
    .S(_07943_));
 FA_X1 _17406_ (.A(_07923_),
    .B(_07944_),
    .CI(_07945_),
    .CO(_07946_),
    .S(_07947_));
 FA_X1 _17407_ (.A(_07948_),
    .B(_07949_),
    .CI(_07950_),
    .CO(_07951_),
    .S(_07952_));
 FA_X1 _17408_ (.A(_07953_),
    .B(_07928_),
    .CI(_07929_),
    .CO(_07954_),
    .S(_07955_));
 FA_X1 _17409_ (.A(_07957_),
    .B(_07958_),
    .CI(_07959_),
    .CO(_07960_),
    .S(_07961_));
 FA_X1 _17410_ (.A(_07962_),
    .B(_07963_),
    .CI(_07964_),
    .CO(_07965_),
    .S(_07966_));
 FA_X1 _17411_ (.A(_07940_),
    .B(_07967_),
    .CI(_07968_),
    .CO(_07969_),
    .S(_07970_));
 FA_X1 _17412_ (.A(_07971_),
    .B(_07973_),
    .CI(_07972_),
    .CO(_07974_),
    .S(_07975_));
 FA_X1 _17413_ (.A(_07976_),
    .B(_07978_),
    .CI(_07977_),
    .CO(_07979_),
    .S(_07980_));
 FA_X1 _17414_ (.A(_07969_),
    .B(_07980_),
    .CI(_07981_),
    .CO(_07982_),
    .S(_07983_));
 FA_X1 _17415_ (.A(_07984_),
    .B(_07985_),
    .CI(_07986_),
    .CO(_07987_),
    .S(_07988_));
 FA_X1 _17416_ (.A(_07989_),
    .B(_07990_),
    .CI(_07991_),
    .CO(_07992_),
    .S(_07993_));
 FA_X1 _17417_ (.A(_07994_),
    .B(_07995_),
    .CI(_07996_),
    .CO(_07997_),
    .S(_07998_));
 FA_X1 _17418_ (.A(_07999_),
    .B(_08000_),
    .CI(_08001_),
    .CO(_08002_),
    .S(_08003_));
 FA_X1 _17419_ (.A(_08004_),
    .B(_08005_),
    .CI(_08006_),
    .CO(_08007_),
    .S(_08008_));
 FA_X1 _17420_ (.A(_08009_),
    .B(_07988_),
    .CI(_08010_),
    .CO(_08011_),
    .S(_08012_));
 FA_X1 _17421_ (.A(_08014_),
    .B(_08013_),
    .CI(_07993_),
    .CO(_08015_),
    .S(_08016_));
 FA_X1 _17422_ (.A(_07990_),
    .B(_08017_),
    .CI(_07991_),
    .CO(_08013_),
    .S(_08018_));
 FA_X1 _17423_ (.A(_08019_),
    .B(_08020_),
    .CI(_08021_),
    .CO(_08022_),
    .S(_08023_));
 FA_X1 _17424_ (.A(_08025_),
    .B(_08024_),
    .CI(_08016_),
    .CO(_08026_),
    .S(_08027_));
 FA_X1 _17425_ (.A(_07947_),
    .B(_07975_),
    .CI(_08028_),
    .CO(_08029_),
    .S(_08030_));
 FA_X1 _17426_ (.A(_08031_),
    .B(_08032_),
    .CI(_08033_),
    .CO(_08028_),
    .S(_08034_));
 FA_X1 _17427_ (.A(_08035_),
    .B(_08036_),
    .CI(_08037_),
    .CO(_08038_),
    .S(_08039_));
 FA_X1 _17428_ (.A(_07953_),
    .B(_08040_),
    .CI(_07928_),
    .CO(_08041_),
    .S(_08042_));
 FA_X1 _17429_ (.A(_08044_),
    .B(_08045_),
    .CI(_08046_),
    .CO(_08047_),
    .S(_08048_));
 FA_X1 _17430_ (.A(_08049_),
    .B(_08050_),
    .CI(_08051_),
    .CO(_08052_),
    .S(_08053_));
 FA_X1 _17431_ (.A(_07967_),
    .B(_08054_),
    .CI(_08055_),
    .CO(_08009_),
    .S(_08056_));
 FA_X1 _17432_ (.A(_08057_),
    .B(_08048_),
    .CI(_08058_),
    .CO(_08059_),
    .S(_08060_));
 FA_X1 _17433_ (.A(_08027_),
    .B(_08062_),
    .CI(_08003_),
    .CO(_08063_),
    .S(_08064_));
 FA_X1 _17434_ (.A(_07984_),
    .B(_08065_),
    .CI(_08066_),
    .CO(_08067_),
    .S(_08068_));
 FA_X1 _17435_ (.A(_08069_),
    .B(_08008_),
    .CI(_08070_),
    .CO(_08071_),
    .S(_08072_));
 FA_X1 _17436_ (.A(_08018_),
    .B(_08073_),
    .CI(_08074_),
    .CO(_08024_),
    .S(_08075_));
 FA_X1 _17437_ (.A(_08017_),
    .B(_07977_),
    .CI(_07991_),
    .CO(_08073_),
    .S(_08076_));
 FA_X1 _17438_ (.A(_08077_),
    .B(_08078_),
    .CI(_08079_),
    .CO(_08080_),
    .S(_08081_));
 FA_X1 _17439_ (.A(_08075_),
    .B(_08082_),
    .CI(_08083_),
    .CO(_08084_),
    .S(_08085_));
 FA_X1 _17440_ (.A(_08086_),
    .B(_08087_),
    .CI(_08064_),
    .CO(_08088_),
    .S(_08089_));
 FA_X1 _17441_ (.A(_08091_),
    .B(_08090_),
    .CI(_08030_),
    .CO(_08092_),
    .S(_08093_));
 FA_X1 _17442_ (.A(_08034_),
    .B(_08094_),
    .CI(_08060_),
    .CO(_08090_),
    .S(_08095_));
 FA_X1 _17443_ (.A(_08096_),
    .B(_08097_),
    .CI(_08098_),
    .CO(_08094_),
    .S(_08099_));
 FA_X1 _17444_ (.A(_08100_),
    .B(_08101_),
    .CI(_08102_),
    .CO(_08103_),
    .S(_08104_));
 FA_X1 _17445_ (.A(_08105_),
    .B(_08040_),
    .CI(_07953_),
    .CO(_08106_),
    .S(_08107_));
 FA_X1 _17446_ (.A(_08109_),
    .B(_08110_),
    .CI(_08056_),
    .CO(_08058_),
    .S(_08111_));
 FA_X1 _17447_ (.A(_08112_),
    .B(_08113_),
    .CI(_08114_),
    .CO(_08115_),
    .S(_08116_));
 FA_X1 _17448_ (.A(_08117_),
    .B(_08118_),
    .CI(_08119_),
    .CO(_08120_),
    .S(_08121_));
 FA_X1 _17449_ (.A(_08123_),
    .B(_08124_),
    .CI(_08085_),
    .CO(_08087_),
    .S(_08125_));
 FA_X1 _17450_ (.A(_08126_),
    .B(_08127_),
    .CI(_08004_),
    .CO(_08128_),
    .S(_08129_));
 FA_X1 _17451_ (.A(_08076_),
    .B(_08130_),
    .CI(_08131_),
    .CO(_08082_),
    .S(_08132_));
 FA_X1 _17452_ (.A(_08133_),
    .B(_08017_),
    .CI(_07977_),
    .CO(_08130_),
    .S(_08134_));
 FA_X1 _17453_ (.A(_08135_),
    .B(_08136_),
    .CI(_08137_),
    .CO(_08138_),
    .S(_08139_));
 FA_X1 _17454_ (.A(_08140_),
    .B(_08132_),
    .CI(_08141_),
    .CO(_08142_),
    .S(_08143_));
 FA_X1 _17455_ (.A(_08144_),
    .B(_08145_),
    .CI(_08146_),
    .CO(_08147_),
    .S(_08148_));
 FA_X1 _17456_ (.A(_08150_),
    .B(_08149_),
    .CI(_08151_),
    .CO(_08152_),
    .S(_08153_));
 FA_X1 _17457_ (.A(_08095_),
    .B(_08155_),
    .CI(_08148_),
    .CO(_08154_),
    .S(_08156_));
 FA_X1 _17458_ (.A(_08099_),
    .B(_08157_),
    .CI(_08121_),
    .CO(_08155_),
    .S(_08158_));
 FA_X1 _17459_ (.A(_08159_),
    .B(_08160_),
    .CI(_08161_),
    .CO(_08157_),
    .S(_08162_));
 FA_X1 _17460_ (.A(_08163_),
    .B(_08164_),
    .CI(_08165_),
    .CO(_08166_),
    .S(_08167_));
 FA_X1 _17461_ (.A(_08105_),
    .B(_08168_),
    .CI(_08040_),
    .CO(_08169_),
    .S(_08170_));
 FA_X1 _17462_ (.A(_08171_),
    .B(_08172_),
    .CI(_08173_),
    .CO(_08122_),
    .S(_08174_));
 FA_X1 _17463_ (.A(_08176_),
    .B(_08177_),
    .CI(_08178_),
    .CO(_08175_),
    .S(_08179_));
 FA_X1 _17464_ (.A(_08180_),
    .B(_08181_),
    .CI(_08182_),
    .CO(_08183_),
    .S(_08184_));
 FA_X1 _17465_ (.A(_08186_),
    .B(_08187_),
    .CI(_08143_),
    .CO(_08188_),
    .S(_08189_));
 FA_X1 _17466_ (.A(_08190_),
    .B(_08191_),
    .CI(_08065_),
    .CO(_08192_),
    .S(_08193_));
 FA_X1 _17467_ (.A(_08134_),
    .B(_08194_),
    .CI(_08195_),
    .CO(_08141_),
    .S(_08196_));
 FA_X1 _17468_ (.A(_07941_),
    .B(_08133_),
    .CI(_07977_),
    .CO(_08194_),
    .S(_08197_));
 FA_X1 _17469_ (.A(_08198_),
    .B(_08199_),
    .CI(_08200_),
    .CO(_08201_),
    .S(_08202_));
 FA_X1 _17470_ (.A(_08196_),
    .B(_08203_),
    .CI(_08204_),
    .CO(_08205_),
    .S(_08206_));
 FA_X1 _17471_ (.A(_08207_),
    .B(_08208_),
    .CI(_08209_),
    .CO(_08210_),
    .S(_08211_));
 FA_X1 _17472_ (.A(_08213_),
    .B(_08212_),
    .CI(_08153_),
    .CO(_08214_),
    .S(_08215_));
 FA_X1 _17473_ (.A(_08216_),
    .B(_08217_),
    .CI(_08218_),
    .CO(_08212_),
    .S(_08219_));
 FA_X1 _17474_ (.A(_08158_),
    .B(_08221_),
    .CI(_08211_),
    .CO(_08220_),
    .S(_08222_));
 FA_X1 _17475_ (.A(_08162_),
    .B(_08223_),
    .CI(_08184_),
    .CO(_08221_),
    .S(_08224_));
 FA_X1 _17476_ (.A(_08225_),
    .B(_08226_),
    .CI(_08227_),
    .CO(_08228_),
    .S(_08229_));
 FA_X1 _17477_ (.A(_08168_),
    .B(_08230_),
    .CI(_08105_),
    .CO(_08231_),
    .S(_08232_));
 FA_X1 _17478_ (.A(_08234_),
    .B(_08235_),
    .CI(_08236_),
    .CO(_08185_),
    .S(_08237_));
 FA_X1 _17479_ (.A(_08238_),
    .B(_08239_),
    .CI(_08240_),
    .CO(_08241_),
    .S(_08242_));
 FA_X1 _17480_ (.A(_08243_),
    .B(_08237_),
    .CI(_08244_),
    .CO(_08245_),
    .S(_08246_));
 FA_X1 _17481_ (.A(_08248_),
    .B(_08249_),
    .CI(_08206_),
    .CO(_08250_),
    .S(_08251_));
 FA_X1 _17482_ (.A(_08197_),
    .B(_08252_),
    .CI(_08253_),
    .CO(_08203_),
    .S(_08254_));
 FA_X1 _17483_ (.A(_07941_),
    .B(_07968_),
    .CI(_08133_),
    .CO(_08252_),
    .S(_08255_));
 FA_X1 _17484_ (.A(_08256_),
    .B(_08257_),
    .CI(_08258_),
    .CO(_08259_),
    .S(_08260_));
 FA_X1 _17485_ (.A(_08261_),
    .B(_08262_),
    .CI(_08259_),
    .CO(_08263_),
    .S(_08264_));
 FA_X1 _17486_ (.A(_08245_),
    .B(_08265_),
    .CI(_08266_),
    .CO(_08267_),
    .S(_08268_));
 FA_X1 _17487_ (.A(_08219_),
    .B(_08269_),
    .CI(_08270_),
    .CO(_08271_),
    .S(_08272_));
 FA_X1 _17488_ (.A(_08273_),
    .B(_08274_),
    .CI(_08275_),
    .CO(_08269_),
    .S(_08276_));
 FA_X1 _17489_ (.A(_08224_),
    .B(_08278_),
    .CI(_08279_),
    .CO(_08277_),
    .S(_08280_));
 FA_X1 _17490_ (.A(_08281_),
    .B(_08282_),
    .CI(_08283_),
    .CO(_08278_),
    .S(_08284_));
 FA_X1 _17491_ (.A(_08285_),
    .B(_07921_),
    .CI(_08233_),
    .CO(_08286_),
    .S(_08287_));
 FA_X1 _17492_ (.A(_08288_),
    .B(_08286_),
    .CI(_08289_),
    .CO(_08290_),
    .S(_08291_));
 FA_X1 _17493_ (.A(_08292_),
    .B(_08293_),
    .CI(_08294_),
    .CO(_08295_),
    .S(_08296_));
 FA_X1 _17494_ (.A(_08255_),
    .B(_08298_),
    .CI(_08299_),
    .CO(_08300_),
    .S(_08301_));
 FA_X1 _17495_ (.A(_08055_),
    .B(_07941_),
    .CI(_07968_),
    .CO(_08298_),
    .S(_08302_));
 FA_X1 _17496_ (.A(_08303_),
    .B(_08304_),
    .CI(_08305_),
    .CO(_08306_),
    .S(_08307_));
 FA_X1 _17497_ (.A(_08308_),
    .B(_08309_),
    .CI(_08306_),
    .CO(_08310_),
    .S(_08311_));
 FA_X1 _17498_ (.A(_08295_),
    .B(_08312_),
    .CI(_08313_),
    .CO(_08314_),
    .S(_08315_));
 FA_X1 _17499_ (.A(_08276_),
    .B(_08316_),
    .CI(_08317_),
    .CO(_08318_),
    .S(_08319_));
 FA_X1 _17500_ (.A(_08320_),
    .B(_08321_),
    .CI(_08322_),
    .CO(_08316_),
    .S(_08323_));
 FA_X1 _17501_ (.A(_08284_),
    .B(_08325_),
    .CI(_08326_),
    .CO(_08324_),
    .S(_08327_));
 FA_X1 _17502_ (.A(_08328_),
    .B(_08329_),
    .CI(_08330_),
    .CO(_08325_),
    .S(_08331_));
 FA_X1 _17503_ (.A(_08332_),
    .B(_08333_),
    .CI(_08230_),
    .CO(_08334_),
    .S(_08335_));
 FA_X1 _17504_ (.A(_08337_),
    .B(_08338_),
    .CI(_08339_),
    .CO(_08340_),
    .S(_08341_));
 FA_X1 _17505_ (.A(_08342_),
    .B(_08343_),
    .CI(_08344_),
    .CO(_08345_),
    .S(_08346_));
 FA_X1 _17506_ (.A(_08302_),
    .B(_08348_),
    .CI(_08349_),
    .CO(_08350_),
    .S(_08351_));
 FA_X1 _17507_ (.A(_08352_),
    .B(_08055_),
    .CI(_07968_),
    .CO(_08348_),
    .S(_08353_));
 FA_X1 _17508_ (.A(_08133_),
    .B(_08354_),
    .CI(_08355_),
    .CO(_08356_),
    .S(_08357_));
 FA_X1 _17509_ (.A(_08358_),
    .B(_08359_),
    .CI(_08360_),
    .CO(_08361_),
    .S(_08362_));
 FA_X1 _17510_ (.A(_08345_),
    .B(_08363_),
    .CI(_08364_),
    .CO(_08365_),
    .S(_08366_));
 FA_X1 _17511_ (.A(_08323_),
    .B(_08367_),
    .CI(_08368_),
    .CO(_08369_),
    .S(_08370_));
 FA_X1 _17512_ (.A(_08371_),
    .B(_08372_),
    .CI(_08373_),
    .CO(_08367_),
    .S(_08374_));
 FA_X1 _17513_ (.A(_08331_),
    .B(_08376_),
    .CI(_08377_),
    .CO(_08375_),
    .S(_08378_));
 FA_X1 _17514_ (.A(_08379_),
    .B(_08380_),
    .CI(_08381_),
    .CO(_08376_),
    .S(_08382_));
 FA_X1 _17515_ (.A(_08383_),
    .B(_08384_),
    .CI(_08385_),
    .CO(_08386_),
    .S(_08387_));
 FA_X1 _17516_ (.A(_08353_),
    .B(_08389_),
    .CI(_08390_),
    .CO(_08391_),
    .S(_08392_));
 FA_X1 _17517_ (.A(_08352_),
    .B(_08055_),
    .CI(_08234_),
    .CO(_08389_),
    .S(_08393_));
 FA_X1 _17518_ (.A(_08005_),
    .B(_08394_),
    .CI(_08395_),
    .CO(_08396_),
    .S(_08397_));
 FA_X1 _17519_ (.A(_08398_),
    .B(_08399_),
    .CI(_08396_),
    .CO(_08400_),
    .S(_08401_));
 FA_X1 _17520_ (.A(_08402_),
    .B(_08403_),
    .CI(_08404_),
    .CO(_08405_),
    .S(_08406_));
 FA_X1 _17521_ (.A(_08374_),
    .B(_08408_),
    .CI(_08409_),
    .CO(_08410_),
    .S(_08411_));
 FA_X1 _17522_ (.A(_08412_),
    .B(_08413_),
    .CI(_08414_),
    .CO(_08408_),
    .S(_08415_));
 FA_X1 _17523_ (.A(_08382_),
    .B(_08417_),
    .CI(_08418_),
    .CO(_08416_),
    .S(_08419_));
 FA_X1 _17524_ (.A(_08420_),
    .B(_08421_),
    .CI(_08422_),
    .CO(_08417_),
    .S(_08423_));
 FA_X1 _17525_ (.A(_08333_),
    .B(_08424_),
    .CI(_08332_),
    .CO(_08388_),
    .S(_08425_));
 FA_X1 _17526_ (.A(_08415_),
    .B(_08427_),
    .CI(_08428_),
    .CO(_08429_),
    .S(_08430_));
 FA_X1 _17527_ (.A(_08431_),
    .B(_08432_),
    .CI(_08433_),
    .CO(_08427_),
    .S(_08434_));
 FA_X1 _17528_ (.A(_08435_),
    .B(_08436_),
    .CI(_08437_),
    .CO(_08432_),
    .S(_08438_));
 FA_X1 _17529_ (.A(_08440_),
    .B(_08441_),
    .CI(_08442_),
    .CO(_08439_),
    .S(_08443_));
 FA_X1 _17530_ (.A(_08444_),
    .B(_08445_),
    .CI(_08397_),
    .CO(_08399_),
    .S(_08446_));
 FA_X1 _17531_ (.A(_08066_),
    .B(_08448_),
    .CI(_08449_),
    .CO(_08450_),
    .S(_08451_));
 FA_X1 _17532_ (.A(_08452_),
    .B(_08453_),
    .CI(_08454_),
    .CO(_08455_),
    .S(_08456_));
 FA_X1 _17533_ (.A(_08434_),
    .B(_08457_),
    .CI(_08458_),
    .CO(_08459_),
    .S(_08460_));
 FA_X1 _17534_ (.A(_08438_),
    .B(_08461_),
    .CI(_08462_),
    .CO(_08457_),
    .S(_08463_));
 FA_X1 _17535_ (.A(_08464_),
    .B(_08465_),
    .CI(_08466_),
    .CO(_08461_),
    .S(_08467_));
 FA_X1 _17536_ (.A(_08469_),
    .B(_08470_),
    .CI(_08471_),
    .CO(_08468_),
    .S(_08472_));
 FA_X1 _17537_ (.A(_08473_),
    .B(_08474_),
    .CI(_08475_),
    .CO(_08476_),
    .S(_08477_));
 FA_X1 _17538_ (.A(_08463_),
    .B(_08478_),
    .CI(_08479_),
    .CO(_08480_),
    .S(_08481_));
 FA_X1 _17539_ (.A(_08467_),
    .B(_08482_),
    .CI(_08483_),
    .CO(_08478_),
    .S(_08484_));
 FA_X1 _17540_ (.A(_08485_),
    .B(_08486_),
    .CI(_08487_),
    .CO(_08482_),
    .S(_08488_));
 FA_X1 _17541_ (.A(_08489_),
    .B(_08490_),
    .CI(_08491_),
    .CO(_08486_),
    .S(_08492_));
 FA_X1 _17542_ (.A(_08234_),
    .B(_08493_),
    .CI(_08494_),
    .CO(_08495_),
    .S(_08496_));
 FA_X1 _17543_ (.A(_08497_),
    .B(_08496_),
    .CI(_08498_),
    .CO(_08499_),
    .S(_08500_));
 FA_X1 _17544_ (.A(_08484_),
    .B(_08503_),
    .CI(_08504_),
    .CO(_08505_),
    .S(_08506_));
 FA_X1 _17545_ (.A(_08488_),
    .B(_08507_),
    .CI(_08499_),
    .CO(_08503_),
    .S(_08508_));
 FA_X1 _17546_ (.A(_08510_),
    .B(_08511_),
    .CI(_08512_),
    .CO(_08509_),
    .S(_08513_));
 FA_X1 _17547_ (.A(_08190_),
    .B(_08515_),
    .CI(_08516_),
    .CO(_08502_),
    .S(_08517_));
 FA_X1 _17548_ (.A(_08518_),
    .B(_08517_),
    .CI(_08519_),
    .CO(_08520_),
    .S(_08521_));
 FA_X1 _17549_ (.A(_08055_),
    .B(_08525_),
    .CI(_08526_),
    .CO(_08527_),
    .S(_08528_));
 FA_X1 _17550_ (.A(_08508_),
    .B(_08529_),
    .CI(_08527_),
    .CO(_08530_),
    .S(_08531_));
 FA_X1 _17551_ (.A(_08532_),
    .B(_08533_),
    .CI(_08528_),
    .CO(_08529_),
    .S(_08534_));
 FA_X1 _17552_ (.A(_08536_),
    .B(_08537_),
    .CI(_08538_),
    .CO(_08519_),
    .S(_08539_));
 FA_X1 _17553_ (.A(_08424_),
    .B(_08540_),
    .CI(_08541_),
    .CO(_08542_),
    .S(_08543_));
 FA_X1 _17554_ (.A(_08534_),
    .B(_08544_),
    .CI(_08545_),
    .CO(_08546_),
    .S(_08547_));
 FA_X1 _17555_ (.A(_08548_),
    .B(_08549_),
    .CI(_08550_),
    .CO(_08551_),
    .S(_08552_));
 HA_X1 _17556_ (.A(_08553_),
    .B(_07347_),
    .CO(_08554_),
    .S(_08555_));
 HA_X1 _17557_ (.A(\temp_imag[0] ),
    .B(_08557_),
    .CO(_07352_),
    .S(_08558_));
 HA_X1 _17558_ (.A(\temp_imag[0] ),
    .B(_08559_),
    .CO(_08556_),
    .S(_08560_));
 HA_X1 _17559_ (.A(_08561_),
    .B(_08562_),
    .CO(_08563_),
    .S(_08564_));
 HA_X1 _17560_ (.A(_07347_),
    .B(_08553_),
    .CO(_08565_),
    .S(_08566_));
 HA_X1 _17561_ (.A(\temp_imag[0] ),
    .B(_08553_),
    .CO(_08567_),
    .S(_08568_));
 HA_X1 _17562_ (.A(_07347_),
    .B(_08569_),
    .CO(_08570_),
    .S(_08571_));
 HA_X1 _17563_ (.A(\temp_imag[0] ),
    .B(_08569_),
    .CO(_08572_),
    .S(_08573_));
 HA_X1 _17564_ (.A(_07347_),
    .B(_08574_),
    .CO(_08575_),
    .S(_08576_));
 HA_X1 _17565_ (.A(\temp_imag[0] ),
    .B(_08574_),
    .CO(_08577_),
    .S(_08578_));
 HA_X1 _17566_ (.A(_07347_),
    .B(_08579_),
    .CO(_08580_),
    .S(_08581_));
 HA_X1 _17567_ (.A(\temp_imag[0] ),
    .B(_08579_),
    .CO(_08582_),
    .S(_08583_));
 HA_X1 _17568_ (.A(_07347_),
    .B(_08584_),
    .CO(_08585_),
    .S(_08586_));
 HA_X1 _17569_ (.A(\temp_imag[0] ),
    .B(_08584_),
    .CO(_08587_),
    .S(_08588_));
 HA_X1 _17570_ (.A(_07347_),
    .B(_08589_),
    .CO(_08590_),
    .S(_08591_));
 HA_X1 _17571_ (.A(\temp_imag[0] ),
    .B(_08589_),
    .CO(_08592_),
    .S(_08593_));
 HA_X1 _17572_ (.A(_07347_),
    .B(_08594_),
    .CO(_08595_),
    .S(_08596_));
 HA_X1 _17573_ (.A(\temp_imag[0] ),
    .B(_08594_),
    .CO(_08597_),
    .S(_08598_));
 HA_X1 _17574_ (.A(_07347_),
    .B(_08599_),
    .CO(_08600_),
    .S(_08601_));
 HA_X1 _17575_ (.A(\temp_imag[0] ),
    .B(_08599_),
    .CO(_08602_),
    .S(_08603_));
 HA_X1 _17576_ (.A(_07347_),
    .B(_08604_),
    .CO(_08605_),
    .S(_08606_));
 HA_X1 _17577_ (.A(\temp_imag[0] ),
    .B(_08604_),
    .CO(_08607_),
    .S(_08608_));
 HA_X1 _17578_ (.A(_07347_),
    .B(_08609_),
    .CO(_08610_),
    .S(_08611_));
 HA_X1 _17579_ (.A(\temp_imag[0] ),
    .B(_08609_),
    .CO(_08612_),
    .S(_08613_));
 HA_X1 _17580_ (.A(_07347_),
    .B(_08614_),
    .CO(_08615_),
    .S(_08616_));
 HA_X1 _17581_ (.A(\temp_imag[0] ),
    .B(_08614_),
    .CO(_08617_),
    .S(_08618_));
 HA_X1 _17582_ (.A(_07347_),
    .B(_08619_),
    .CO(_08620_),
    .S(_08621_));
 HA_X1 _17583_ (.A(\temp_imag[0] ),
    .B(net522),
    .CO(_08622_),
    .S(_08623_));
 HA_X1 _17584_ (.A(_07347_),
    .B(_08624_),
    .CO(_08625_),
    .S(_08626_));
 HA_X1 _17585_ (.A(\temp_imag[0] ),
    .B(_08624_),
    .CO(_08627_),
    .S(_08628_));
 HA_X1 _17586_ (.A(_07347_),
    .B(_08629_),
    .CO(_08630_),
    .S(_08631_));
 HA_X1 _17587_ (.A(\temp_imag[0] ),
    .B(net521),
    .CO(_08632_),
    .S(_08633_));
 HA_X1 _17588_ (.A(_08634_),
    .B(_07355_),
    .CO(_08635_),
    .S(_08636_));
 HA_X1 _17589_ (.A(\temp_real[0] ),
    .B(_08638_),
    .CO(_07360_),
    .S(_08639_));
 HA_X1 _17590_ (.A(\temp_real[0] ),
    .B(_08640_),
    .CO(_08637_),
    .S(_08641_));
 HA_X1 _17591_ (.A(_08642_),
    .B(_08643_),
    .CO(_08644_),
    .S(_08645_));
 HA_X1 _17592_ (.A(_07355_),
    .B(_08634_),
    .CO(_08646_),
    .S(_08647_));
 HA_X1 _17593_ (.A(\temp_real[0] ),
    .B(_08634_),
    .CO(_08648_),
    .S(_08649_));
 HA_X1 _17594_ (.A(_07355_),
    .B(_08650_),
    .CO(_08651_),
    .S(_08652_));
 HA_X1 _17595_ (.A(\temp_real[0] ),
    .B(_08650_),
    .CO(_08653_),
    .S(_08654_));
 HA_X1 _17596_ (.A(_07355_),
    .B(_08655_),
    .CO(_08656_),
    .S(_08657_));
 HA_X1 _17597_ (.A(\temp_real[0] ),
    .B(_08655_),
    .CO(_08658_),
    .S(_08659_));
 HA_X1 _17598_ (.A(_07355_),
    .B(_08660_),
    .CO(_08661_),
    .S(_08662_));
 HA_X1 _17599_ (.A(\temp_real[0] ),
    .B(_08660_),
    .CO(_08663_),
    .S(_08664_));
 HA_X1 _17600_ (.A(_07355_),
    .B(_08665_),
    .CO(_08666_),
    .S(_08667_));
 HA_X1 _17601_ (.A(\temp_real[0] ),
    .B(_08665_),
    .CO(_08668_),
    .S(_08669_));
 HA_X1 _17602_ (.A(_07355_),
    .B(_08670_),
    .CO(_08671_),
    .S(_08672_));
 HA_X1 _17603_ (.A(\temp_real[0] ),
    .B(_08670_),
    .CO(_08673_),
    .S(_08674_));
 HA_X1 _17604_ (.A(_07355_),
    .B(_08675_),
    .CO(_08676_),
    .S(_08677_));
 HA_X1 _17605_ (.A(\temp_real[0] ),
    .B(_08675_),
    .CO(_08678_),
    .S(_08679_));
 HA_X1 _17606_ (.A(_07355_),
    .B(_08680_),
    .CO(_08681_),
    .S(_08682_));
 HA_X1 _17607_ (.A(\temp_real[0] ),
    .B(_08680_),
    .CO(_08683_),
    .S(_08684_));
 HA_X1 _17608_ (.A(_07355_),
    .B(_08685_),
    .CO(_08686_),
    .S(_08687_));
 HA_X1 _17609_ (.A(\temp_real[0] ),
    .B(_08685_),
    .CO(_08688_),
    .S(_08689_));
 HA_X1 _17610_ (.A(_07355_),
    .B(_08690_),
    .CO(_08691_),
    .S(_08692_));
 HA_X1 _17611_ (.A(\temp_real[0] ),
    .B(_08690_),
    .CO(_08693_),
    .S(_08694_));
 HA_X1 _17612_ (.A(_07355_),
    .B(_08695_),
    .CO(_08696_),
    .S(_08697_));
 HA_X1 _17613_ (.A(\temp_real[0] ),
    .B(_08695_),
    .CO(_08698_),
    .S(_08699_));
 HA_X1 _17614_ (.A(_07355_),
    .B(_08700_),
    .CO(_08701_),
    .S(_08702_));
 HA_X1 _17615_ (.A(\temp_real[0] ),
    .B(_08700_),
    .CO(_08703_),
    .S(_08704_));
 HA_X1 _17616_ (.A(_07355_),
    .B(_08705_),
    .CO(_08706_),
    .S(_08707_));
 HA_X1 _17617_ (.A(\temp_real[0] ),
    .B(_08705_),
    .CO(_08708_),
    .S(_08709_));
 HA_X1 _17618_ (.A(_07355_),
    .B(_08710_),
    .CO(_08711_),
    .S(_08712_));
 HA_X1 _17619_ (.A(\temp_real[0] ),
    .B(_08710_),
    .CO(_08713_),
    .S(_08714_));
 HA_X1 _17620_ (.A(_08715_),
    .B(net398),
    .CO(_08716_),
    .S(_08717_));
 HA_X1 _17621_ (.A(_07367_),
    .B(_08718_),
    .CO(_08719_),
    .S(_08720_));
 HA_X1 _17622_ (.A(_08721_),
    .B(_08722_),
    .CO(_08723_),
    .S(_08724_));
 HA_X1 _17623_ (.A(_07367_),
    .B(_08725_),
    .CO(_08726_),
    .S(_08727_));
 HA_X1 _17624_ (.A(_08715_),
    .B(net384),
    .CO(_08728_),
    .S(_08729_));
 HA_X1 _17625_ (.A(_08730_),
    .B(_08731_),
    .CO(_08732_),
    .S(_08733_));
 HA_X1 _17626_ (.A(_08721_),
    .B(_08734_),
    .CO(_08735_),
    .S(_08736_));
 HA_X1 _17627_ (.A(_07367_),
    .B(_08737_),
    .CO(_08738_),
    .S(_08739_));
 HA_X1 _17628_ (.A(_08715_),
    .B(_08740_),
    .CO(_08741_),
    .S(_08742_));
 HA_X1 _17629_ (.A(_08743_),
    .B(_08744_),
    .CO(_08745_),
    .S(_08746_));
 HA_X1 _17630_ (.A(_08730_),
    .B(_08747_),
    .CO(_08748_),
    .S(_08749_));
 HA_X1 _17631_ (.A(_08721_),
    .B(_08750_),
    .CO(_08751_),
    .S(_08752_));
 HA_X1 _17632_ (.A(_07367_),
    .B(_08753_),
    .CO(_08754_),
    .S(_08755_));
 HA_X1 _17633_ (.A(_08715_),
    .B(net385),
    .CO(_08756_),
    .S(_08757_));
 HA_X1 _17634_ (.A(_07367_),
    .B(_08758_),
    .CO(_08759_),
    .S(_08760_));
 HA_X1 _17635_ (.A(_08715_),
    .B(_08761_),
    .CO(_08762_),
    .S(_08763_));
 HA_X1 _17636_ (.A(_08764_),
    .B(_08765_),
    .CO(_08766_),
    .S(_08767_));
 HA_X1 _17637_ (.A(_08743_),
    .B(_08768_),
    .CO(_08769_),
    .S(_08770_));
 HA_X1 _17638_ (.A(_08730_),
    .B(_08771_),
    .CO(_08772_),
    .S(_08773_));
 HA_X1 _17639_ (.A(_08721_),
    .B(_08774_),
    .CO(_08775_),
    .S(_08776_));
 HA_X1 _17640_ (.A(_08777_),
    .B(_08778_),
    .CO(_08779_),
    .S(_08780_));
 HA_X1 _17641_ (.A(_08764_),
    .B(_08781_),
    .CO(_08782_),
    .S(_08783_));
 HA_X1 _17642_ (.A(_08743_),
    .B(_08784_),
    .CO(_08785_),
    .S(_08786_));
 HA_X1 _17643_ (.A(_08730_),
    .B(_08787_),
    .CO(_08788_),
    .S(_08789_));
 HA_X1 _17644_ (.A(_08721_),
    .B(_08790_),
    .CO(_08791_),
    .S(_08792_));
 HA_X1 _17645_ (.A(_07367_),
    .B(_08793_),
    .CO(_08794_),
    .S(_08795_));
 HA_X1 _17646_ (.A(_08715_),
    .B(net386),
    .CO(_08796_),
    .S(_08797_));
 HA_X1 _17647_ (.A(_08777_),
    .B(_08798_),
    .CO(_08799_),
    .S(_08800_));
 HA_X1 _17648_ (.A(_08764_),
    .B(_08801_),
    .CO(_08802_),
    .S(_08803_));
 HA_X1 _17649_ (.A(_08743_),
    .B(_08804_),
    .CO(_08805_),
    .S(_08806_));
 HA_X1 _17650_ (.A(_08730_),
    .B(_08807_),
    .CO(_08808_),
    .S(_08809_));
 HA_X1 _17651_ (.A(_08721_),
    .B(_08810_),
    .CO(_08811_),
    .S(_08812_));
 HA_X1 _17652_ (.A(_07367_),
    .B(_08813_),
    .CO(_08814_),
    .S(_08815_));
 HA_X1 _17653_ (.A(_08715_),
    .B(_08816_),
    .CO(_08817_),
    .S(_08818_));
 HA_X1 _17654_ (.A(_08819_),
    .B(_08820_),
    .CO(_08821_),
    .S(_08822_));
 HA_X1 _17655_ (.A(_08777_),
    .B(_08823_),
    .CO(_08824_),
    .S(_08825_));
 HA_X1 _17656_ (.A(_08764_),
    .B(_08826_),
    .CO(_08827_),
    .S(_08828_));
 HA_X1 _17657_ (.A(_08743_),
    .B(_08829_),
    .CO(_08830_),
    .S(_08831_));
 HA_X1 _17658_ (.A(_08721_),
    .B(_08832_),
    .CO(_08833_),
    .S(_08834_));
 HA_X1 _17659_ (.A(_07367_),
    .B(_08835_),
    .CO(_08836_),
    .S(_08837_));
 HA_X1 _17660_ (.A(_08715_),
    .B(net387),
    .CO(_08838_),
    .S(_08839_));
 HA_X1 _17661_ (.A(_08764_),
    .B(_08840_),
    .CO(_08841_),
    .S(_08842_));
 HA_X1 _17662_ (.A(_08743_),
    .B(_08843_),
    .CO(_08844_),
    .S(_08845_));
 HA_X1 _17663_ (.A(_08721_),
    .B(_08846_),
    .CO(_08847_),
    .S(_08848_));
 HA_X1 _17664_ (.A(_08777_),
    .B(_08849_),
    .CO(_08850_),
    .S(_08851_));
 HA_X1 _17665_ (.A(_07367_),
    .B(_08852_),
    .CO(_08853_),
    .S(_08854_));
 HA_X1 _17666_ (.A(_08715_),
    .B(_08855_),
    .CO(_08856_),
    .S(_08857_));
 HA_X1 _17667_ (.A(_08730_),
    .B(_08858_),
    .CO(_08859_),
    .S(_08860_));
 HA_X1 _17668_ (.A(_08721_),
    .B(_08861_),
    .CO(_08862_),
    .S(_08863_));
 HA_X1 _17669_ (.A(_07367_),
    .B(_08864_),
    .CO(_08865_),
    .S(_08866_));
 HA_X1 _17670_ (.A(_08715_),
    .B(net388),
    .CO(_08867_),
    .S(_08868_));
 HA_X1 _17671_ (.A(_08777_),
    .B(_08869_),
    .CO(_08870_),
    .S(_08871_));
 HA_X1 _17672_ (.A(_08764_),
    .B(_08872_),
    .CO(_08873_),
    .S(_08874_));
 HA_X1 _17673_ (.A(_08743_),
    .B(_08875_),
    .CO(_08876_),
    .S(_08877_));
 HA_X1 _17674_ (.A(_08730_),
    .B(_08878_),
    .CO(_08879_),
    .S(_08880_));
 HA_X1 _17675_ (.A(_08730_),
    .B(_08881_),
    .CO(_08882_),
    .S(_08883_));
 HA_X1 _17676_ (.A(_08721_),
    .B(_08884_),
    .CO(_08885_),
    .S(_08886_));
 HA_X1 _17677_ (.A(_07367_),
    .B(_08887_),
    .CO(_08888_),
    .S(_08889_));
 HA_X1 _17678_ (.A(_08715_),
    .B(_08890_),
    .CO(_08891_),
    .S(_08892_));
 HA_X1 _17679_ (.A(_08777_),
    .B(_08893_),
    .CO(_08894_),
    .S(_08895_));
 HA_X1 _17680_ (.A(_08764_),
    .B(_08896_),
    .CO(_08897_),
    .S(_08898_));
 HA_X1 _17681_ (.A(_08743_),
    .B(_08899_),
    .CO(_08900_),
    .S(_08901_));
 HA_X1 _17682_ (.A(_08721_),
    .B(_08902_),
    .CO(_08903_),
    .S(_08904_));
 HA_X1 _17683_ (.A(_07367_),
    .B(_08905_),
    .CO(_08906_),
    .S(_08907_));
 HA_X1 _17684_ (.A(_08743_),
    .B(_08908_),
    .CO(_08909_),
    .S(_08910_));
 HA_X1 _17685_ (.A(_08730_),
    .B(_08911_),
    .CO(_08912_),
    .S(_08913_));
 HA_X1 _17686_ (.A(_08715_),
    .B(net389),
    .CO(_08914_),
    .S(_08915_));
 HA_X1 _17687_ (.A(_08777_),
    .B(_08916_),
    .CO(_08917_),
    .S(_08918_));
 HA_X1 _17688_ (.A(_08764_),
    .B(_08919_),
    .CO(_08920_),
    .S(_08921_));
 HA_X1 _17689_ (.A(_08777_),
    .B(_08922_),
    .CO(_08923_),
    .S(_08924_));
 HA_X1 _17690_ (.A(_08764_),
    .B(_08925_),
    .CO(_08926_),
    .S(_08927_));
 HA_X1 _17691_ (.A(_08743_),
    .B(_08928_),
    .CO(_08929_),
    .S(_08930_));
 HA_X1 _17692_ (.A(_08730_),
    .B(_08931_),
    .CO(_08932_),
    .S(_08933_));
 HA_X1 _17693_ (.A(_08721_),
    .B(_08934_),
    .CO(_08935_),
    .S(_08936_));
 HA_X1 _17694_ (.A(_07367_),
    .B(_08937_),
    .CO(_08938_),
    .S(_08939_));
 HA_X1 _17695_ (.A(_08715_),
    .B(_08940_),
    .CO(_08941_),
    .S(_08942_));
 HA_X1 _17696_ (.A(_08777_),
    .B(_08943_),
    .CO(_08944_),
    .S(_08945_));
 HA_X1 _17697_ (.A(_08764_),
    .B(_08946_),
    .CO(_08947_),
    .S(_08948_));
 HA_X1 _17698_ (.A(_08743_),
    .B(_08949_),
    .CO(_08950_),
    .S(_08951_));
 HA_X1 _17699_ (.A(_08730_),
    .B(_08952_),
    .CO(_08953_),
    .S(_08954_));
 HA_X1 _17700_ (.A(_08721_),
    .B(_08955_),
    .CO(_08956_),
    .S(_08957_));
 HA_X1 _17701_ (.A(_07367_),
    .B(_08958_),
    .CO(_08959_),
    .S(_08960_));
 HA_X1 _17702_ (.A(_08715_),
    .B(net390),
    .CO(_08961_),
    .S(_08962_));
 HA_X1 _17703_ (.A(_08777_),
    .B(_08963_),
    .CO(_08964_),
    .S(_08965_));
 HA_X1 _17704_ (.A(_08764_),
    .B(_08966_),
    .CO(_08967_),
    .S(_08968_));
 HA_X1 _17705_ (.A(_08743_),
    .B(_08969_),
    .CO(_08970_),
    .S(_08971_));
 HA_X1 _17706_ (.A(_08730_),
    .B(_08972_),
    .CO(_08973_),
    .S(_08974_));
 HA_X1 _17707_ (.A(_08721_),
    .B(_08975_),
    .CO(_08976_),
    .S(_08977_));
 HA_X1 _17708_ (.A(_07367_),
    .B(_08978_),
    .CO(_08979_),
    .S(_08980_));
 HA_X1 _17709_ (.A(_08715_),
    .B(_08981_),
    .CO(_08982_),
    .S(_08983_));
 HA_X1 _17710_ (.A(_08715_),
    .B(net391),
    .CO(_08984_),
    .S(_08985_));
 HA_X1 _17711_ (.A(_08721_),
    .B(_08986_),
    .CO(_08987_),
    .S(_08988_));
 HA_X1 _17712_ (.A(_07367_),
    .B(_08989_),
    .CO(_08990_),
    .S(_08991_));
 HA_X1 _17713_ (.A(_08743_),
    .B(_08992_),
    .CO(_08993_),
    .S(_08994_));
 HA_X1 _17714_ (.A(_08730_),
    .B(_08995_),
    .CO(_08996_),
    .S(_08997_));
 HA_X1 _17715_ (.A(_08777_),
    .B(_08998_),
    .CO(_08999_),
    .S(_09000_));
 HA_X1 _17716_ (.A(_08764_),
    .B(_09001_),
    .CO(_09002_),
    .S(_09003_));
 HA_X1 _17717_ (.A(_07367_),
    .B(_09004_),
    .CO(_09005_),
    .S(_09006_));
 HA_X1 _17718_ (.A(net42),
    .B(_09007_),
    .CO(_09008_),
    .S(_09009_));
 HA_X1 _17719_ (.A(_08777_),
    .B(_09010_),
    .CO(_09011_),
    .S(_09012_));
 HA_X1 _17720_ (.A(_08764_),
    .B(_09013_),
    .CO(_09014_),
    .S(_09015_));
 HA_X1 _17721_ (.A(_08743_),
    .B(_09016_),
    .CO(_09017_),
    .S(_09018_));
 HA_X1 _17722_ (.A(_08730_),
    .B(_09019_),
    .CO(_09020_),
    .S(_09021_));
 HA_X1 _17723_ (.A(_08721_),
    .B(_09022_),
    .CO(_09023_),
    .S(_09024_));
 HA_X1 _17724_ (.A(net42),
    .B(net392),
    .CO(_09025_),
    .S(_09026_));
 HA_X1 _17725_ (.A(_08721_),
    .B(_09027_),
    .CO(_09028_),
    .S(_09029_));
 HA_X1 _17726_ (.A(_07367_),
    .B(_09030_),
    .CO(_09031_),
    .S(_09032_));
 HA_X1 _17727_ (.A(_08777_),
    .B(_09033_),
    .CO(_09034_),
    .S(_09035_));
 HA_X1 _17728_ (.A(_08764_),
    .B(_09036_),
    .CO(_09037_),
    .S(_09038_));
 HA_X1 _17729_ (.A(_08743_),
    .B(_09039_),
    .CO(_09040_),
    .S(_09041_));
 HA_X1 _17730_ (.A(_08730_),
    .B(_09042_),
    .CO(_09043_),
    .S(_09044_));
 HA_X1 _17731_ (.A(_08730_),
    .B(_09045_),
    .CO(_09046_),
    .S(_09047_));
 HA_X1 _17732_ (.A(_08721_),
    .B(_09048_),
    .CO(_09049_),
    .S(_09050_));
 HA_X1 _17733_ (.A(_07367_),
    .B(_09051_),
    .CO(_09052_),
    .S(_09053_));
 HA_X1 _17734_ (.A(net42),
    .B(_09054_),
    .CO(_09055_),
    .S(_09056_));
 HA_X1 _17735_ (.A(_08777_),
    .B(_09057_),
    .CO(_09058_),
    .S(_09059_));
 HA_X1 _17736_ (.A(_08764_),
    .B(_09060_),
    .CO(_09061_),
    .S(_09062_));
 HA_X1 _17737_ (.A(_08743_),
    .B(_09063_),
    .CO(_09064_),
    .S(_09065_));
 HA_X1 _17738_ (.A(_08743_),
    .B(_09066_),
    .CO(_09067_),
    .S(_09068_));
 HA_X1 _17739_ (.A(_08730_),
    .B(_09069_),
    .CO(_09070_),
    .S(_09071_));
 HA_X1 _17740_ (.A(_08721_),
    .B(_09072_),
    .CO(_09073_),
    .S(_09074_));
 HA_X1 _17741_ (.A(_09075_),
    .B(_07367_),
    .CO(_09076_),
    .S(_09077_));
 HA_X1 _17742_ (.A(net42),
    .B(net393),
    .CO(_09078_),
    .S(_09079_));
 HA_X1 _17743_ (.A(_08777_),
    .B(_09080_),
    .CO(_09081_),
    .S(_09082_));
 HA_X1 _17744_ (.A(_08764_),
    .B(_09083_),
    .CO(_09084_),
    .S(_09085_));
 HA_X1 _17745_ (.A(_08764_),
    .B(_09086_),
    .CO(_09087_),
    .S(_09088_));
 HA_X1 _17746_ (.A(_08743_),
    .B(_09089_),
    .CO(_09090_),
    .S(_09091_));
 HA_X1 _17747_ (.A(_08730_),
    .B(_09092_),
    .CO(_09093_),
    .S(_09094_));
 HA_X1 _17748_ (.A(_08721_),
    .B(_09095_),
    .CO(_09096_),
    .S(_09097_));
 HA_X1 _17749_ (.A(_09098_),
    .B(_07367_),
    .CO(_09099_),
    .S(_09100_));
 HA_X1 _17750_ (.A(_09101_),
    .B(net42),
    .CO(_09102_),
    .S(_09103_));
 HA_X1 _17751_ (.A(_08777_),
    .B(_09104_),
    .CO(_09105_),
    .S(_09106_));
 HA_X1 _17752_ (.A(_08777_),
    .B(_09107_),
    .CO(_09108_),
    .S(_09109_));
 HA_X1 _17753_ (.A(_08764_),
    .B(_09110_),
    .CO(_09111_),
    .S(_09112_));
 HA_X1 _17754_ (.A(_08743_),
    .B(_09113_),
    .CO(_09114_),
    .S(_09115_));
 HA_X1 _17755_ (.A(_08730_),
    .B(_09116_),
    .CO(_09117_),
    .S(_09118_));
 HA_X1 _17756_ (.A(_08721_),
    .B(_09119_),
    .CO(_09120_),
    .S(_09121_));
 HA_X1 _17757_ (.A(_07367_),
    .B(_09122_),
    .CO(_09123_),
    .S(_09124_));
 HA_X1 _17758_ (.A(net42),
    .B(net394),
    .CO(_09125_),
    .S(_09126_));
 HA_X1 _17759_ (.A(_08777_),
    .B(_09127_),
    .CO(_09128_),
    .S(_09129_));
 HA_X1 _17760_ (.A(_08764_),
    .B(_09130_),
    .CO(_09131_),
    .S(_09132_));
 HA_X1 _17761_ (.A(_08743_),
    .B(_09133_),
    .CO(_09134_),
    .S(_09135_));
 HA_X1 _17762_ (.A(_08730_),
    .B(_09136_),
    .CO(_09137_),
    .S(_09138_));
 HA_X1 _17763_ (.A(_08721_),
    .B(_09139_),
    .CO(_09140_),
    .S(_09141_));
 HA_X1 _17764_ (.A(_07367_),
    .B(_09142_),
    .CO(_09143_),
    .S(_09144_));
 HA_X1 _17765_ (.A(net42),
    .B(_09145_),
    .CO(_09146_),
    .S(_09147_));
 HA_X1 _17766_ (.A(net42),
    .B(net395),
    .CO(_09148_),
    .S(_09149_));
 HA_X1 _17767_ (.A(_08777_),
    .B(_09150_),
    .CO(_09151_),
    .S(_09152_));
 HA_X1 _17768_ (.A(_08764_),
    .B(_09153_),
    .CO(_09154_),
    .S(_09155_));
 HA_X1 _17769_ (.A(_08743_),
    .B(_09156_),
    .CO(_09157_),
    .S(_09158_));
 HA_X1 _17770_ (.A(_08730_),
    .B(_09159_),
    .CO(_09160_),
    .S(_09161_));
 HA_X1 _17771_ (.A(_08721_),
    .B(_09162_),
    .CO(_09163_),
    .S(_09164_));
 HA_X1 _17772_ (.A(_07367_),
    .B(_09165_),
    .CO(_09166_),
    .S(_09167_));
 HA_X1 _17773_ (.A(_07367_),
    .B(_09168_),
    .CO(_09169_),
    .S(_09170_));
 HA_X1 _17774_ (.A(net42),
    .B(_09171_),
    .CO(_09172_),
    .S(_09173_));
 HA_X1 _17775_ (.A(_08764_),
    .B(_09174_),
    .CO(_09175_),
    .S(_09176_));
 HA_X1 _17776_ (.A(_08743_),
    .B(_09177_),
    .CO(_09178_),
    .S(_09179_));
 HA_X1 _17777_ (.A(_08730_),
    .B(_09180_),
    .CO(_09181_),
    .S(_09182_));
 HA_X1 _17778_ (.A(_08721_),
    .B(_09183_),
    .CO(_09184_),
    .S(_09185_));
 HA_X1 _17779_ (.A(_08819_),
    .B(_09186_),
    .CO(_09187_),
    .S(_09188_));
 HA_X1 _17780_ (.A(_08777_),
    .B(_09189_),
    .CO(_09190_),
    .S(_09191_));
 HA_X1 _17781_ (.A(_08721_),
    .B(_09192_),
    .CO(_09193_),
    .S(_09194_));
 HA_X1 _17782_ (.A(_07367_),
    .B(_09195_),
    .CO(_09196_),
    .S(_09197_));
 HA_X1 _17783_ (.A(net42),
    .B(net396),
    .CO(_09198_),
    .S(_09199_));
 HA_X1 _17784_ (.A(_08819_),
    .B(_09200_),
    .CO(_09201_),
    .S(_09202_));
 HA_X1 _17785_ (.A(_08777_),
    .B(_09203_),
    .CO(_09204_),
    .S(_09205_));
 HA_X1 _17786_ (.A(_08764_),
    .B(_09206_),
    .CO(_09207_),
    .S(_09208_));
 HA_X1 _17787_ (.A(_08743_),
    .B(_09209_),
    .CO(_09210_),
    .S(_09211_));
 HA_X1 _17788_ (.A(_08730_),
    .B(_09212_),
    .CO(_09213_),
    .S(_09214_));
 HA_X1 _17789_ (.A(_08730_),
    .B(_09215_),
    .CO(_09216_),
    .S(_09217_));
 HA_X1 _17790_ (.A(_08721_),
    .B(_09218_),
    .CO(_09219_),
    .S(_09220_));
 HA_X1 _17791_ (.A(_07367_),
    .B(_09221_),
    .CO(_09222_),
    .S(_09223_));
 HA_X1 _17792_ (.A(net42),
    .B(_09224_),
    .CO(_09225_),
    .S(_09226_));
 HA_X1 _17793_ (.A(_08819_),
    .B(_09227_),
    .CO(_09228_),
    .S(_09229_));
 HA_X1 _17794_ (.A(_08777_),
    .B(_09230_),
    .CO(_09231_),
    .S(_09232_));
 HA_X1 _17795_ (.A(_08764_),
    .B(_09233_),
    .CO(_09234_),
    .S(_09235_));
 HA_X1 _17796_ (.A(_08743_),
    .B(_09236_),
    .CO(_09237_),
    .S(_09238_));
 HA_X1 _17797_ (.A(net42),
    .B(net397),
    .CO(_09239_),
    .S(_09240_));
 HA_X1 _17798_ (.A(_08721_),
    .B(_09241_),
    .CO(_09242_),
    .S(_09243_));
 HA_X1 _17799_ (.A(_07367_),
    .B(_09244_),
    .CO(_09245_),
    .S(_09246_));
 HA_X1 _17800_ (.A(_08743_),
    .B(_09247_),
    .CO(_09248_),
    .S(_09249_));
 HA_X1 _17801_ (.A(_08730_),
    .B(_09250_),
    .CO(_09251_),
    .S(_09252_));
 HA_X1 _17802_ (.A(_08777_),
    .B(_09253_),
    .CO(_09254_),
    .S(_09255_));
 HA_X1 _17803_ (.A(_08764_),
    .B(_09256_),
    .CO(_09257_),
    .S(_09258_));
 HA_X1 _17804_ (.A(_08819_),
    .B(_09259_),
    .CO(_09260_),
    .S(_09261_));
 HA_X1 _17805_ (.A(_07367_),
    .B(_09262_),
    .CO(_09263_),
    .S(_09264_));
 HA_X1 _17806_ (.A(\butterfly_count[2] ),
    .B(net42),
    .CO(_09265_),
    .S(_09266_));
 HA_X1 _17807_ (.A(_08764_),
    .B(_09267_),
    .CO(_09268_),
    .S(_09269_));
 HA_X1 _17808_ (.A(_08743_),
    .B(_09270_),
    .CO(_09271_),
    .S(_09272_));
 HA_X1 _17809_ (.A(_08730_),
    .B(_09273_),
    .CO(_09274_),
    .S(_09275_));
 HA_X1 _17810_ (.A(_08721_),
    .B(_09276_),
    .CO(_09277_),
    .S(_09278_));
 HA_X1 _17811_ (.A(_08819_),
    .B(_09279_),
    .CO(_09280_),
    .S(_09281_));
 HA_X1 _17812_ (.A(_08777_),
    .B(_09282_),
    .CO(_09283_),
    .S(_09284_));
 HA_X1 _17813_ (.A(_09285_),
    .B(_09286_),
    .CO(_09287_),
    .S(_09288_));
 HA_X1 _17814_ (.A(\butterfly_count[1] ),
    .B(net42),
    .CO(_09289_),
    .S(_09290_));
 HA_X1 _17815_ (.A(_08721_),
    .B(_09291_),
    .CO(_09292_),
    .S(_09293_));
 HA_X1 _17816_ (.A(_07367_),
    .B(_09294_),
    .CO(_09295_),
    .S(_09296_));
 HA_X1 _17817_ (.A(_08777_),
    .B(_09297_),
    .CO(_09298_),
    .S(_09299_));
 HA_X1 _17818_ (.A(_08764_),
    .B(_09300_),
    .CO(_09301_),
    .S(_09302_));
 HA_X1 _17819_ (.A(_08743_),
    .B(_09303_),
    .CO(_09304_),
    .S(_09305_));
 HA_X1 _17820_ (.A(_08730_),
    .B(_09306_),
    .CO(_09307_),
    .S(_09308_));
 HA_X1 _17821_ (.A(_09309_),
    .B(_09310_),
    .CO(_09311_),
    .S(_09312_));
 HA_X1 _17822_ (.A(_09313_),
    .B(_09314_),
    .CO(_09315_),
    .S(_09316_));
 HA_X1 _17823_ (.A(_09318_),
    .B(_09317_),
    .CO(_09319_),
    .S(_09320_));
 HA_X1 _17824_ (.A(_09321_),
    .B(_09322_),
    .CO(_09323_),
    .S(_09324_));
 HA_X1 _17825_ (.A(_09325_),
    .B(_09326_),
    .CO(_09327_),
    .S(_09328_));
 HA_X1 _17826_ (.A(_09329_),
    .B(_09330_),
    .CO(_09331_),
    .S(_09332_));
 HA_X1 _17827_ (.A(_07367_),
    .B(_07368_),
    .CO(_09333_),
    .S(_09334_));
 HA_X1 _17828_ (.A(_09335_),
    .B(_09286_),
    .CO(_09336_),
    .S(_09337_));
 HA_X1 _17829_ (.A(\butterfly_count[0] ),
    .B(net42),
    .CO(_09338_),
    .S(_09339_));
 HA_X1 _17830_ (.A(_09340_),
    .B(_09341_),
    .CO(_09342_),
    .S(_09343_));
 HA_X1 _17831_ (.A(_09340_),
    .B(_09341_),
    .CO(_09325_),
    .S(_09344_));
 HA_X1 _17832_ (.A(\stage[2] ),
    .B(_09341_),
    .CO(_09345_),
    .S(_09346_));
 HA_X1 _17833_ (.A(_09341_),
    .B(\stage[2] ),
    .CO(_09309_),
    .S(_09347_));
 HA_X1 _17834_ (.A(\butterfly_in_group[0] ),
    .B(_09348_),
    .CO(_09349_),
    .S(_00042_));
 HA_X1 _17835_ (.A(\butterfly_in_group[1] ),
    .B(_09350_),
    .CO(_09351_),
    .S(_09352_));
 HA_X1 _17836_ (.A(_09352_),
    .B(_09353_),
    .CO(_09354_),
    .S(_09355_));
 HA_X1 _17837_ (.A(_09355_),
    .B(_09349_),
    .CO(_09356_),
    .S(_00043_));
 HA_X1 _17838_ (.A(_09286_),
    .B(_00042_),
    .CO(_07364_),
    .S(_00044_));
 HA_X1 _17839_ (.A(_09335_),
    .B(_09285_),
    .CO(_09357_),
    .S(_09358_));
 HA_X1 _17840_ (.A(\butterfly_count[0] ),
    .B(\butterfly_count[1] ),
    .CO(_09359_),
    .S(_09360_));
 HA_X1 _17841_ (.A(_09361_),
    .B(_09362_),
    .CO(_09363_),
    .S(_09364_));
 HA_X1 _17842_ (.A(_09361_),
    .B(_09362_),
    .CO(_09365_),
    .S(_09366_));
 HA_X1 _17843_ (.A(_09361_),
    .B(\stage[1] ),
    .CO(_09367_),
    .S(_09368_));
 HA_X1 _17844_ (.A(\stage[0] ),
    .B(_09362_),
    .CO(_09369_),
    .S(_09370_));
 HA_X1 _17845_ (.A(\stage[0] ),
    .B(_09362_),
    .CO(_09371_),
    .S(_09372_));
 HA_X1 _17846_ (.A(\stage[0] ),
    .B(\stage[1] ),
    .CO(_09341_),
    .S(_09373_));
 HA_X1 _17847_ (.A(\stage[0] ),
    .B(\stage[1] ),
    .CO(_09374_),
    .S(_09375_));
 HA_X1 _17848_ (.A(_09376_),
    .B(_09377_),
    .CO(_09378_),
    .S(_09379_));
 HA_X1 _17849_ (.A(\sample_count[0] ),
    .B(\sample_count[1] ),
    .CO(_09380_),
    .S(_09381_));
 HA_X1 _17850_ (.A(\sample_count[2] ),
    .B(_09380_),
    .CO(_09382_),
    .S(_09383_));
 HA_X1 _17851_ (.A(_09384_),
    .B(_09385_),
    .CO(_09386_),
    .S(_09387_));
 HA_X1 _17852_ (.A(_09388_),
    .B(_09387_),
    .CO(_09389_),
    .S(_07404_));
 HA_X1 _17853_ (.A(_09390_),
    .B(_07449_),
    .CO(_09391_),
    .S(_09392_));
 HA_X1 _17854_ (.A(_07380_),
    .B(_07481_),
    .CO(_07405_),
    .S(_07439_));
 HA_X1 _17855_ (.A(_09384_),
    .B(_07377_),
    .CO(_07414_),
    .S(_09393_));
 HA_X1 _17856_ (.A(_09394_),
    .B(_09395_),
    .CO(_09396_),
    .S(_07431_));
 HA_X1 _17857_ (.A(_09397_),
    .B(_09398_),
    .CO(_07432_),
    .S(_07463_));
 HA_X1 _17858_ (.A(_07603_),
    .B(_07671_),
    .CO(_09399_),
    .S(_07459_));
 HA_X1 _17859_ (.A(_09393_),
    .B(_07529_),
    .CO(_07440_),
    .S(_09400_));
 HA_X1 _17860_ (.A(_07444_),
    .B(_09401_),
    .CO(_07454_),
    .S(_09402_));
 HA_X1 _17861_ (.A(_09404_),
    .B(_09405_),
    .CO(_07464_),
    .S(_07516_));
 HA_X1 _17862_ (.A(_07653_),
    .B(_07718_),
    .CO(_09406_),
    .S(_07513_));
 HA_X1 _17863_ (.A(_07621_),
    .B(_07533_),
    .CO(_09407_),
    .S(_09408_));
 HA_X1 _17864_ (.A(_07485_),
    .B(_07578_),
    .CO(_09409_),
    .S(_09410_));
 HA_X1 _17865_ (.A(_09407_),
    .B(_09410_),
    .CO(_09411_),
    .S(_09412_));
 HA_X1 _17866_ (.A(_07671_),
    .B(_07578_),
    .CO(_09414_),
    .S(_09415_));
 HA_X1 _17867_ (.A(_09408_),
    .B(_09414_),
    .CO(_09413_),
    .S(_09416_));
 HA_X1 _17868_ (.A(_07484_),
    .B(_07531_),
    .CO(_09417_),
    .S(_09418_));
 HA_X1 _17869_ (.A(_09420_),
    .B(_07547_),
    .CO(_07508_),
    .S(_09421_));
 HA_X1 _17870_ (.A(_09384_),
    .B(_07472_),
    .CO(_09403_),
    .S(_09422_));
 HA_X1 _17871_ (.A(_09423_),
    .B(_09424_),
    .CO(_07518_),
    .S(_07563_));
 HA_X1 _17872_ (.A(_09425_),
    .B(_09416_),
    .CO(_09419_),
    .S(_09426_));
 HA_X1 _17873_ (.A(_07718_),
    .B(_07621_),
    .CO(_09427_),
    .S(_09428_));
 HA_X1 _17874_ (.A(_09427_),
    .B(_09415_),
    .CO(_09425_),
    .S(_09429_));
 HA_X1 _17875_ (.A(_07532_),
    .B(_07576_),
    .CO(_09430_),
    .S(_09431_));
 HA_X1 _17876_ (.A(_09421_),
    .B(_09422_),
    .CO(_07544_),
    .S(_07594_));
 HA_X1 _17877_ (.A(_07548_),
    .B(_09433_),
    .CO(_07555_),
    .S(_09434_));
 HA_X1 _17878_ (.A(_09435_),
    .B(_09436_),
    .CO(_07564_),
    .S(_07607_));
 HA_X1 _17879_ (.A(_09437_),
    .B(_09429_),
    .CO(_09432_),
    .S(_09438_));
 HA_X1 _17880_ (.A(_07559_),
    .B(_07671_),
    .CO(_09439_),
    .S(_09440_));
 HA_X1 _17881_ (.A(_09439_),
    .B(_09428_),
    .CO(_09437_),
    .S(_09441_));
 HA_X1 _17882_ (.A(_07577_),
    .B(_07619_),
    .CO(_09442_),
    .S(_09443_));
 HA_X1 _17883_ (.A(_09445_),
    .B(_09430_),
    .CO(_09446_),
    .S(_07585_));
 HA_X1 _17884_ (.A(_07473_),
    .B(_09434_),
    .CO(_07595_),
    .S(_07642_));
 HA_X1 _17885_ (.A(_09384_),
    .B(_07372_),
    .CO(_09433_),
    .S(_09447_));
 HA_X1 _17886_ (.A(_07599_),
    .B(_07648_),
    .CO(_07610_),
    .S(_07644_));
 HA_X1 _17887_ (.A(_09448_),
    .B(_09449_),
    .CO(_07608_),
    .S(_07656_));
 HA_X1 _17888_ (.A(_09450_),
    .B(_09441_),
    .CO(_09444_),
    .S(_09451_));
 HA_X1 _17889_ (.A(_07603_),
    .B(_07718_),
    .CO(_09452_),
    .S(_09453_));
 HA_X1 _17890_ (.A(_09452_),
    .B(_09440_),
    .CO(_09450_),
    .S(_09454_));
 HA_X1 _17891_ (.A(_07620_),
    .B(_07669_),
    .CO(_09455_),
    .S(_09456_));
 HA_X1 _17892_ (.A(_09458_),
    .B(_09442_),
    .CO(_07628_),
    .S(_07633_));
 HA_X1 _17893_ (.A(_07485_),
    .B(_09447_),
    .CO(_07643_),
    .S(_09459_));
 HA_X1 _17894_ (.A(_07649_),
    .B(_07698_),
    .CO(_09460_),
    .S(_09461_));
 HA_X1 _17895_ (.A(_09463_),
    .B(_09464_),
    .CO(_07657_),
    .S(_07706_));
 HA_X1 _17896_ (.A(_07670_),
    .B(_07716_),
    .CO(_09466_),
    .S(_09467_));
 HA_X1 _17897_ (.A(_09468_),
    .B(_09454_),
    .CO(_09457_),
    .S(_09469_));
 HA_X1 _17898_ (.A(_07676_),
    .B(_09455_),
    .CO(_07679_),
    .S(_07684_));
 HA_X1 _17899_ (.A(_07630_),
    .B(_07680_),
    .CO(_09470_),
    .S(_09471_));
 HA_X1 _17900_ (.A(_07699_),
    .B(_09472_),
    .CO(_09473_),
    .S(_09474_));
 HA_X1 _17901_ (.A(_07378_),
    .B(_07533_),
    .CO(_09462_),
    .S(_09475_));
 HA_X1 _17902_ (.A(_07658_),
    .B(_07708_),
    .CO(_09465_),
    .S(_09476_));
 HA_X1 _17903_ (.A(_09477_),
    .B(_09478_),
    .CO(_07707_),
    .S(_07749_));
 HA_X1 _17904_ (.A(_09467_),
    .B(_09469_),
    .CO(_07675_),
    .S(_07721_));
 HA_X1 _17905_ (.A(_07717_),
    .B(_07759_),
    .CO(_09480_),
    .S(_09481_));
 HA_X1 _17906_ (.A(_09482_),
    .B(_09453_),
    .CO(_09468_),
    .S(_09483_));
 HA_X1 _17907_ (.A(_07723_),
    .B(_09466_),
    .CO(_07726_),
    .S(_07731_));
 HA_X1 _17908_ (.A(_07681_),
    .B(_07727_),
    .CO(_09484_),
    .S(_09485_));
 HA_X1 _17909_ (.A(_09474_),
    .B(_09475_),
    .CO(_07738_),
    .S(_07780_));
 HA_X1 _17910_ (.A(_07372_),
    .B(_07378_),
    .CO(_07746_),
    .S(_09486_));
 HA_X1 _17911_ (.A(_09487_),
    .B(_09488_),
    .CO(_09489_),
    .S(_09490_));
 HA_X1 _17912_ (.A(_07709_),
    .B(_07751_),
    .CO(_09479_),
    .S(_09491_));
 HA_X1 _17913_ (.A(_09492_),
    .B(_09493_),
    .CO(_07750_),
    .S(_07788_));
 HA_X1 _17914_ (.A(_09481_),
    .B(_09483_),
    .CO(_07722_),
    .S(_07763_));
 HA_X1 _17915_ (.A(_07760_),
    .B(_07798_),
    .CO(_09495_),
    .S(_09496_));
 HA_X1 _17916_ (.A(_07559_),
    .B(_07653_),
    .CO(_09482_),
    .S(_09497_));
 HA_X1 _17917_ (.A(_07765_),
    .B(_09480_),
    .CO(_07768_),
    .S(_07773_));
 HA_X1 _17918_ (.A(_07728_),
    .B(_07769_),
    .CO(_09498_),
    .S(_09499_));
 HA_X1 _17919_ (.A(_07578_),
    .B(_09490_),
    .CO(_07781_),
    .S(_07819_));
 HA_X1 _17920_ (.A(_07748_),
    .B(_09486_),
    .CO(_09488_),
    .S(_09500_));
 HA_X1 _17921_ (.A(_09500_),
    .B(_09501_),
    .CO(_09502_),
    .S(_09503_));
 HA_X1 _17922_ (.A(_07752_),
    .B(_07790_),
    .CO(_09494_),
    .S(_09504_));
 HA_X1 _17923_ (.A(_09505_),
    .B(_09506_),
    .CO(_07789_),
    .S(_07825_));
 HA_X1 _17924_ (.A(_09496_),
    .B(_09497_),
    .CO(_07764_),
    .S(_07802_));
 HA_X1 _17925_ (.A(_07603_),
    .B(_07653_),
    .CO(_07874_),
    .S(_07912_));
 HA_X1 _17926_ (.A(_07799_),
    .B(_07830_),
    .CO(_09508_),
    .S(_09509_));
 HA_X1 _17927_ (.A(_07804_),
    .B(_09495_),
    .CO(_07807_),
    .S(_07812_));
 HA_X1 _17928_ (.A(_07770_),
    .B(_07808_),
    .CO(_09510_),
    .S(_09511_));
 HA_X1 _17929_ (.A(_07621_),
    .B(_09503_),
    .CO(_07820_),
    .S(_07849_));
 HA_X1 _17930_ (.A(_07378_),
    .B(_09512_),
    .CO(_09501_),
    .S(_09513_));
 HA_X1 _17931_ (.A(_07791_),
    .B(_07827_),
    .CO(_09507_),
    .S(_09514_));
 HA_X1 _17932_ (.A(_09515_),
    .B(_09516_),
    .CO(_07826_),
    .S(_09517_));
 HA_X1 _17933_ (.A(_09514_),
    .B(_09518_),
    .CO(_09519_),
    .S(_07851_));
 HA_X1 _17934_ (.A(_07603_),
    .B(_09509_),
    .CO(_07803_),
    .S(_09520_));
 HA_X1 _17935_ (.A(_07559_),
    .B(_07912_),
    .CO(_09521_),
    .S(_09522_));
 HA_X1 _17936_ (.A(_07874_),
    .B(_07832_),
    .CO(_07896_),
    .S(_07901_));
 HA_X1 _17937_ (.A(_07831_),
    .B(_07875_),
    .CO(_09523_),
    .S(_09524_));
 HA_X1 _17938_ (.A(_09526_),
    .B(_09508_),
    .CO(_07839_),
    .S(_07844_));
 HA_X1 _17939_ (.A(_07809_),
    .B(_07840_),
    .CO(_09527_),
    .S(_09528_));
 HA_X1 _17940_ (.A(_07671_),
    .B(_09513_),
    .CO(_07850_),
    .S(_07870_));
 HA_X1 _17941_ (.A(_07828_),
    .B(_09529_),
    .CO(_09518_),
    .S(_09530_));
 HA_X1 _17942_ (.A(_09532_),
    .B(_09533_),
    .CO(_09531_),
    .S(_09534_));
 HA_X1 _17943_ (.A(_09530_),
    .B(_09535_),
    .CO(_09536_),
    .S(_07872_));
 HA_X1 _17944_ (.A(_07653_),
    .B(_09524_),
    .CO(_09525_),
    .S(_09537_));
 HA_X1 _17945_ (.A(_09536_),
    .B(_09537_),
    .CO(_09538_),
    .S(_07868_));
 HA_X1 _17946_ (.A(_09538_),
    .B(_09523_),
    .CO(_07861_),
    .S(_07865_));
 HA_X1 _17947_ (.A(_07841_),
    .B(_07862_),
    .CO(_09539_),
    .S(_09540_));
 HA_X1 _17948_ (.A(_07718_),
    .B(_09541_),
    .CO(_07871_),
    .S(_07892_));
 HA_X1 _17949_ (.A(_09542_),
    .B(_09543_),
    .CO(_09535_),
    .S(_09544_));
 HA_X1 _17950_ (.A(_09545_),
    .B(_09534_),
    .CO(_09543_),
    .S(_09546_));
 HA_X1 _17951_ (.A(_09547_),
    .B(_09548_),
    .CO(_09545_),
    .S(_09549_));
 HA_X1 _17952_ (.A(_09544_),
    .B(_09550_),
    .CO(_09551_),
    .S(_07894_));
 HA_X1 _17953_ (.A(_09521_),
    .B(_07876_),
    .CO(_09552_),
    .S(_09553_));
 HA_X1 _17954_ (.A(_09551_),
    .B(_09553_),
    .CO(_09554_),
    .S(_09555_));
 HA_X1 _17955_ (.A(_09554_),
    .B(_09552_),
    .CO(_07883_),
    .S(_09556_));
 HA_X1 _17956_ (.A(_07863_),
    .B(_07884_),
    .CO(_09557_),
    .S(_09558_));
 HA_X1 _17957_ (.A(_07559_),
    .B(_09486_),
    .CO(_07893_),
    .S(_09559_));
 HA_X1 _17958_ (.A(_09546_),
    .B(_09560_),
    .CO(_09550_),
    .S(_09561_));
 HA_X1 _17959_ (.A(_07885_),
    .B(_09563_),
    .CO(_09564_),
    .S(_09565_));
 HA_X1 _17960_ (.A(_07888_),
    .B(_07898_),
    .CO(_09563_),
    .S(_09566_));
 HA_X1 _17961_ (.A(_09567_),
    .B(_09549_),
    .CO(_09560_),
    .S(_09568_));
 HA_X1 _17962_ (.A(_07378_),
    .B(_07603_),
    .CO(_09562_),
    .S(_09569_));
 HA_X1 _17963_ (.A(_09566_),
    .B(_09570_),
    .CO(_09571_),
    .S(_09572_));
 HA_X1 _17964_ (.A(_07899_),
    .B(_09573_),
    .CO(_09570_),
    .S(_09574_));
 HA_X1 _17965_ (.A(_07902_),
    .B(_09575_),
    .CO(_09573_),
    .S(_09576_));
 HA_X1 _17966_ (.A(_09568_),
    .B(_09569_),
    .CO(_07913_),
    .S(_09577_));
 HA_X1 _17967_ (.A(_09578_),
    .B(_09579_),
    .CO(_09567_),
    .S(_09580_));
 HA_X1 _17968_ (.A(_09577_),
    .B(_09581_),
    .CO(_09582_),
    .S(_09583_));
 HA_X1 _17969_ (.A(_08019_),
    .B(_08336_),
    .CO(_09584_),
    .S(_07919_));
 HA_X1 _17970_ (.A(_07929_),
    .B(_07930_),
    .CO(_09585_),
    .S(_08112_));
 HA_X1 _17971_ (.A(_07914_),
    .B(_07915_),
    .CO(_08051_),
    .S(_09586_));
 HA_X1 _17972_ (.A(_08043_),
    .B(_07933_),
    .CO(_09587_),
    .S(_07924_));
 HA_X1 _17973_ (.A(_08077_),
    .B(_08426_),
    .CO(_07920_),
    .S(_09588_));
 HA_X1 _17974_ (.A(_08108_),
    .B(_07956_),
    .CO(_07925_),
    .S(_07948_));
 HA_X1 _17975_ (.A(_07928_),
    .B(_07929_),
    .CO(_09589_),
    .S(_08176_));
 HA_X1 _17976_ (.A(_07933_),
    .B(_07914_),
    .CO(_08114_),
    .S(_09590_));
 HA_X1 _17977_ (.A(_07927_),
    .B(_07951_),
    .CO(_09591_),
    .S(_07945_));
 HA_X1 _17978_ (.A(_09592_),
    .B(_09593_),
    .CO(_09594_),
    .S(_07934_));
 HA_X1 _17979_ (.A(_07916_),
    .B(_09592_),
    .CO(_07936_),
    .S(_07962_));
 HA_X1 _17980_ (.A(_07953_),
    .B(_07928_),
    .CO(_09595_),
    .S(_08238_));
 HA_X1 _17981_ (.A(_07956_),
    .B(_07933_),
    .CO(_08178_),
    .S(_09596_));
 HA_X1 _17982_ (.A(_08352_),
    .B(_08054_),
    .CO(_08069_),
    .S(_08173_));
 HA_X1 _17983_ (.A(_08173_),
    .B(_07943_),
    .CO(_09597_),
    .S(_07959_));
 HA_X1 _17984_ (.A(_09588_),
    .B(_08233_),
    .CO(_07944_),
    .S(_08031_));
 HA_X1 _17985_ (.A(_07921_),
    .B(_08043_),
    .CO(_07949_),
    .S(_08035_));
 HA_X1 _17986_ (.A(_07952_),
    .B(_08038_),
    .CO(_07971_),
    .S(_08033_));
 HA_X1 _17987_ (.A(_07915_),
    .B(_07916_),
    .CO(_07964_),
    .S(_08049_));
 HA_X1 _17988_ (.A(_07953_),
    .B(_08040_),
    .CO(_09598_),
    .S(_08288_));
 HA_X1 _17989_ (.A(_07956_),
    .B(_08043_),
    .CO(_08240_),
    .S(_09599_));
 HA_X1 _17990_ (.A(_08234_),
    .B(_07970_),
    .CO(_09600_),
    .S(_08046_));
 HA_X1 _17991_ (.A(_08285_),
    .B(_08135_),
    .CO(_08032_),
    .S(_08096_));
 HA_X1 _17992_ (.A(_08108_),
    .B(_08233_),
    .CO(_08036_),
    .S(_08100_));
 HA_X1 _17993_ (.A(_08039_),
    .B(_08103_),
    .CO(_08061_),
    .S(_08098_));
 HA_X1 _17994_ (.A(_08105_),
    .B(_08040_),
    .CO(_09602_),
    .S(_08337_));
 HA_X1 _17995_ (.A(_08108_),
    .B(_08043_),
    .CO(_08289_),
    .S(_09603_));
 HA_X1 _17996_ (.A(_08071_),
    .B(_09604_),
    .CO(_09601_),
    .S(_09605_));
 HA_X1 _17997_ (.A(_08336_),
    .B(_08198_),
    .CO(_08097_),
    .S(_08159_));
 HA_X1 _17998_ (.A(_08285_),
    .B(_07921_),
    .CO(_08101_),
    .S(_08163_));
 HA_X1 _17999_ (.A(_08104_),
    .B(_08166_),
    .CO(_08117_),
    .S(_08161_));
 HA_X1 _18000_ (.A(_08105_),
    .B(_08168_),
    .CO(_09607_),
    .S(_08383_));
 HA_X1 _18001_ (.A(_08108_),
    .B(_07921_),
    .CO(_08339_),
    .S(_09608_));
 HA_X1 _18002_ (.A(_09609_),
    .B(_09610_),
    .CO(_09606_),
    .S(_09611_));
 HA_X1 _18003_ (.A(_09612_),
    .B(_08068_),
    .CO(_09609_),
    .S(_09613_));
 HA_X1 _18004_ (.A(_08147_),
    .B(_08084_),
    .CO(_09615_),
    .S(_08151_));
 HA_X1 _18005_ (.A(_08426_),
    .B(_08256_),
    .CO(_08160_),
    .S(_09616_));
 HA_X1 _18006_ (.A(_08336_),
    .B(_08233_),
    .CO(_08164_),
    .S(_08225_));
 HA_X1 _18007_ (.A(_08167_),
    .B(_08228_),
    .CO(_08180_),
    .S(_09617_));
 HA_X1 _18008_ (.A(_08168_),
    .B(_08230_),
    .CO(_09618_),
    .S(_09619_));
 HA_X1 _18009_ (.A(_07921_),
    .B(_08233_),
    .CO(_08385_),
    .S(_09620_));
 HA_X1 _18010_ (.A(_09621_),
    .B(_09613_),
    .CO(_09614_),
    .S(_09622_));
 HA_X1 _18011_ (.A(_09623_),
    .B(_08129_),
    .CO(_09621_),
    .S(_09624_));
 HA_X1 _18012_ (.A(_08210_),
    .B(_08142_),
    .CO(_08213_),
    .S(_08218_));
 HA_X1 _18013_ (.A(_09616_),
    .B(_09617_),
    .CO(_08223_),
    .S(_08281_));
 HA_X1 _18014_ (.A(_08285_),
    .B(_08426_),
    .CO(_08226_),
    .S(_09626_));
 HA_X1 _18015_ (.A(_08229_),
    .B(_09627_),
    .CO(_08247_),
    .S(_09628_));
 HA_X1 _18016_ (.A(_09629_),
    .B(_09624_),
    .CO(_09625_),
    .S(_09630_));
 HA_X1 _18017_ (.A(_08267_),
    .B(_08205_),
    .CO(_08270_),
    .S(_08275_));
 HA_X1 _18018_ (.A(_08215_),
    .B(_08271_),
    .CO(_09631_),
    .S(_09632_));
 HA_X1 _18019_ (.A(_08303_),
    .B(_09628_),
    .CO(_08282_),
    .S(_08328_));
 HA_X1 _18020_ (.A(_09626_),
    .B(_09633_),
    .CO(_09627_),
    .S(_09634_));
 HA_X1 _18021_ (.A(_09634_),
    .B(_09635_),
    .CO(_08297_),
    .S(_09636_));
 HA_X1 _18022_ (.A(_09637_),
    .B(_09638_),
    .CO(_08244_),
    .S(_08293_));
 HA_X1 _18023_ (.A(_08332_),
    .B(_08333_),
    .CO(_09639_),
    .S(_09640_));
 HA_X1 _18024_ (.A(_08285_),
    .B(_08336_),
    .CO(_09641_),
    .S(_09642_));
 HA_X1 _18025_ (.A(_09643_),
    .B(_09630_),
    .CO(_08266_),
    .S(_08312_));
 HA_X1 _18026_ (.A(_09644_),
    .B(_08193_),
    .CO(_09629_),
    .S(_09645_));
 HA_X1 _18027_ (.A(_08314_),
    .B(_09646_),
    .CO(_08317_),
    .S(_08322_));
 HA_X1 _18028_ (.A(_08272_),
    .B(_08318_),
    .CO(_09647_),
    .S(_09648_));
 HA_X1 _18029_ (.A(_07985_),
    .B(_09636_),
    .CO(_08329_),
    .S(_08379_));
 HA_X1 _18030_ (.A(_08336_),
    .B(_08287_),
    .CO(_09635_),
    .S(_09649_));
 HA_X1 _18031_ (.A(_09649_),
    .B(_09650_),
    .CO(_08347_),
    .S(_09651_));
 HA_X1 _18032_ (.A(_09652_),
    .B(_09653_),
    .CO(_08294_),
    .S(_08343_));
 HA_X1 _18033_ (.A(_08333_),
    .B(_08424_),
    .CO(_09654_),
    .S(_08522_));
 HA_X1 _18034_ (.A(_08336_),
    .B(_08426_),
    .CO(_09655_),
    .S(_09656_));
 HA_X1 _18035_ (.A(_09657_),
    .B(_09645_),
    .CO(_08313_),
    .S(_08363_));
 HA_X1 _18036_ (.A(_08352_),
    .B(_08234_),
    .CO(_08447_),
    .S(_09658_));
 HA_X1 _18037_ (.A(_07967_),
    .B(_08234_),
    .CO(_09644_),
    .S(_09659_));
 HA_X1 _18038_ (.A(_08365_),
    .B(_09660_),
    .CO(_08368_),
    .S(_08373_));
 HA_X1 _18039_ (.A(_08319_),
    .B(_08369_),
    .CO(_09661_),
    .S(_09662_));
 HA_X1 _18040_ (.A(_08005_),
    .B(_09651_),
    .CO(_08380_),
    .S(_08420_));
 HA_X1 _18041_ (.A(_08426_),
    .B(_09663_),
    .CO(_09650_),
    .S(_09664_));
 HA_X1 _18042_ (.A(_09665_),
    .B(_09666_),
    .CO(_08344_),
    .S(_09667_));
 HA_X1 _18043_ (.A(_09668_),
    .B(_09669_),
    .CO(_08407_),
    .S(_08422_));
 HA_X1 _18044_ (.A(_09670_),
    .B(_09659_),
    .CO(_08364_),
    .S(_08403_));
 HA_X1 _18045_ (.A(_08405_),
    .B(_09671_),
    .CO(_08409_),
    .S(_08414_));
 HA_X1 _18046_ (.A(_08370_),
    .B(_08410_),
    .CO(_09672_),
    .S(_09673_));
 HA_X1 _18047_ (.A(_08066_),
    .B(_09664_),
    .CO(_08421_),
    .S(_08440_));
 HA_X1 _18048_ (.A(_09674_),
    .B(_09675_),
    .CO(_09676_),
    .S(_09677_));
 HA_X1 _18049_ (.A(_09619_),
    .B(_08338_),
    .CO(_09678_),
    .S(_09679_));
 HA_X1 _18050_ (.A(_09680_),
    .B(_09681_),
    .CO(_09682_),
    .S(_08442_));
 HA_X1 _18051_ (.A(_08054_),
    .B(_09683_),
    .CO(_08404_),
    .S(_09684_));
 HA_X1 _18052_ (.A(_09685_),
    .B(_09684_),
    .CO(_09686_),
    .S(_08437_));
 HA_X1 _18053_ (.A(_09686_),
    .B(_09687_),
    .CO(_08428_),
    .S(_08433_));
 HA_X1 _18054_ (.A(_08411_),
    .B(_08429_),
    .CO(_09688_),
    .S(_09689_));
 HA_X1 _18055_ (.A(_08127_),
    .B(_09690_),
    .CO(_08441_),
    .S(_08469_));
 HA_X1 _18056_ (.A(_09691_),
    .B(_09692_),
    .CO(_09693_),
    .S(_09694_));
 HA_X1 _18057_ (.A(_09641_),
    .B(_09663_),
    .CO(_09695_),
    .S(_09696_));
 HA_X1 _18058_ (.A(_09697_),
    .B(_09698_),
    .CO(_09699_),
    .S(_08471_));
 HA_X1 _18059_ (.A(_09700_),
    .B(_08456_),
    .CO(_09701_),
    .S(_08466_));
 HA_X1 _18060_ (.A(_09701_),
    .B(_08455_),
    .CO(_08458_),
    .S(_08462_));
 HA_X1 _18061_ (.A(_08430_),
    .B(_08459_),
    .CO(_09702_),
    .S(_09703_));
 HA_X1 _18062_ (.A(_08426_),
    .B(_08190_),
    .CO(_08470_),
    .S(_09704_));
 HA_X1 _18063_ (.A(_09705_),
    .B(_09696_),
    .CO(_09698_),
    .S(_09706_));
 HA_X1 _18064_ (.A(_09640_),
    .B(_09655_),
    .CO(_09705_),
    .S(_09707_));
 HA_X1 _18065_ (.A(_09706_),
    .B(_09707_),
    .CO(_08473_),
    .S(_09708_));
 HA_X1 _18066_ (.A(_09658_),
    .B(_09709_),
    .CO(_08453_),
    .S(_09710_));
 HA_X1 _18067_ (.A(_09710_),
    .B(_08495_),
    .CO(_09711_),
    .S(_09712_));
 HA_X1 _18068_ (.A(_09713_),
    .B(_09712_),
    .CO(_09714_),
    .S(_09715_));
 HA_X1 _18069_ (.A(_09714_),
    .B(_09711_),
    .CO(_08479_),
    .S(_09716_));
 HA_X1 _18070_ (.A(_08460_),
    .B(_08480_),
    .CO(_09717_),
    .S(_09718_));
 HA_X1 _18071_ (.A(_08522_),
    .B(_09719_),
    .CO(_08501_),
    .S(_09720_));
 HA_X1 _18072_ (.A(_08426_),
    .B(_08536_),
    .CO(_09721_),
    .S(_09722_));
 HA_X1 _18073_ (.A(_08496_),
    .B(_08498_),
    .CO(_09723_),
    .S(_09724_));
 HA_X1 _18074_ (.A(_08497_),
    .B(_09724_),
    .CO(_09725_),
    .S(_09726_));
 HA_X1 _18075_ (.A(_09725_),
    .B(_09723_),
    .CO(_08504_),
    .S(_09727_));
 HA_X1 _18076_ (.A(_08481_),
    .B(_08505_),
    .CO(_09728_),
    .S(_09729_));
 HA_X1 _18077_ (.A(_09730_),
    .B(_09731_),
    .CO(_08514_),
    .S(_09732_));
 HA_X1 _18078_ (.A(_08523_),
    .B(_08524_),
    .CO(_08526_),
    .S(_09733_));
 HA_X1 _18079_ (.A(_08522_),
    .B(_09733_),
    .CO(_08525_),
    .S(_09734_));
 HA_X1 _18080_ (.A(_08506_),
    .B(_08530_),
    .CO(_09735_),
    .S(_09736_));
 HA_X1 _18081_ (.A(_09737_),
    .B(_08521_),
    .CO(_08535_),
    .S(_08548_));
 HA_X1 _18082_ (.A(_08540_),
    .B(_08541_),
    .CO(_09738_),
    .S(_09739_));
 HA_X1 _18083_ (.A(_08424_),
    .B(_09739_),
    .CO(_09740_),
    .S(_09741_));
 HA_X1 _18084_ (.A(_09740_),
    .B(_09738_),
    .CO(_08545_),
    .S(_09742_));
 HA_X1 _18085_ (.A(_08531_),
    .B(_08546_),
    .CO(_09744_),
    .S(_09745_));
 HA_X1 _18086_ (.A(_08518_),
    .B(_09746_),
    .CO(_09743_),
    .S(_09747_));
 HA_X1 _18087_ (.A(_09748_),
    .B(_09749_),
    .CO(_08541_),
    .S(_09750_));
 DFF_X1 _18088_ (.D(_00016_),
    .CK(clknet_leaf_36_clk),
    .Q(_00003_),
    .QN(_07340_));
 DFF_X2 _18089_ (.D(_00017_),
    .CK(clknet_leaf_2_clk),
    .Q(_00004_),
    .QN(_07341_));
 DFF_X1 _18090_ (.D(_00018_),
    .CK(clknet_leaf_37_clk),
    .Q(_00005_),
    .QN(_07342_));
 DFF_X1 _18091_ (.D(_00013_),
    .CK(clknet_leaf_74_clk),
    .Q(_00000_),
    .QN(_07343_));
 DFF_X2 _18092_ (.D(_00014_),
    .CK(clknet_leaf_79_clk),
    .Q(_00001_),
    .QN(_07344_));
 DFF_X1 _18093_ (.D(_00015_),
    .CK(clknet_leaf_74_clk),
    .Q(_00002_),
    .QN(_07339_));
 DFF_X1 _18094_ (.D(_00047_),
    .CK(clknet_leaf_66_clk),
    .Q(_00046_),
    .QN(_07345_));
 DFF_X1 _18095_ (.D(_00006_),
    .CK(clknet_leaf_66_clk),
    .Q(_00021_),
    .QN(_00032_));
 DFF_X1 _18096_ (.D(_00048_),
    .CK(clknet_leaf_65_clk),
    .Q(_00022_),
    .QN(_00037_));
 DFF_X1 _18097_ (.D(_00008_),
    .CK(clknet_leaf_67_clk),
    .Q(_00024_),
    .QN(_00033_));
 DFF_X1 _18098_ (.D(_00007_),
    .CK(clknet_leaf_67_clk),
    .Q(_00023_),
    .QN(_00035_));
 DFF_X1 _18099_ (.D(_00049_),
    .CK(clknet_leaf_67_clk),
    .Q(_00025_),
    .QN(_00036_));
 DFF_X1 _18100_ (.D(_00050_),
    .CK(clknet_leaf_67_clk),
    .Q(_00045_),
    .QN(_00034_));
 CLKBUF_X3 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_0_clk));
 LOGIC1_X1 _17620__319 (.Z(net398));
 DFF_X1 \bit_rev_idx[0]$_SDFFE_PN0P_  (.D(_00051_),
    .CK(clknet_leaf_2_clk),
    .Q(\bit_rev_idx[0] ),
    .QN(_00039_));
 DFF_X2 \bit_rev_idx[1]$_SDFFE_PN0P_  (.D(_00052_),
    .CK(clknet_leaf_2_clk),
    .Q(\bit_rev_idx[1] ),
    .QN(_00027_));
 DFF_X1 \bit_rev_idx[2]$_SDFFE_PN0P_  (.D(_00053_),
    .CK(clknet_leaf_2_clk),
    .Q(\bit_rev_idx[2] ),
    .QN(_00029_));
 DFF_X2 \busy$_SDFFE_PN0P_  (.D(_00054_),
    .CK(clknet_leaf_79_clk),
    .Q(net88),
    .QN(_07338_));
 DFF_X2 \butterfly_count[0]$_SDFFE_PN0P_  (.D(_00055_),
    .CK(clknet_leaf_78_clk),
    .Q(\butterfly_count[0] ),
    .QN(_09335_));
 DFF_X2 \butterfly_count[1]$_SDFFE_PN0P_  (.D(_00056_),
    .CK(clknet_leaf_78_clk),
    .Q(\butterfly_count[1] ),
    .QN(_09285_));
 DFF_X1 \butterfly_count[2]$_SDFFE_PN0P_  (.D(_00057_),
    .CK(clknet_leaf_77_clk),
    .Q(\butterfly_count[2] ),
    .QN(_00040_));
 DFF_X1 \butterfly_in_group[0]$_DFFE_PP_  (.D(_00058_),
    .CK(clknet_leaf_77_clk),
    .Q(\butterfly_in_group[0] ),
    .QN(_07337_));
 DFF_X2 \butterfly_in_group[1]$_DFFE_PP_  (.D(_00059_),
    .CK(clknet_leaf_77_clk),
    .Q(\butterfly_in_group[1] ),
    .QN(_07336_));
 DFF_X1 \butterfly_in_group[2]$_DFFE_PP_  (.D(_00060_),
    .CK(clknet_leaf_77_clk),
    .Q(\butterfly_in_group[2] ),
    .QN(_07335_));
 DFF_X1 \data_out_imag[0]$_SDFFE_PN0P_  (.D(_00061_),
    .CK(clknet_3_0__leaf_clk),
    .Q(net89),
    .QN(_07334_));
 DFF_X1 \data_out_imag[100]$_SDFFE_PN0P_  (.D(_00062_),
    .CK(clknet_leaf_0_clk),
    .Q(net90),
    .QN(_07333_));
 DFF_X2 \data_out_imag[101]$_SDFFE_PN0P_  (.D(_00063_),
    .CK(clknet_leaf_0_clk),
    .Q(net91),
    .QN(_07332_));
 DFF_X1 \data_out_imag[102]$_SDFFE_PN0P_  (.D(_00064_),
    .CK(clknet_leaf_81_clk),
    .Q(net92),
    .QN(_07331_));
 DFF_X1 \data_out_imag[103]$_SDFFE_PN0P_  (.D(_00065_),
    .CK(clknet_leaf_82_clk),
    .Q(net95),
    .QN(_07330_));
 DFF_X1 \data_out_imag[104]$_SDFFE_PN0P_  (.D(_00066_),
    .CK(clknet_leaf_0_clk),
    .Q(net96),
    .QN(_07329_));
 DFF_X1 \data_out_imag[105]$_SDFFE_PN0P_  (.D(_00067_),
    .CK(clknet_leaf_0_clk),
    .Q(net99),
    .QN(_07328_));
 DFF_X1 \data_out_imag[106]$_SDFFE_PN0P_  (.D(_00068_),
    .CK(clknet_leaf_81_clk),
    .Q(net100),
    .QN(_07327_));
 DFF_X1 \data_out_imag[107]$_SDFFE_PN0P_  (.D(_00069_),
    .CK(clknet_leaf_81_clk),
    .Q(net102),
    .QN(_07326_));
 DFF_X1 \data_out_imag[108]$_SDFFE_PN0P_  (.D(_00070_),
    .CK(clknet_leaf_80_clk),
    .Q(net103),
    .QN(_07325_));
 DFF_X1 \data_out_imag[109]$_SDFFE_PN0P_  (.D(_00071_),
    .CK(clknet_leaf_81_clk),
    .Q(net105),
    .QN(_07324_));
 DFF_X1 \data_out_imag[10]$_SDFFE_PN0P_  (.D(_00072_),
    .CK(clknet_leaf_0_clk),
    .Q(net106),
    .QN(_07323_));
 DFF_X1 \data_out_imag[110]$_SDFFE_PN0P_  (.D(_00073_),
    .CK(clknet_leaf_80_clk),
    .Q(net108),
    .QN(_07322_));
 DFF_X2 \data_out_imag[111]$_SDFFE_PN0P_  (.D(_00074_),
    .CK(clknet_leaf_1_clk),
    .Q(net109),
    .QN(_07321_));
 DFF_X1 \data_out_imag[112]$_SDFFE_PN0P_  (.D(_00075_),
    .CK(clknet_leaf_80_clk),
    .Q(net110),
    .QN(_07320_));
 DFF_X1 \data_out_imag[113]$_SDFFE_PN0P_  (.D(_00076_),
    .CK(clknet_leaf_81_clk),
    .Q(net111),
    .QN(_07319_));
 DFF_X2 \data_out_imag[114]$_SDFFE_PN0P_  (.D(_00077_),
    .CK(clknet_leaf_1_clk),
    .Q(net112),
    .QN(_07318_));
 DFF_X2 \data_out_imag[115]$_SDFFE_PN0P_  (.D(_00078_),
    .CK(clknet_leaf_1_clk),
    .Q(net113),
    .QN(_07317_));
 DFF_X2 \data_out_imag[116]$_SDFFE_PN0P_  (.D(_00079_),
    .CK(clknet_leaf_0_clk),
    .Q(net114),
    .QN(_07316_));
 DFF_X2 \data_out_imag[117]$_SDFFE_PN0P_  (.D(_00080_),
    .CK(clknet_leaf_0_clk),
    .Q(net115),
    .QN(_07315_));
 DFF_X1 \data_out_imag[118]$_SDFFE_PN0P_  (.D(_00081_),
    .CK(clknet_leaf_81_clk),
    .Q(net116),
    .QN(_07314_));
 DFF_X1 \data_out_imag[119]$_SDFFE_PN0P_  (.D(_00082_),
    .CK(clknet_leaf_80_clk),
    .Q(net117),
    .QN(_07313_));
 DFF_X1 \data_out_imag[11]$_SDFFE_PN0P_  (.D(_00083_),
    .CK(clknet_leaf_80_clk),
    .Q(net118),
    .QN(_07312_));
 DFF_X1 \data_out_imag[120]$_SDFFE_PN0P_  (.D(_00084_),
    .CK(clknet_leaf_80_clk),
    .Q(net119),
    .QN(_07311_));
 DFF_X1 \data_out_imag[121]$_SDFFE_PN0P_  (.D(_00085_),
    .CK(clknet_leaf_81_clk),
    .Q(net120),
    .QN(_07310_));
 DFF_X1 \data_out_imag[122]$_SDFFE_PN0P_  (.D(_00086_),
    .CK(clknet_leaf_8_clk),
    .Q(net121),
    .QN(_07309_));
 DFF_X1 \data_out_imag[123]$_SDFFE_PN0P_  (.D(_00087_),
    .CK(clknet_leaf_80_clk),
    .Q(net122),
    .QN(_07308_));
 DFF_X1 \data_out_imag[124]$_SDFFE_PN0P_  (.D(_00088_),
    .CK(clknet_leaf_8_clk),
    .Q(net123),
    .QN(_07307_));
 DFF_X1 \data_out_imag[125]$_SDFFE_PN0P_  (.D(_00089_),
    .CK(clknet_leaf_9_clk),
    .Q(net124),
    .QN(_07306_));
 DFF_X1 \data_out_imag[126]$_SDFFE_PN0P_  (.D(_00090_),
    .CK(clknet_leaf_19_clk),
    .Q(net126),
    .QN(_07305_));
 DFF_X1 \data_out_imag[127]$_SDFFE_PN0P_  (.D(_00091_),
    .CK(clknet_leaf_19_clk),
    .Q(net127),
    .QN(_07304_));
 DFF_X1 \data_out_imag[12]$_SDFFE_PN0P_  (.D(_00092_),
    .CK(clknet_leaf_19_clk),
    .Q(net128),
    .QN(_07303_));
 DFF_X1 \data_out_imag[13]$_SDFFE_PN0P_  (.D(_00093_),
    .CK(clknet_leaf_20_clk),
    .Q(net134),
    .QN(_07302_));
 DFF_X1 \data_out_imag[14]$_SDFFE_PN0P_  (.D(_00094_),
    .CK(clknet_leaf_27_clk),
    .Q(net135),
    .QN(_07301_));
 DFF_X1 \data_out_imag[15]$_SDFFE_PN0P_  (.D(_00095_),
    .CK(clknet_leaf_30_clk),
    .Q(net136),
    .QN(_07300_));
 DFF_X1 \data_out_imag[16]$_SDFFE_PN0P_  (.D(_00096_),
    .CK(clknet_leaf_31_clk),
    .Q(net141),
    .QN(_07299_));
 DFF_X1 \data_out_imag[17]$_SDFFE_PN0P_  (.D(_00097_),
    .CK(clknet_leaf_29_clk),
    .Q(net142),
    .QN(_07298_));
 DFF_X1 \data_out_imag[18]$_SDFFE_PN0P_  (.D(_00098_),
    .CK(clknet_leaf_31_clk),
    .Q(net145),
    .QN(_07297_));
 DFF_X1 \data_out_imag[19]$_SDFFE_PN0P_  (.D(_00099_),
    .CK(clknet_leaf_30_clk),
    .Q(net146),
    .QN(_07296_));
 DFF_X1 \data_out_imag[1]$_SDFFE_PN0P_  (.D(_00100_),
    .CK(clknet_leaf_29_clk),
    .Q(net147),
    .QN(_07295_));
 DFF_X1 \data_out_imag[20]$_SDFFE_PN0P_  (.D(_00101_),
    .CK(clknet_leaf_28_clk),
    .Q(net148),
    .QN(_07294_));
 DFF_X1 \data_out_imag[21]$_SDFFE_PN0P_  (.D(_00102_),
    .CK(clknet_leaf_28_clk),
    .Q(net150),
    .QN(_07293_));
 DFF_X1 \data_out_imag[22]$_SDFFE_PN0P_  (.D(_00103_),
    .CK(clknet_leaf_27_clk),
    .Q(net155),
    .QN(_07292_));
 DFF_X1 \data_out_imag[23]$_SDFFE_PN0P_  (.D(_00104_),
    .CK(clknet_leaf_22_clk),
    .Q(net157),
    .QN(_07291_));
 DFF_X1 \data_out_imag[24]$_SDFFE_PN0P_  (.D(_00105_),
    .CK(clknet_leaf_20_clk),
    .Q(net159),
    .QN(_07290_));
 DFF_X1 \data_out_imag[25]$_SDFFE_PN0P_  (.D(_00106_),
    .CK(clknet_leaf_21_clk),
    .Q(net160),
    .QN(_07289_));
 DFF_X1 \data_out_imag[26]$_SDFFE_PN0P_  (.D(_00107_),
    .CK(clknet_leaf_20_clk),
    .Q(net161),
    .QN(_07288_));
 DFF_X1 \data_out_imag[27]$_SDFFE_PN0P_  (.D(_00108_),
    .CK(clknet_leaf_20_clk),
    .Q(net162),
    .QN(_07287_));
 DFF_X1 \data_out_imag[28]$_SDFFE_PN0P_  (.D(_00109_),
    .CK(clknet_leaf_20_clk),
    .Q(net163),
    .QN(_07286_));
 DFF_X1 \data_out_imag[29]$_SDFFE_PN0P_  (.D(_00110_),
    .CK(clknet_leaf_21_clk),
    .Q(net164),
    .QN(_07285_));
 DFF_X1 \data_out_imag[2]$_SDFFE_PN0P_  (.D(_00111_),
    .CK(clknet_leaf_31_clk),
    .Q(net165),
    .QN(_07284_));
 DFF_X1 \data_out_imag[30]$_SDFFE_PN0P_  (.D(_00112_),
    .CK(clknet_leaf_27_clk),
    .Q(net166),
    .QN(_07283_));
 DFF_X1 \data_out_imag[31]$_SDFFE_PN0P_  (.D(_00113_),
    .CK(clknet_leaf_31_clk),
    .Q(net167),
    .QN(_07282_));
 DFF_X1 \data_out_imag[32]$_SDFFE_PN0P_  (.D(_00114_),
    .CK(clknet_leaf_28_clk),
    .Q(net168),
    .QN(_07281_));
 DFF_X1 \data_out_imag[33]$_SDFFE_PN0P_  (.D(_00115_),
    .CK(clknet_leaf_28_clk),
    .Q(net169),
    .QN(_07280_));
 DFF_X1 \data_out_imag[34]$_SDFFE_PN0P_  (.D(_00116_),
    .CK(clknet_leaf_31_clk),
    .Q(net170),
    .QN(_07279_));
 DFF_X1 \data_out_imag[35]$_SDFFE_PN0P_  (.D(_00117_),
    .CK(clknet_leaf_31_clk),
    .Q(net171),
    .QN(_07278_));
 DFF_X1 \data_out_imag[36]$_SDFFE_PN0P_  (.D(_00118_),
    .CK(clknet_leaf_29_clk),
    .Q(net172),
    .QN(_07277_));
 DFF_X1 \data_out_imag[37]$_SDFFE_PN0P_  (.D(_00119_),
    .CK(clknet_leaf_28_clk),
    .Q(net173),
    .QN(_07276_));
 DFF_X1 \data_out_imag[38]$_SDFFE_PN0P_  (.D(_00120_),
    .CK(clknet_leaf_27_clk),
    .Q(net174),
    .QN(_07275_));
 DFF_X1 \data_out_imag[39]$_SDFFE_PN0P_  (.D(_00121_),
    .CK(clknet_leaf_21_clk),
    .Q(net175),
    .QN(_07274_));
 DFF_X1 \data_out_imag[3]$_SDFFE_PN0P_  (.D(_00122_),
    .CK(clknet_leaf_28_clk),
    .Q(net176),
    .QN(_07273_));
 DFF_X1 \data_out_imag[40]$_SDFFE_PN0P_  (.D(_00123_),
    .CK(clknet_leaf_21_clk),
    .Q(net177),
    .QN(_07272_));
 DFF_X1 \data_out_imag[41]$_SDFFE_PN0P_  (.D(_00124_),
    .CK(clknet_leaf_21_clk),
    .Q(net178),
    .QN(_07271_));
 DFF_X1 \data_out_imag[42]$_SDFFE_PN0P_  (.D(_00125_),
    .CK(clknet_leaf_21_clk),
    .Q(net179),
    .QN(_07270_));
 DFF_X1 \data_out_imag[43]$_SDFFE_PN0P_  (.D(_00126_),
    .CK(clknet_leaf_20_clk),
    .Q(net180),
    .QN(_07269_));
 DFF_X1 \data_out_imag[44]$_SDFFE_PN0P_  (.D(_00127_),
    .CK(clknet_leaf_20_clk),
    .Q(net181),
    .QN(_07268_));
 DFF_X1 \data_out_imag[45]$_SDFFE_PN0P_  (.D(_00128_),
    .CK(clknet_leaf_21_clk),
    .Q(net182),
    .QN(_07267_));
 DFF_X1 \data_out_imag[46]$_SDFFE_PN0P_  (.D(_00129_),
    .CK(clknet_leaf_27_clk),
    .Q(net183),
    .QN(_07266_));
 DFF_X1 \data_out_imag[47]$_SDFFE_PN0P_  (.D(_00130_),
    .CK(clknet_leaf_30_clk),
    .Q(net184),
    .QN(_07265_));
 DFF_X1 \data_out_imag[48]$_SDFFE_PN0P_  (.D(_00131_),
    .CK(clknet_leaf_30_clk),
    .Q(net185),
    .QN(_07264_));
 DFF_X1 \data_out_imag[49]$_SDFFE_PN0P_  (.D(_00132_),
    .CK(clknet_leaf_29_clk),
    .Q(net186),
    .QN(_07263_));
 DFF_X1 \data_out_imag[4]$_SDFFE_PN0P_  (.D(_00133_),
    .CK(clknet_leaf_28_clk),
    .Q(net187),
    .QN(_07262_));
 DFF_X1 \data_out_imag[50]$_SDFFE_PN0P_  (.D(_00134_),
    .CK(clknet_leaf_30_clk),
    .Q(net188),
    .QN(_07261_));
 DFF_X1 \data_out_imag[51]$_SDFFE_PN0P_  (.D(_00135_),
    .CK(clknet_leaf_29_clk),
    .Q(net189),
    .QN(_07260_));
 DFF_X1 \data_out_imag[52]$_SDFFE_PN0P_  (.D(_00136_),
    .CK(clknet_leaf_26_clk),
    .Q(net190),
    .QN(_07259_));
 DFF_X1 \data_out_imag[53]$_SDFFE_PN0P_  (.D(_00137_),
    .CK(clknet_leaf_29_clk),
    .Q(net191),
    .QN(_07258_));
 DFF_X1 \data_out_imag[54]$_SDFFE_PN0P_  (.D(_00138_),
    .CK(clknet_leaf_22_clk),
    .Q(net192),
    .QN(_07257_));
 DFF_X1 \data_out_imag[55]$_SDFFE_PN0P_  (.D(_00139_),
    .CK(clknet_leaf_22_clk),
    .Q(net193),
    .QN(_07256_));
 DFF_X1 \data_out_imag[56]$_SDFFE_PN0P_  (.D(_00140_),
    .CK(clknet_leaf_18_clk),
    .Q(net194),
    .QN(_07255_));
 DFF_X1 \data_out_imag[57]$_SDFFE_PN0P_  (.D(_00141_),
    .CK(clknet_leaf_19_clk),
    .Q(net195),
    .QN(_07254_));
 DFF_X1 \data_out_imag[58]$_SDFFE_PN0P_  (.D(_00142_),
    .CK(clknet_leaf_18_clk),
    .Q(net196),
    .QN(_07253_));
 DFF_X1 \data_out_imag[59]$_SDFFE_PN0P_  (.D(_00143_),
    .CK(clknet_leaf_18_clk),
    .Q(net197),
    .QN(_07252_));
 DFF_X1 \data_out_imag[5]$_SDFFE_PN0P_  (.D(_00144_),
    .CK(clknet_leaf_17_clk),
    .Q(net198),
    .QN(_07251_));
 DFF_X1 \data_out_imag[60]$_SDFFE_PN0P_  (.D(_00145_),
    .CK(clknet_leaf_17_clk),
    .Q(net199),
    .QN(_07250_));
 DFF_X1 \data_out_imag[61]$_SDFFE_PN0P_  (.D(_00146_),
    .CK(clknet_leaf_17_clk),
    .Q(net200),
    .QN(_07249_));
 DFF_X1 \data_out_imag[62]$_SDFFE_PN0P_  (.D(_00147_),
    .CK(clknet_leaf_17_clk),
    .Q(net201),
    .QN(_07248_));
 DFF_X1 \data_out_imag[63]$_SDFFE_PN0P_  (.D(_00148_),
    .CK(clknet_leaf_18_clk),
    .Q(net202),
    .QN(_07247_));
 DFF_X1 \data_out_imag[64]$_SDFFE_PN0P_  (.D(_00149_),
    .CK(clknet_leaf_18_clk),
    .Q(net203),
    .QN(_07246_));
 DFF_X1 \data_out_imag[65]$_SDFFE_PN0P_  (.D(_00150_),
    .CK(clknet_leaf_11_clk),
    .Q(net204),
    .QN(_07245_));
 DFF_X1 \data_out_imag[66]$_SDFFE_PN0P_  (.D(_00151_),
    .CK(clknet_leaf_10_clk),
    .Q(net205),
    .QN(_07244_));
 DFF_X1 \data_out_imag[67]$_SDFFE_PN0P_  (.D(_00152_),
    .CK(clknet_leaf_10_clk),
    .Q(net206),
    .QN(_07243_));
 DFF_X1 \data_out_imag[68]$_SDFFE_PN0P_  (.D(_00153_),
    .CK(clknet_leaf_9_clk),
    .Q(net207),
    .QN(_07242_));
 DFF_X1 \data_out_imag[69]$_SDFFE_PN0P_  (.D(_00154_),
    .CK(clknet_leaf_9_clk),
    .Q(net208),
    .QN(_07241_));
 DFF_X1 \data_out_imag[6]$_SDFFE_PN0P_  (.D(_00155_),
    .CK(clknet_leaf_9_clk),
    .Q(net209),
    .QN(_07240_));
 DFF_X1 \data_out_imag[70]$_SDFFE_PN0P_  (.D(_00156_),
    .CK(clknet_leaf_9_clk),
    .Q(net210),
    .QN(_07239_));
 DFF_X1 \data_out_imag[71]$_SDFFE_PN0P_  (.D(_00157_),
    .CK(clknet_leaf_9_clk),
    .Q(net211),
    .QN(_07238_));
 DFF_X1 \data_out_imag[72]$_SDFFE_PN0P_  (.D(_00158_),
    .CK(clknet_leaf_9_clk),
    .Q(net212),
    .QN(_07237_));
 DFF_X1 \data_out_imag[73]$_SDFFE_PN0P_  (.D(_00159_),
    .CK(clknet_leaf_9_clk),
    .Q(net213),
    .QN(_07236_));
 DFF_X1 \data_out_imag[74]$_SDFFE_PN0P_  (.D(_00160_),
    .CK(clknet_leaf_10_clk),
    .Q(net214),
    .QN(_07235_));
 DFF_X1 \data_out_imag[75]$_SDFFE_PN0P_  (.D(_00161_),
    .CK(clknet_leaf_10_clk),
    .Q(net215),
    .QN(_07234_));
 DFF_X1 \data_out_imag[76]$_SDFFE_PN0P_  (.D(_00162_),
    .CK(clknet_leaf_10_clk),
    .Q(net216),
    .QN(_07233_));
 DFF_X1 \data_out_imag[77]$_SDFFE_PN0P_  (.D(_00163_),
    .CK(clknet_leaf_10_clk),
    .Q(net217),
    .QN(_07232_));
 DFF_X1 \data_out_imag[78]$_SDFFE_PN0P_  (.D(_00164_),
    .CK(clknet_leaf_11_clk),
    .Q(net218),
    .QN(_07231_));
 DFF_X1 \data_out_imag[79]$_SDFFE_PN0P_  (.D(_00165_),
    .CK(clknet_leaf_11_clk),
    .Q(net219),
    .QN(_07230_));
 DFF_X1 \data_out_imag[7]$_SDFFE_PN0P_  (.D(_00166_),
    .CK(clknet_leaf_11_clk),
    .Q(net220),
    .QN(_07229_));
 DFF_X1 \data_out_imag[80]$_SDFFE_PN0P_  (.D(_00167_),
    .CK(clknet_leaf_12_clk),
    .Q(net221),
    .QN(_07228_));
 DFF_X1 \data_out_imag[81]$_SDFFE_PN0P_  (.D(_00168_),
    .CK(clknet_leaf_11_clk),
    .Q(net222),
    .QN(_07227_));
 DFF_X1 \data_out_imag[82]$_SDFFE_PN0P_  (.D(_00169_),
    .CK(clknet_leaf_11_clk),
    .Q(net223),
    .QN(_07226_));
 DFF_X1 \data_out_imag[83]$_SDFFE_PN0P_  (.D(_00170_),
    .CK(clknet_leaf_11_clk),
    .Q(net224),
    .QN(_07225_));
 DFF_X1 \data_out_imag[84]$_SDFFE_PN0P_  (.D(_00171_),
    .CK(clknet_leaf_16_clk),
    .Q(net225),
    .QN(_07224_));
 DFF_X1 \data_out_imag[85]$_SDFFE_PN0P_  (.D(_00172_),
    .CK(clknet_leaf_11_clk),
    .Q(net226),
    .QN(_07223_));
 DFF_X1 \data_out_imag[86]$_SDFFE_PN0P_  (.D(_00173_),
    .CK(clknet_leaf_12_clk),
    .Q(net227),
    .QN(_07222_));
 DFF_X1 \data_out_imag[87]$_SDFFE_PN0P_  (.D(_00174_),
    .CK(clknet_leaf_16_clk),
    .Q(net228),
    .QN(_07221_));
 DFF_X1 \data_out_imag[88]$_SDFFE_PN0P_  (.D(_00175_),
    .CK(clknet_leaf_17_clk),
    .Q(net229),
    .QN(_07220_));
 DFF_X1 \data_out_imag[89]$_SDFFE_PN0P_  (.D(_00176_),
    .CK(clknet_leaf_16_clk),
    .Q(net230),
    .QN(_07219_));
 DFF_X1 \data_out_imag[8]$_SDFFE_PN0P_  (.D(_00177_),
    .CK(clknet_leaf_17_clk),
    .Q(net231),
    .QN(_07218_));
 DFF_X1 \data_out_imag[90]$_SDFFE_PN0P_  (.D(_00178_),
    .CK(clknet_leaf_16_clk),
    .Q(net232),
    .QN(_07217_));
 DFF_X1 \data_out_imag[91]$_SDFFE_PN0P_  (.D(_00179_),
    .CK(clknet_leaf_17_clk),
    .Q(net233),
    .QN(_07216_));
 DFF_X1 \data_out_imag[92]$_SDFFE_PN0P_  (.D(_00180_),
    .CK(clknet_leaf_16_clk),
    .Q(net234),
    .QN(_07215_));
 DFF_X1 \data_out_imag[93]$_SDFFE_PN0P_  (.D(_00181_),
    .CK(clknet_leaf_18_clk),
    .Q(net235),
    .QN(_07214_));
 DFF_X1 \data_out_imag[94]$_SDFFE_PN0P_  (.D(_00182_),
    .CK(clknet_leaf_17_clk),
    .Q(net236),
    .QN(_07213_));
 DFF_X1 \data_out_imag[95]$_SDFFE_PN0P_  (.D(_00183_),
    .CK(clknet_leaf_16_clk),
    .Q(net237),
    .QN(_07212_));
 DFF_X1 \data_out_imag[96]$_SDFFE_PN0P_  (.D(_00184_),
    .CK(clknet_leaf_27_clk),
    .Q(net238),
    .QN(_07211_));
 DFF_X1 \data_out_imag[97]$_SDFFE_PN0P_  (.D(_00185_),
    .CK(clknet_leaf_12_clk),
    .Q(net239),
    .QN(_07210_));
 DFF_X1 \data_out_imag[98]$_SDFFE_PN0P_  (.D(_00186_),
    .CK(clknet_leaf_16_clk),
    .Q(net240),
    .QN(_07209_));
 DFF_X1 \data_out_imag[99]$_SDFFE_PN0P_  (.D(_00187_),
    .CK(clknet_leaf_12_clk),
    .Q(net241),
    .QN(_07208_));
 DFF_X1 \data_out_imag[9]$_SDFFE_PN0P_  (.D(_00188_),
    .CK(clknet_leaf_27_clk),
    .Q(net242),
    .QN(_07207_));
 DFF_X1 \data_out_real[0]$_SDFFE_PN0P_  (.D(_00189_),
    .CK(clknet_leaf_32_clk),
    .Q(net243),
    .QN(_07206_));
 DFF_X1 \data_out_real[100]$_SDFFE_PN0P_  (.D(_00190_),
    .CK(clknet_leaf_62_clk),
    .Q(net244),
    .QN(_07205_));
 DFF_X1 \data_out_real[101]$_SDFFE_PN0P_  (.D(_00191_),
    .CK(clknet_leaf_62_clk),
    .Q(net245),
    .QN(_07204_));
 DFF_X1 \data_out_real[102]$_SDFFE_PN0P_  (.D(_00192_),
    .CK(clknet_leaf_62_clk),
    .Q(net246),
    .QN(_07203_));
 DFF_X1 \data_out_real[103]$_SDFFE_PN0P_  (.D(_00193_),
    .CK(clknet_leaf_61_clk),
    .Q(net247),
    .QN(_07202_));
 DFF_X1 \data_out_real[104]$_SDFFE_PN0P_  (.D(_00194_),
    .CK(clknet_leaf_61_clk),
    .Q(net248),
    .QN(_07201_));
 DFF_X1 \data_out_real[105]$_SDFFE_PN0P_  (.D(_00195_),
    .CK(clknet_leaf_62_clk),
    .Q(net249),
    .QN(_07200_));
 DFF_X1 \data_out_real[106]$_SDFFE_PN0P_  (.D(_00196_),
    .CK(clknet_leaf_61_clk),
    .Q(net250),
    .QN(_07199_));
 DFF_X1 \data_out_real[107]$_SDFFE_PN0P_  (.D(_00197_),
    .CK(clknet_leaf_57_clk),
    .Q(net251),
    .QN(_07198_));
 DFF_X1 \data_out_real[108]$_SDFFE_PN0P_  (.D(_00198_),
    .CK(clknet_leaf_61_clk),
    .Q(net252),
    .QN(_07197_));
 DFF_X1 \data_out_real[109]$_SDFFE_PN0P_  (.D(_00199_),
    .CK(clknet_leaf_61_clk),
    .Q(net253),
    .QN(_07196_));
 DFF_X1 \data_out_real[10]$_SDFFE_PN0P_  (.D(_00200_),
    .CK(clknet_leaf_57_clk),
    .Q(net254),
    .QN(_07195_));
 DFF_X1 \data_out_real[110]$_SDFFE_PN0P_  (.D(_00201_),
    .CK(clknet_leaf_58_clk),
    .Q(net255),
    .QN(_07194_));
 DFF_X1 \data_out_real[111]$_SDFFE_PN0P_  (.D(_00202_),
    .CK(clknet_leaf_58_clk),
    .Q(net256),
    .QN(_07193_));
 DFF_X1 \data_out_real[112]$_SDFFE_PN0P_  (.D(_00203_),
    .CK(clknet_leaf_59_clk),
    .Q(net257),
    .QN(_07192_));
 DFF_X1 \data_out_real[113]$_SDFFE_PN0P_  (.D(_00204_),
    .CK(clknet_leaf_59_clk),
    .Q(net258),
    .QN(_07191_));
 DFF_X1 \data_out_real[114]$_SDFFE_PN0P_  (.D(_00205_),
    .CK(clknet_leaf_58_clk),
    .Q(net259),
    .QN(_07190_));
 DFF_X1 \data_out_real[115]$_SDFFE_PN0P_  (.D(_00206_),
    .CK(clknet_leaf_59_clk),
    .Q(net260),
    .QN(_07189_));
 DFF_X1 \data_out_real[116]$_SDFFE_PN0P_  (.D(_00207_),
    .CK(clknet_leaf_58_clk),
    .Q(net261),
    .QN(_07188_));
 DFF_X1 \data_out_real[117]$_SDFFE_PN0P_  (.D(_00208_),
    .CK(clknet_leaf_59_clk),
    .Q(net262),
    .QN(_07187_));
 DFF_X1 \data_out_real[118]$_SDFFE_PN0P_  (.D(_00209_),
    .CK(clknet_leaf_58_clk),
    .Q(net263),
    .QN(_07186_));
 DFF_X1 \data_out_real[119]$_SDFFE_PN0P_  (.D(_00210_),
    .CK(clknet_leaf_58_clk),
    .Q(net264),
    .QN(_07185_));
 DFF_X1 \data_out_real[11]$_SDFFE_PN0P_  (.D(_00211_),
    .CK(clknet_leaf_56_clk),
    .Q(net265),
    .QN(_07184_));
 DFF_X1 \data_out_real[120]$_SDFFE_PN0P_  (.D(_00212_),
    .CK(clknet_leaf_56_clk),
    .Q(net266),
    .QN(_07183_));
 DFF_X1 \data_out_real[121]$_SDFFE_PN0P_  (.D(_00213_),
    .CK(clknet_leaf_56_clk),
    .Q(net267),
    .QN(_07182_));
 DFF_X1 \data_out_real[122]$_SDFFE_PN0P_  (.D(_00214_),
    .CK(clknet_leaf_55_clk),
    .Q(net268),
    .QN(_07181_));
 DFF_X1 \data_out_real[123]$_SDFFE_PN0P_  (.D(_00215_),
    .CK(clknet_leaf_55_clk),
    .Q(net269),
    .QN(_07180_));
 DFF_X1 \data_out_real[124]$_SDFFE_PN0P_  (.D(_00216_),
    .CK(clknet_leaf_56_clk),
    .Q(net270),
    .QN(_07179_));
 DFF_X1 \data_out_real[125]$_SDFFE_PN0P_  (.D(_00217_),
    .CK(clknet_leaf_55_clk),
    .Q(net271),
    .QN(_07178_));
 DFF_X1 \data_out_real[126]$_SDFFE_PN0P_  (.D(_00218_),
    .CK(clknet_leaf_56_clk),
    .Q(net272),
    .QN(_07177_));
 DFF_X1 \data_out_real[127]$_SDFFE_PN0P_  (.D(_00219_),
    .CK(clknet_leaf_55_clk),
    .Q(net273),
    .QN(_07176_));
 DFF_X1 \data_out_real[12]$_SDFFE_PN0P_  (.D(_00220_),
    .CK(clknet_leaf_55_clk),
    .Q(net274),
    .QN(_07175_));
 DFF_X1 \data_out_real[13]$_SDFFE_PN0P_  (.D(_00221_),
    .CK(clknet_leaf_55_clk),
    .Q(net275),
    .QN(_07174_));
 DFF_X1 \data_out_real[14]$_SDFFE_PN0P_  (.D(_00222_),
    .CK(clknet_leaf_54_clk),
    .Q(net276),
    .QN(_07173_));
 DFF_X1 \data_out_real[15]$_SDFFE_PN0P_  (.D(_00223_),
    .CK(clknet_leaf_54_clk),
    .Q(net277),
    .QN(_07172_));
 DFF_X1 \data_out_real[16]$_SDFFE_PN0P_  (.D(_00224_),
    .CK(clknet_leaf_50_clk),
    .Q(net278),
    .QN(_07171_));
 DFF_X1 \data_out_real[17]$_SDFFE_PN0P_  (.D(_00225_),
    .CK(clknet_leaf_50_clk),
    .Q(net279),
    .QN(_07170_));
 DFF_X1 \data_out_real[18]$_SDFFE_PN0P_  (.D(_00226_),
    .CK(clknet_leaf_50_clk),
    .Q(net280),
    .QN(_07169_));
 DFF_X1 \data_out_real[19]$_SDFFE_PN0P_  (.D(_00227_),
    .CK(clknet_leaf_50_clk),
    .Q(net281),
    .QN(_07168_));
 DFF_X1 \data_out_real[1]$_SDFFE_PN0P_  (.D(_00228_),
    .CK(clknet_leaf_49_clk),
    .Q(net282),
    .QN(_07167_));
 DFF_X1 \data_out_real[20]$_SDFFE_PN0P_  (.D(_00229_),
    .CK(clknet_leaf_49_clk),
    .Q(net283),
    .QN(_07166_));
 DFF_X1 \data_out_real[21]$_SDFFE_PN0P_  (.D(_00230_),
    .CK(clknet_leaf_48_clk),
    .Q(net284),
    .QN(_07165_));
 DFF_X1 \data_out_real[22]$_SDFFE_PN0P_  (.D(_00231_),
    .CK(clknet_leaf_44_clk),
    .Q(net285),
    .QN(_07164_));
 DFF_X1 \data_out_real[23]$_SDFFE_PN0P_  (.D(_00232_),
    .CK(clknet_leaf_45_clk),
    .Q(net286),
    .QN(_07163_));
 DFF_X1 \data_out_real[24]$_SDFFE_PN0P_  (.D(_00233_),
    .CK(clknet_leaf_45_clk),
    .Q(net287),
    .QN(_07162_));
 DFF_X1 \data_out_real[25]$_SDFFE_PN0P_  (.D(_00234_),
    .CK(clknet_leaf_32_clk),
    .Q(net288),
    .QN(_07161_));
 DFF_X1 \data_out_real[26]$_SDFFE_PN0P_  (.D(_00235_),
    .CK(clknet_leaf_46_clk),
    .Q(net289),
    .QN(_07160_));
 DFF_X1 \data_out_real[27]$_SDFFE_PN0P_  (.D(_00236_),
    .CK(clknet_leaf_49_clk),
    .Q(net290),
    .QN(_07159_));
 DFF_X1 \data_out_real[28]$_SDFFE_PN0P_  (.D(_00237_),
    .CK(clknet_leaf_48_clk),
    .Q(net291),
    .QN(_07158_));
 DFF_X1 \data_out_real[29]$_SDFFE_PN0P_  (.D(_00238_),
    .CK(clknet_leaf_48_clk),
    .Q(net292),
    .QN(_07157_));
 DFF_X1 \data_out_real[2]$_SDFFE_PN0P_  (.D(_00239_),
    .CK(clknet_leaf_32_clk),
    .Q(net293),
    .QN(_07156_));
 DFF_X1 \data_out_real[30]$_SDFFE_PN0P_  (.D(_00240_),
    .CK(clknet_leaf_49_clk),
    .Q(net294),
    .QN(_07155_));
 DFF_X1 \data_out_real[31]$_SDFFE_PN0P_  (.D(_00241_),
    .CK(clknet_leaf_31_clk),
    .Q(net295),
    .QN(_07154_));
 DFF_X1 \data_out_real[32]$_SDFFE_PN0P_  (.D(_00242_),
    .CK(clknet_leaf_46_clk),
    .Q(net296),
    .QN(_07153_));
 DFF_X1 \data_out_real[33]$_SDFFE_PN0P_  (.D(_00243_),
    .CK(clknet_leaf_48_clk),
    .Q(net297),
    .QN(_07152_));
 DFF_X1 \data_out_real[34]$_SDFFE_PN0P_  (.D(_00244_),
    .CK(clknet_leaf_32_clk),
    .Q(net298),
    .QN(_07151_));
 DFF_X1 \data_out_real[35]$_SDFFE_PN0P_  (.D(_00245_),
    .CK(clknet_leaf_47_clk),
    .Q(net299),
    .QN(_07150_));
 DFF_X1 \data_out_real[36]$_SDFFE_PN0P_  (.D(_00246_),
    .CK(clknet_leaf_46_clk),
    .Q(net300),
    .QN(_07149_));
 DFF_X1 \data_out_real[37]$_SDFFE_PN0P_  (.D(_00247_),
    .CK(clknet_leaf_47_clk),
    .Q(net301),
    .QN(_07148_));
 DFF_X1 \data_out_real[38]$_SDFFE_PN0P_  (.D(_00248_),
    .CK(clknet_leaf_32_clk),
    .Q(net302),
    .QN(_07147_));
 DFF_X1 \data_out_real[39]$_SDFFE_PN0P_  (.D(_00249_),
    .CK(clknet_leaf_46_clk),
    .Q(net303),
    .QN(_07146_));
 DFF_X1 \data_out_real[3]$_SDFFE_PN0P_  (.D(_00250_),
    .CK(clknet_leaf_47_clk),
    .Q(net304),
    .QN(_07145_));
 DFF_X1 \data_out_real[40]$_SDFFE_PN0P_  (.D(_00251_),
    .CK(clknet_leaf_45_clk),
    .Q(net305),
    .QN(_07144_));
 DFF_X1 \data_out_real[41]$_SDFFE_PN0P_  (.D(_00252_),
    .CK(clknet_leaf_44_clk),
    .Q(net306),
    .QN(_07143_));
 DFF_X1 \data_out_real[42]$_SDFFE_PN0P_  (.D(_00253_),
    .CK(clknet_leaf_46_clk),
    .Q(net307),
    .QN(_07142_));
 DFF_X1 \data_out_real[43]$_SDFFE_PN0P_  (.D(_00254_),
    .CK(clknet_leaf_55_clk),
    .Q(net308),
    .QN(_07141_));
 DFF_X1 \data_out_real[44]$_SDFFE_PN0P_  (.D(_00255_),
    .CK(clknet_leaf_49_clk),
    .Q(net309),
    .QN(_07140_));
 DFF_X1 \data_out_real[45]$_SDFFE_PN0P_  (.D(_00256_),
    .CK(clknet_leaf_49_clk),
    .Q(net310),
    .QN(_07139_));
 DFF_X1 \data_out_real[46]$_SDFFE_PN0P_  (.D(_00257_),
    .CK(clknet_leaf_49_clk),
    .Q(net311),
    .QN(_07138_));
 DFF_X1 \data_out_real[47]$_SDFFE_PN0P_  (.D(_00258_),
    .CK(clknet_leaf_32_clk),
    .Q(net312),
    .QN(_07137_));
 DFF_X1 \data_out_real[48]$_SDFFE_PN0P_  (.D(_00259_),
    .CK(clknet_leaf_47_clk),
    .Q(net313),
    .QN(_07136_));
 DFF_X1 \data_out_real[49]$_SDFFE_PN0P_  (.D(_00260_),
    .CK(clknet_leaf_48_clk),
    .Q(net314),
    .QN(_07135_));
 DFF_X1 \data_out_real[4]$_SDFFE_PN0P_  (.D(_00261_),
    .CK(clknet_leaf_46_clk),
    .Q(net315),
    .QN(_07134_));
 DFF_X1 \data_out_real[50]$_SDFFE_PN0P_  (.D(_00262_),
    .CK(clknet_leaf_45_clk),
    .Q(net316),
    .QN(_07133_));
 DFF_X1 \data_out_real[51]$_SDFFE_PN0P_  (.D(_00263_),
    .CK(clknet_leaf_48_clk),
    .Q(net317),
    .QN(_07132_));
 DFF_X1 \data_out_real[52]$_SDFFE_PN0P_  (.D(_00264_),
    .CK(clknet_leaf_46_clk),
    .Q(net318),
    .QN(_07131_));
 DFF_X1 \data_out_real[53]$_SDFFE_PN0P_  (.D(_00265_),
    .CK(clknet_leaf_48_clk),
    .Q(net319),
    .QN(_07130_));
 DFF_X1 \data_out_real[54]$_SDFFE_PN0P_  (.D(_00266_),
    .CK(clknet_leaf_45_clk),
    .Q(net320),
    .QN(_07129_));
 DFF_X1 \data_out_real[55]$_SDFFE_PN0P_  (.D(_00267_),
    .CK(clknet_leaf_45_clk),
    .Q(net321),
    .QN(_07128_));
 DFF_X1 \data_out_real[56]$_SDFFE_PN0P_  (.D(_00268_),
    .CK(clknet_leaf_45_clk),
    .Q(net322),
    .QN(_07127_));
 DFF_X1 \data_out_real[57]$_SDFFE_PN0P_  (.D(_00269_),
    .CK(clknet_leaf_45_clk),
    .Q(net323),
    .QN(_07126_));
 DFF_X1 \data_out_real[58]$_SDFFE_PN0P_  (.D(_00270_),
    .CK(clknet_leaf_59_clk),
    .Q(net324),
    .QN(_07125_));
 DFF_X1 \data_out_real[59]$_SDFFE_PN0P_  (.D(_00271_),
    .CK(clknet_leaf_56_clk),
    .Q(net325),
    .QN(_07124_));
 DFF_X1 \data_out_real[5]$_SDFFE_PN0P_  (.D(_00272_),
    .CK(clknet_leaf_59_clk),
    .Q(net326),
    .QN(_07123_));
 DFF_X1 \data_out_real[60]$_SDFFE_PN0P_  (.D(_00273_),
    .CK(clknet_leaf_59_clk),
    .Q(net327),
    .QN(_07122_));
 DFF_X1 \data_out_real[61]$_SDFFE_PN0P_  (.D(_00274_),
    .CK(clknet_leaf_60_clk),
    .Q(net328),
    .QN(_07121_));
 DFF_X1 \data_out_real[62]$_SDFFE_PN0P_  (.D(_00275_),
    .CK(clknet_leaf_56_clk),
    .Q(net329),
    .QN(_07120_));
 DFF_X1 \data_out_real[63]$_SDFFE_PN0P_  (.D(_00276_),
    .CK(clknet_leaf_57_clk),
    .Q(net330),
    .QN(_07119_));
 DFF_X1 \data_out_real[64]$_SDFFE_PN0P_  (.D(_00277_),
    .CK(clknet_leaf_59_clk),
    .Q(net331),
    .QN(_07118_));
 DFF_X1 \data_out_real[65]$_SDFFE_PN0P_  (.D(_00278_),
    .CK(clknet_leaf_56_clk),
    .Q(net332),
    .QN(_07117_));
 DFF_X1 \data_out_real[66]$_SDFFE_PN0P_  (.D(_00279_),
    .CK(clknet_leaf_60_clk),
    .Q(net333),
    .QN(_07116_));
 DFF_X1 \data_out_real[67]$_SDFFE_PN0P_  (.D(_00280_),
    .CK(clknet_leaf_57_clk),
    .Q(net334),
    .QN(_07115_));
 DFF_X1 \data_out_real[68]$_SDFFE_PN0P_  (.D(_00281_),
    .CK(clknet_leaf_60_clk),
    .Q(net335),
    .QN(_07114_));
 DFF_X1 \data_out_real[69]$_SDFFE_PN0P_  (.D(_00282_),
    .CK(clknet_leaf_58_clk),
    .Q(net336),
    .QN(_07113_));
 DFF_X1 \data_out_real[6]$_SDFFE_PN0P_  (.D(_00283_),
    .CK(clknet_leaf_60_clk),
    .Q(net337),
    .QN(_07112_));
 DFF_X1 \data_out_real[70]$_SDFFE_PN0P_  (.D(_00284_),
    .CK(clknet_leaf_57_clk),
    .Q(net338),
    .QN(_07111_));
 DFF_X1 \data_out_real[71]$_SDFFE_PN0P_  (.D(_00285_),
    .CK(clknet_leaf_54_clk),
    .Q(net339),
    .QN(_07110_));
 DFF_X1 \data_out_real[72]$_SDFFE_PN0P_  (.D(_00286_),
    .CK(clknet_leaf_60_clk),
    .Q(net340),
    .QN(_07109_));
 DFF_X1 \data_out_real[73]$_SDFFE_PN0P_  (.D(_00287_),
    .CK(clknet_leaf_54_clk),
    .Q(net341),
    .QN(_07108_));
 DFF_X1 \data_out_real[74]$_SDFFE_PN0P_  (.D(_00288_),
    .CK(clknet_leaf_57_clk),
    .Q(net342),
    .QN(_07107_));
 DFF_X1 \data_out_real[75]$_SDFFE_PN0P_  (.D(_00289_),
    .CK(clknet_leaf_60_clk),
    .Q(net343),
    .QN(_07106_));
 DFF_X1 \data_out_real[76]$_SDFFE_PN0P_  (.D(_00290_),
    .CK(clknet_leaf_57_clk),
    .Q(net344),
    .QN(_07105_));
 DFF_X1 \data_out_real[77]$_SDFFE_PN0P_  (.D(_00291_),
    .CK(clknet_leaf_54_clk),
    .Q(net345),
    .QN(_07104_));
 DFF_X1 \data_out_real[78]$_SDFFE_PN0P_  (.D(_00292_),
    .CK(clknet_leaf_60_clk),
    .Q(net346),
    .QN(_07103_));
 DFF_X1 \data_out_real[79]$_SDFFE_PN0P_  (.D(_00293_),
    .CK(clknet_leaf_61_clk),
    .Q(net347),
    .QN(_07102_));
 DFF_X1 \data_out_real[7]$_SDFFE_PN0P_  (.D(_00294_),
    .CK(clknet_leaf_61_clk),
    .Q(net348),
    .QN(_07101_));
 DFF_X1 \data_out_real[80]$_SDFFE_PN0P_  (.D(_00295_),
    .CK(clknet_leaf_53_clk),
    .Q(net349),
    .QN(_07100_));
 DFF_X1 \data_out_real[81]$_SDFFE_PN0P_  (.D(_00296_),
    .CK(clknet_leaf_63_clk),
    .Q(net350),
    .QN(_07099_));
 DFF_X1 \data_out_real[82]$_SDFFE_PN0P_  (.D(_00297_),
    .CK(clknet_leaf_62_clk),
    .Q(net351),
    .QN(_07098_));
 DFF_X1 \data_out_real[83]$_SDFFE_PN0P_  (.D(_00298_),
    .CK(clknet_leaf_54_clk),
    .Q(net352),
    .QN(_07097_));
 DFF_X1 \data_out_real[84]$_SDFFE_PN0P_  (.D(_00299_),
    .CK(clknet_leaf_54_clk),
    .Q(net353),
    .QN(_07096_));
 DFF_X1 \data_out_real[85]$_SDFFE_PN0P_  (.D(_00300_),
    .CK(clknet_leaf_62_clk),
    .Q(net354),
    .QN(_07095_));
 DFF_X1 \data_out_real[86]$_SDFFE_PN0P_  (.D(_00301_),
    .CK(clknet_leaf_63_clk),
    .Q(net355),
    .QN(_07094_));
 DFF_X1 \data_out_real[87]$_SDFFE_PN0P_  (.D(_00302_),
    .CK(clknet_leaf_63_clk),
    .Q(net356),
    .QN(_07093_));
 DFF_X1 \data_out_real[88]$_SDFFE_PN0P_  (.D(_00303_),
    .CK(clknet_leaf_66_clk),
    .Q(net357),
    .QN(_07092_));
 DFF_X2 \data_out_real[89]$_SDFFE_PN0P_  (.D(_00304_),
    .CK(clknet_leaf_67_clk),
    .Q(net358),
    .QN(_07091_));
 DFF_X2 \data_out_real[8]$_SDFFE_PN0P_  (.D(_00305_),
    .CK(clknet_leaf_68_clk),
    .Q(net359),
    .QN(_07090_));
 DFF_X2 \data_out_real[90]$_SDFFE_PN0P_  (.D(_00306_),
    .CK(clknet_leaf_67_clk),
    .Q(net360),
    .QN(_07089_));
 DFF_X1 \data_out_real[91]$_SDFFE_PN0P_  (.D(_00307_),
    .CK(clknet_leaf_65_clk),
    .Q(net361),
    .QN(_07088_));
 DFF_X2 \data_out_real[92]$_SDFFE_PN0P_  (.D(_00308_),
    .CK(clknet_leaf_65_clk),
    .Q(net362),
    .QN(_07087_));
 DFF_X2 \data_out_real[93]$_SDFFE_PN0P_  (.D(_00309_),
    .CK(clknet_leaf_68_clk),
    .Q(net363),
    .QN(_07086_));
 DFF_X2 \data_out_real[94]$_SDFFE_PN0P_  (.D(_00310_),
    .CK(clknet_leaf_76_clk),
    .Q(net364),
    .QN(_07085_));
 DFF_X2 \data_out_real[95]$_SDFFE_PN0P_  (.D(_00311_),
    .CK(clknet_leaf_74_clk),
    .Q(net365),
    .QN(_07084_));
 DFF_X2 \data_out_real[96]$_SDFFE_PN0P_  (.D(_00312_),
    .CK(clknet_leaf_76_clk),
    .Q(net366),
    .QN(_07083_));
 DFF_X2 \data_out_real[97]$_SDFFE_PN0P_  (.D(_00313_),
    .CK(clknet_leaf_76_clk),
    .Q(net367),
    .QN(_07082_));
 DFF_X2 \data_out_real[98]$_SDFFE_PN0P_  (.D(_00314_),
    .CK(clknet_leaf_75_clk),
    .Q(net368),
    .QN(_07081_));
 DFF_X2 \data_out_real[99]$_SDFFE_PN0P_  (.D(_00315_),
    .CK(clknet_leaf_76_clk),
    .Q(net369),
    .QN(_07080_));
 DFF_X2 \data_out_real[9]$_SDFFE_PN0P_  (.D(_00316_),
    .CK(clknet_leaf_79_clk),
    .Q(net370),
    .QN(_07079_));
 DFF_X2 \data_ready$_SDFFE_PN1P_  (.D(_00317_),
    .CK(clknet_leaf_79_clk),
    .Q(net371),
    .QN(_07078_));
 DFF_X2 \data_valid_out$_SDFFE_PN0P_  (.D(_00318_),
    .CK(clknet_leaf_1_clk),
    .Q(net372),
    .QN(_07077_));
 DFF_X1 \group[0]$_DFFE_PP_  (.D(_00319_),
    .CK(clknet_leaf_77_clk),
    .Q(\group[0] ),
    .QN(_07076_));
 DFF_X1 \group[1]$_DFFE_PP_  (.D(_00320_),
    .CK(clknet_leaf_77_clk),
    .Q(\group[1] ),
    .QN(_07075_));
 DFF_X1 \group[2]$_DFFE_PP_  (.D(_00321_),
    .CK(clknet_leaf_77_clk),
    .Q(\group[2] ),
    .QN(_07074_));
 DFF_X1 \idx1[0]$_DFFE_PP_  (.D(_00013_),
    .CK(clknet_leaf_74_clk),
    .Q(\idx1[0] ),
    .QN(_00038_));
 DFF_X1 \idx1[1]$_DFFE_PP_  (.D(_00014_),
    .CK(clknet_leaf_79_clk),
    .Q(\idx1[1] ),
    .QN(_00026_));
 DFF_X1 \idx1[2]$_DFFE_PP_  (.D(_00015_),
    .CK(clknet_leaf_74_clk),
    .Q(\idx1[2] ),
    .QN(_00028_));
 DFF_X1 \idx2[0]$_DFFE_PP_  (.D(_00016_),
    .CK(clknet_leaf_36_clk),
    .Q(\idx2[0] ),
    .QN(_00030_));
 DFF_X2 \idx2[1]$_DFFE_PP_  (.D(_00017_),
    .CK(clknet_leaf_37_clk),
    .Q(\idx2[1] ),
    .QN(_07073_));
 DFF_X1 \idx2[2]$_DFFE_PP_  (.D(_00018_),
    .CK(clknet_leaf_37_clk),
    .Q(\idx2[2] ),
    .QN(_07072_));
 DFF_X1 \sample_count[0]$_SDFFE_PN0P_  (.D(_00322_),
    .CK(clknet_leaf_2_clk),
    .Q(\sample_count[0] ),
    .QN(_09376_));
 DFF_X1 \sample_count[1]$_SDFFE_PN0P_  (.D(_00323_),
    .CK(clknet_leaf_2_clk),
    .Q(\sample_count[1] ),
    .QN(_09377_));
 DFF_X1 \sample_count[2]$_SDFFE_PN0P_  (.D(_00324_),
    .CK(clknet_leaf_2_clk),
    .Q(\sample_count[2] ),
    .QN(_07071_));
 DFF_X2 \samples_imag[0][0]$_DFFE_PP_  (.D(_00325_),
    .CK(clknet_leaf_3_clk),
    .Q(\samples_imag[0][0] ),
    .QN(_07070_));
 DFF_X2 \samples_imag[0][10]$_DFFE_PP_  (.D(_00326_),
    .CK(clknet_leaf_6_clk),
    .Q(\samples_imag[0][10] ),
    .QN(_07069_));
 DFF_X2 \samples_imag[0][11]$_DFFE_PP_  (.D(_00327_),
    .CK(clknet_leaf_7_clk),
    .Q(\samples_imag[0][11] ),
    .QN(_07068_));
 DFF_X2 \samples_imag[0][12]$_DFFE_PP_  (.D(_00328_),
    .CK(clknet_leaf_6_clk),
    .Q(\samples_imag[0][12] ),
    .QN(_07067_));
 DFF_X2 \samples_imag[0][13]$_DFFE_PP_  (.D(_00329_),
    .CK(clknet_leaf_6_clk),
    .Q(\samples_imag[0][13] ),
    .QN(_07066_));
 DFF_X2 \samples_imag[0][14]$_DFFE_PP_  (.D(_00330_),
    .CK(clknet_leaf_4_clk),
    .Q(\samples_imag[0][14] ),
    .QN(_07065_));
 DFF_X2 \samples_imag[0][15]$_DFFE_PP_  (.D(_00331_),
    .CK(clknet_leaf_3_clk),
    .Q(\samples_imag[0][15] ),
    .QN(_07064_));
 DFF_X2 \samples_imag[0][1]$_DFFE_PP_  (.D(_00332_),
    .CK(clknet_leaf_4_clk),
    .Q(\samples_imag[0][1] ),
    .QN(_07063_));
 DFF_X2 \samples_imag[0][2]$_DFFE_PP_  (.D(_00333_),
    .CK(clknet_leaf_37_clk),
    .Q(\samples_imag[0][2] ),
    .QN(_07062_));
 DFF_X2 \samples_imag[0][3]$_DFFE_PP_  (.D(_00334_),
    .CK(clknet_leaf_3_clk),
    .Q(\samples_imag[0][3] ),
    .QN(_07061_));
 DFF_X2 \samples_imag[0][4]$_DFFE_PP_  (.D(_00335_),
    .CK(clknet_leaf_4_clk),
    .Q(\samples_imag[0][4] ),
    .QN(_07060_));
 DFF_X2 \samples_imag[0][5]$_DFFE_PP_  (.D(_00336_),
    .CK(clknet_leaf_4_clk),
    .Q(\samples_imag[0][5] ),
    .QN(_07059_));
 DFF_X2 \samples_imag[0][6]$_DFFE_PP_  (.D(_00337_),
    .CK(clknet_leaf_5_clk),
    .Q(\samples_imag[0][6] ),
    .QN(_07058_));
 DFF_X2 \samples_imag[0][7]$_DFFE_PP_  (.D(_00338_),
    .CK(clknet_leaf_5_clk),
    .Q(\samples_imag[0][7] ),
    .QN(_07057_));
 DFF_X2 \samples_imag[0][8]$_DFFE_PP_  (.D(_00339_),
    .CK(clknet_leaf_5_clk),
    .Q(\samples_imag[0][8] ),
    .QN(_07056_));
 DFF_X1 \samples_imag[0][9]$_DFFE_PP_  (.D(_00340_),
    .CK(clknet_leaf_6_clk),
    .Q(\samples_imag[0][9] ),
    .QN(_07055_));
 DFF_X1 \samples_imag[1][0]$_DFFE_PP_  (.D(_00341_),
    .CK(clknet_leaf_30_clk),
    .Q(\samples_imag[1][0] ),
    .QN(_07054_));
 DFF_X1 \samples_imag[1][10]$_DFFE_PP_  (.D(_00342_),
    .CK(clknet_leaf_19_clk),
    .Q(\samples_imag[1][10] ),
    .QN(_07053_));
 DFF_X1 \samples_imag[1][11]$_DFFE_PP_  (.D(_00343_),
    .CK(clknet_leaf_19_clk),
    .Q(\samples_imag[1][11] ),
    .QN(_07052_));
 DFF_X1 \samples_imag[1][12]$_DFFE_PP_  (.D(_00344_),
    .CK(clknet_leaf_23_clk),
    .Q(\samples_imag[1][12] ),
    .QN(_07051_));
 DFF_X1 \samples_imag[1][13]$_DFFE_PP_  (.D(_00345_),
    .CK(clknet_leaf_23_clk),
    .Q(\samples_imag[1][13] ),
    .QN(_07050_));
 DFF_X1 \samples_imag[1][14]$_DFFE_PP_  (.D(_00346_),
    .CK(clknet_leaf_26_clk),
    .Q(\samples_imag[1][14] ),
    .QN(_07049_));
 DFF_X2 \samples_imag[1][15]$_DFFE_PP_  (.D(_00347_),
    .CK(clknet_leaf_33_clk),
    .Q(\samples_imag[1][15] ),
    .QN(_07048_));
 DFF_X1 \samples_imag[1][1]$_DFFE_PP_  (.D(_00348_),
    .CK(clknet_leaf_25_clk),
    .Q(\samples_imag[1][1] ),
    .QN(_07047_));
 DFF_X1 \samples_imag[1][2]$_DFFE_PP_  (.D(_00349_),
    .CK(clknet_leaf_33_clk),
    .Q(\samples_imag[1][2] ),
    .QN(_07046_));
 DFF_X1 \samples_imag[1][3]$_DFFE_PP_  (.D(_00350_),
    .CK(clknet_leaf_34_clk),
    .Q(\samples_imag[1][3] ),
    .QN(_07045_));
 DFF_X1 \samples_imag[1][4]$_DFFE_PP_  (.D(_00351_),
    .CK(clknet_leaf_34_clk),
    .Q(\samples_imag[1][4] ),
    .QN(_07044_));
 DFF_X1 \samples_imag[1][5]$_DFFE_PP_  (.D(_00352_),
    .CK(clknet_leaf_25_clk),
    .Q(\samples_imag[1][5] ),
    .QN(_07043_));
 DFF_X2 \samples_imag[1][6]$_DFFE_PP_  (.D(_00353_),
    .CK(clknet_leaf_25_clk),
    .Q(\samples_imag[1][6] ),
    .QN(_07042_));
 DFF_X1 \samples_imag[1][7]$_DFFE_PP_  (.D(_00354_),
    .CK(clknet_leaf_22_clk),
    .Q(\samples_imag[1][7] ),
    .QN(_07041_));
 DFF_X1 \samples_imag[1][8]$_DFFE_PP_  (.D(_00355_),
    .CK(clknet_leaf_23_clk),
    .Q(\samples_imag[1][8] ),
    .QN(_07040_));
 DFF_X1 \samples_imag[1][9]$_DFFE_PP_  (.D(_00356_),
    .CK(clknet_leaf_23_clk),
    .Q(\samples_imag[1][9] ),
    .QN(_07039_));
 DFF_X2 \samples_imag[2][0]$_DFFE_PP_  (.D(_00357_),
    .CK(clknet_leaf_26_clk),
    .Q(\samples_imag[2][0] ),
    .QN(_07038_));
 DFF_X1 \samples_imag[2][10]$_DFFE_PP_  (.D(_00358_),
    .CK(clknet_leaf_23_clk),
    .Q(\samples_imag[2][10] ),
    .QN(_07037_));
 DFF_X1 \samples_imag[2][11]$_DFFE_PP_  (.D(_00359_),
    .CK(clknet_leaf_23_clk),
    .Q(\samples_imag[2][11] ),
    .QN(_07036_));
 DFF_X1 \samples_imag[2][12]$_DFFE_PP_  (.D(_00360_),
    .CK(clknet_leaf_23_clk),
    .Q(\samples_imag[2][12] ),
    .QN(_07035_));
 DFF_X1 \samples_imag[2][13]$_DFFE_PP_  (.D(_00361_),
    .CK(clknet_leaf_22_clk),
    .Q(\samples_imag[2][13] ),
    .QN(_07034_));
 DFF_X2 \samples_imag[2][14]$_DFFE_PP_  (.D(_00362_),
    .CK(clknet_leaf_22_clk),
    .Q(\samples_imag[2][14] ),
    .QN(_07033_));
 DFF_X2 \samples_imag[2][15]$_DFFE_PP_  (.D(_00363_),
    .CK(clknet_leaf_34_clk),
    .Q(\samples_imag[2][15] ),
    .QN(_07032_));
 DFF_X2 \samples_imag[2][1]$_DFFE_PP_  (.D(_00364_),
    .CK(clknet_leaf_26_clk),
    .Q(\samples_imag[2][1] ),
    .QN(_07031_));
 DFF_X2 \samples_imag[2][2]$_DFFE_PP_  (.D(_00365_),
    .CK(clknet_leaf_34_clk),
    .Q(\samples_imag[2][2] ),
    .QN(_07030_));
 DFF_X2 \samples_imag[2][3]$_DFFE_PP_  (.D(_00366_),
    .CK(clknet_leaf_34_clk),
    .Q(\samples_imag[2][3] ),
    .QN(_07029_));
 DFF_X2 \samples_imag[2][4]$_DFFE_PP_  (.D(_00367_),
    .CK(clknet_leaf_34_clk),
    .Q(\samples_imag[2][4] ),
    .QN(_07028_));
 DFF_X1 \samples_imag[2][5]$_DFFE_PP_  (.D(_00368_),
    .CK(clknet_leaf_26_clk),
    .Q(\samples_imag[2][5] ),
    .QN(_07027_));
 DFF_X2 \samples_imag[2][6]$_DFFE_PP_  (.D(_00369_),
    .CK(clknet_leaf_25_clk),
    .Q(\samples_imag[2][6] ),
    .QN(_07026_));
 DFF_X2 \samples_imag[2][7]$_DFFE_PP_  (.D(_00370_),
    .CK(clknet_leaf_22_clk),
    .Q(\samples_imag[2][7] ),
    .QN(_07025_));
 DFF_X1 \samples_imag[2][8]$_DFFE_PP_  (.D(_00371_),
    .CK(clknet_leaf_24_clk),
    .Q(\samples_imag[2][8] ),
    .QN(_07024_));
 DFF_X1 \samples_imag[2][9]$_DFFE_PP_  (.D(_00372_),
    .CK(clknet_leaf_24_clk),
    .Q(\samples_imag[2][9] ),
    .QN(_07023_));
 DFF_X1 \samples_imag[3][0]$_DFFE_PP_  (.D(_00373_),
    .CK(clknet_leaf_30_clk),
    .Q(\samples_imag[3][0] ),
    .QN(_07022_));
 DFF_X1 \samples_imag[3][10]$_DFFE_PP_  (.D(_00374_),
    .CK(clknet_leaf_23_clk),
    .Q(\samples_imag[3][10] ),
    .QN(_07021_));
 DFF_X1 \samples_imag[3][11]$_DFFE_PP_  (.D(_00375_),
    .CK(clknet_leaf_18_clk),
    .Q(\samples_imag[3][11] ),
    .QN(_07020_));
 DFF_X1 \samples_imag[3][12]$_DFFE_PP_  (.D(_00376_),
    .CK(clknet_leaf_15_clk),
    .Q(\samples_imag[3][12] ),
    .QN(_07019_));
 DFF_X1 \samples_imag[3][13]$_DFFE_PP_  (.D(_00377_),
    .CK(clknet_leaf_15_clk),
    .Q(\samples_imag[3][13] ),
    .QN(_07018_));
 DFF_X2 \samples_imag[3][14]$_DFFE_PP_  (.D(_00378_),
    .CK(clknet_leaf_18_clk),
    .Q(\samples_imag[3][14] ),
    .QN(_07017_));
 DFF_X2 \samples_imag[3][15]$_DFFE_PP_  (.D(_00379_),
    .CK(clknet_leaf_33_clk),
    .Q(\samples_imag[3][15] ),
    .QN(_07016_));
 DFF_X1 \samples_imag[3][1]$_DFFE_PP_  (.D(_00380_),
    .CK(clknet_leaf_26_clk),
    .Q(\samples_imag[3][1] ),
    .QN(_07015_));
 DFF_X2 \samples_imag[3][2]$_DFFE_PP_  (.D(_00381_),
    .CK(clknet_leaf_33_clk),
    .Q(\samples_imag[3][2] ),
    .QN(_07014_));
 DFF_X1 \samples_imag[3][3]$_DFFE_PP_  (.D(_00382_),
    .CK(clknet_leaf_34_clk),
    .Q(\samples_imag[3][3] ),
    .QN(_07013_));
 DFF_X1 \samples_imag[3][4]$_DFFE_PP_  (.D(_00383_),
    .CK(clknet_leaf_25_clk),
    .Q(\samples_imag[3][4] ),
    .QN(_07012_));
 DFF_X1 \samples_imag[3][5]$_DFFE_PP_  (.D(_00384_),
    .CK(clknet_leaf_26_clk),
    .Q(\samples_imag[3][5] ),
    .QN(_07011_));
 DFF_X2 \samples_imag[3][6]$_DFFE_PP_  (.D(_00385_),
    .CK(clknet_leaf_25_clk),
    .Q(\samples_imag[3][6] ),
    .QN(_07010_));
 DFF_X1 \samples_imag[3][7]$_DFFE_PP_  (.D(_00386_),
    .CK(clknet_leaf_24_clk),
    .Q(\samples_imag[3][7] ),
    .QN(_07009_));
 DFF_X1 \samples_imag[3][8]$_DFFE_PP_  (.D(_00387_),
    .CK(clknet_leaf_24_clk),
    .Q(\samples_imag[3][8] ),
    .QN(_07008_));
 DFF_X1 \samples_imag[3][9]$_DFFE_PP_  (.D(_00388_),
    .CK(clknet_leaf_24_clk),
    .Q(\samples_imag[3][9] ),
    .QN(_07007_));
 DFF_X2 \samples_imag[4][0]$_DFFE_PP_  (.D(_00389_),
    .CK(clknet_leaf_15_clk),
    .Q(\samples_imag[4][0] ),
    .QN(_07006_));
 DFF_X1 \samples_imag[4][10]$_DFFE_PP_  (.D(_00390_),
    .CK(clknet_leaf_13_clk),
    .Q(\samples_imag[4][10] ),
    .QN(_07005_));
 DFF_X1 \samples_imag[4][11]$_DFFE_PP_  (.D(_00391_),
    .CK(clknet_leaf_13_clk),
    .Q(\samples_imag[4][11] ),
    .QN(_07004_));
 DFF_X1 \samples_imag[4][12]$_DFFE_PP_  (.D(_00392_),
    .CK(clknet_leaf_13_clk),
    .Q(\samples_imag[4][12] ),
    .QN(_07003_));
 DFF_X1 \samples_imag[4][13]$_DFFE_PP_  (.D(_00393_),
    .CK(clknet_leaf_12_clk),
    .Q(\samples_imag[4][13] ),
    .QN(_07002_));
 DFF_X2 \samples_imag[4][14]$_DFFE_PP_  (.D(_00394_),
    .CK(clknet_leaf_15_clk),
    .Q(\samples_imag[4][14] ),
    .QN(_07001_));
 DFF_X2 \samples_imag[4][15]$_DFFE_PP_  (.D(_00395_),
    .CK(clknet_leaf_35_clk),
    .Q(\samples_imag[4][15] ),
    .QN(_07000_));
 DFF_X2 \samples_imag[4][1]$_DFFE_PP_  (.D(_00396_),
    .CK(clknet_leaf_15_clk),
    .Q(\samples_imag[4][1] ),
    .QN(_06999_));
 DFF_X2 \samples_imag[4][2]$_DFFE_PP_  (.D(_00397_),
    .CK(clknet_leaf_35_clk),
    .Q(\samples_imag[4][2] ),
    .QN(_06998_));
 DFF_X2 \samples_imag[4][3]$_DFFE_PP_  (.D(_00398_),
    .CK(clknet_leaf_35_clk),
    .Q(\samples_imag[4][3] ),
    .QN(_06997_));
 DFF_X2 \samples_imag[4][4]$_DFFE_PP_  (.D(_00399_),
    .CK(clknet_leaf_13_clk),
    .Q(\samples_imag[4][4] ),
    .QN(_06996_));
 DFF_X2 \samples_imag[4][5]$_DFFE_PP_  (.D(_00400_),
    .CK(clknet_leaf_13_clk),
    .Q(\samples_imag[4][5] ),
    .QN(_06995_));
 DFF_X1 \samples_imag[4][6]$_DFFE_PP_  (.D(_00401_),
    .CK(clknet_leaf_13_clk),
    .Q(\samples_imag[4][6] ),
    .QN(_06994_));
 DFF_X1 \samples_imag[4][7]$_DFFE_PP_  (.D(_00402_),
    .CK(clknet_leaf_5_clk),
    .Q(\samples_imag[4][7] ),
    .QN(_06993_));
 DFF_X1 \samples_imag[4][8]$_DFFE_PP_  (.D(_00403_),
    .CK(clknet_leaf_5_clk),
    .Q(\samples_imag[4][8] ),
    .QN(_06992_));
 DFF_X1 \samples_imag[4][9]$_DFFE_PP_  (.D(_00404_),
    .CK(clknet_leaf_5_clk),
    .Q(\samples_imag[4][9] ),
    .QN(_06991_));
 DFF_X2 \samples_imag[5][0]$_DFFE_PP_  (.D(_00405_),
    .CK(clknet_leaf_14_clk),
    .Q(\samples_imag[5][0] ),
    .QN(_06990_));
 DFF_X1 \samples_imag[5][10]$_DFFE_PP_  (.D(_00406_),
    .CK(clknet_leaf_14_clk),
    .Q(\samples_imag[5][10] ),
    .QN(_06989_));
 DFF_X1 \samples_imag[5][11]$_DFFE_PP_  (.D(_00407_),
    .CK(clknet_leaf_15_clk),
    .Q(\samples_imag[5][11] ),
    .QN(_06988_));
 DFF_X1 \samples_imag[5][12]$_DFFE_PP_  (.D(_00408_),
    .CK(clknet_leaf_16_clk),
    .Q(\samples_imag[5][12] ),
    .QN(_06987_));
 DFF_X1 \samples_imag[5][13]$_DFFE_PP_  (.D(_00409_),
    .CK(clknet_leaf_15_clk),
    .Q(\samples_imag[5][13] ),
    .QN(_06986_));
 DFF_X1 \samples_imag[5][14]$_DFFE_PP_  (.D(_00410_),
    .CK(clknet_leaf_15_clk),
    .Q(\samples_imag[5][14] ),
    .QN(_06985_));
 DFF_X1 \samples_imag[5][15]$_DFFE_PP_  (.D(_00411_),
    .CK(clknet_leaf_35_clk),
    .Q(\samples_imag[5][15] ),
    .QN(_06984_));
 DFF_X1 \samples_imag[5][1]$_DFFE_PP_  (.D(_00412_),
    .CK(clknet_leaf_12_clk),
    .Q(\samples_imag[5][1] ),
    .QN(_06983_));
 DFF_X2 \samples_imag[5][2]$_DFFE_PP_  (.D(_00413_),
    .CK(clknet_leaf_35_clk),
    .Q(\samples_imag[5][2] ),
    .QN(_06982_));
 DFF_X2 \samples_imag[5][3]$_DFFE_PP_  (.D(_00414_),
    .CK(clknet_leaf_35_clk),
    .Q(\samples_imag[5][3] ),
    .QN(_06981_));
 DFF_X2 \samples_imag[5][4]$_DFFE_PP_  (.D(_00415_),
    .CK(clknet_leaf_14_clk),
    .Q(\samples_imag[5][4] ),
    .QN(_06980_));
 DFF_X2 \samples_imag[5][5]$_DFFE_PP_  (.D(_00416_),
    .CK(clknet_leaf_14_clk),
    .Q(\samples_imag[5][5] ),
    .QN(_06979_));
 DFF_X1 \samples_imag[5][6]$_DFFE_PP_  (.D(_00417_),
    .CK(clknet_leaf_12_clk),
    .Q(\samples_imag[5][6] ),
    .QN(_06978_));
 DFF_X2 \samples_imag[5][7]$_DFFE_PP_  (.D(_00418_),
    .CK(clknet_leaf_14_clk),
    .Q(\samples_imag[5][7] ),
    .QN(_06977_));
 DFF_X2 \samples_imag[5][8]$_DFFE_PP_  (.D(_00419_),
    .CK(clknet_leaf_14_clk),
    .Q(\samples_imag[5][8] ),
    .QN(_06976_));
 DFF_X2 \samples_imag[5][9]$_DFFE_PP_  (.D(_00420_),
    .CK(clknet_leaf_14_clk),
    .Q(\samples_imag[5][9] ),
    .QN(_06975_));
 DFF_X1 \samples_imag[6][0]$_DFFE_PP_  (.D(_00421_),
    .CK(clknet_leaf_5_clk),
    .Q(\samples_imag[6][0] ),
    .QN(_06974_));
 DFF_X2 \samples_imag[6][10]$_DFFE_PP_  (.D(_00422_),
    .CK(clknet_leaf_82_clk),
    .Q(\samples_imag[6][10] ),
    .QN(_06973_));
 DFF_X2 \samples_imag[6][11]$_DFFE_PP_  (.D(_00423_),
    .CK(clknet_leaf_7_clk),
    .Q(\samples_imag[6][11] ),
    .QN(_06972_));
 DFF_X2 \samples_imag[6][12]$_DFFE_PP_  (.D(_00424_),
    .CK(clknet_leaf_8_clk),
    .Q(\samples_imag[6][12] ),
    .QN(_06971_));
 DFF_X2 \samples_imag[6][13]$_DFFE_PP_  (.D(_00425_),
    .CK(clknet_leaf_7_clk),
    .Q(\samples_imag[6][13] ),
    .QN(_06970_));
 DFF_X2 \samples_imag[6][14]$_DFFE_PP_  (.D(_00426_),
    .CK(clknet_leaf_7_clk),
    .Q(\samples_imag[6][14] ),
    .QN(_06969_));
 DFF_X2 \samples_imag[6][15]$_DFFE_PP_  (.D(_00427_),
    .CK(clknet_leaf_36_clk),
    .Q(\samples_imag[6][15] ),
    .QN(_06968_));
 DFF_X2 \samples_imag[6][1]$_DFFE_PP_  (.D(_00428_),
    .CK(clknet_leaf_6_clk),
    .Q(\samples_imag[6][1] ),
    .QN(_06967_));
 DFF_X1 \samples_imag[6][2]$_DFFE_PP_  (.D(_00429_),
    .CK(clknet_leaf_36_clk),
    .Q(\samples_imag[6][2] ),
    .QN(_06966_));
 DFF_X1 \samples_imag[6][3]$_DFFE_PP_  (.D(_00430_),
    .CK(clknet_leaf_4_clk),
    .Q(\samples_imag[6][3] ),
    .QN(_06965_));
 DFF_X2 \samples_imag[6][4]$_DFFE_PP_  (.D(_00431_),
    .CK(clknet_leaf_3_clk),
    .Q(\samples_imag[6][4] ),
    .QN(_06964_));
 DFF_X2 \samples_imag[6][5]$_DFFE_PP_  (.D(_00432_),
    .CK(clknet_leaf_3_clk),
    .Q(\samples_imag[6][5] ),
    .QN(_06963_));
 DFF_X2 \samples_imag[6][6]$_DFFE_PP_  (.D(_00433_),
    .CK(clknet_leaf_82_clk),
    .Q(\samples_imag[6][6] ),
    .QN(_06962_));
 DFF_X2 \samples_imag[6][7]$_DFFE_PP_  (.D(_00434_),
    .CK(clknet_leaf_82_clk),
    .Q(\samples_imag[6][7] ),
    .QN(_06961_));
 DFF_X2 \samples_imag[6][8]$_DFFE_PP_  (.D(_00435_),
    .CK(clknet_leaf_82_clk),
    .Q(\samples_imag[6][8] ),
    .QN(_06960_));
 DFF_X2 \samples_imag[6][9]$_DFFE_PP_  (.D(_00436_),
    .CK(clknet_leaf_82_clk),
    .Q(\samples_imag[6][9] ),
    .QN(_06959_));
 DFF_X2 \samples_imag[7][0]$_DFFE_PP_  (.D(_00437_),
    .CK(clknet_leaf_7_clk),
    .Q(\samples_imag[7][0] ),
    .QN(_06958_));
 DFF_X1 \samples_imag[7][10]$_DFFE_PP_  (.D(_00438_),
    .CK(clknet_leaf_7_clk),
    .Q(\samples_imag[7][10] ),
    .QN(_06957_));
 DFF_X2 \samples_imag[7][11]$_DFFE_PP_  (.D(_00439_),
    .CK(clknet_leaf_8_clk),
    .Q(\samples_imag[7][11] ),
    .QN(_06956_));
 DFF_X2 \samples_imag[7][12]$_DFFE_PP_  (.D(_00440_),
    .CK(clknet_leaf_8_clk),
    .Q(\samples_imag[7][12] ),
    .QN(_06955_));
 DFF_X2 \samples_imag[7][13]$_DFFE_PP_  (.D(_00441_),
    .CK(clknet_leaf_8_clk),
    .Q(\samples_imag[7][13] ),
    .QN(_06954_));
 DFF_X2 \samples_imag[7][14]$_DFFE_PP_  (.D(_00442_),
    .CK(clknet_leaf_10_clk),
    .Q(\samples_imag[7][14] ),
    .QN(_06953_));
 DFF_X2 \samples_imag[7][15]$_DFFE_PP_  (.D(_00443_),
    .CK(clknet_leaf_36_clk),
    .Q(\samples_imag[7][15] ),
    .QN(_06952_));
 DFF_X2 \samples_imag[7][1]$_DFFE_PP_  (.D(_00444_),
    .CK(clknet_leaf_7_clk),
    .Q(\samples_imag[7][1] ),
    .QN(_06951_));
 DFF_X2 \samples_imag[7][2]$_DFFE_PP_  (.D(_00445_),
    .CK(clknet_leaf_36_clk),
    .Q(\samples_imag[7][2] ),
    .QN(_06950_));
 DFF_X2 \samples_imag[7][3]$_DFFE_PP_  (.D(_00446_),
    .CK(clknet_leaf_4_clk),
    .Q(\samples_imag[7][3] ),
    .QN(_06949_));
 DFF_X2 \samples_imag[7][4]$_DFFE_PP_  (.D(_00447_),
    .CK(clknet_leaf_4_clk),
    .Q(\samples_imag[7][4] ),
    .QN(_06948_));
 DFF_X2 \samples_imag[7][5]$_DFFE_PP_  (.D(_00448_),
    .CK(clknet_leaf_4_clk),
    .Q(\samples_imag[7][5] ),
    .QN(_06947_));
 DFF_X2 \samples_imag[7][6]$_DFFE_PP_  (.D(_00449_),
    .CK(clknet_leaf_8_clk),
    .Q(\samples_imag[7][6] ),
    .QN(_06946_));
 DFF_X2 \samples_imag[7][7]$_DFFE_PP_  (.D(_00450_),
    .CK(clknet_leaf_82_clk),
    .Q(\samples_imag[7][7] ),
    .QN(_06945_));
 DFF_X2 \samples_imag[7][8]$_DFFE_PP_  (.D(_00451_),
    .CK(clknet_leaf_82_clk),
    .Q(\samples_imag[7][8] ),
    .QN(_06944_));
 DFF_X2 \samples_imag[7][9]$_DFFE_PP_  (.D(_00452_),
    .CK(clknet_leaf_6_clk),
    .Q(\samples_imag[7][9] ),
    .QN(_06943_));
 DFF_X1 \samples_real[0][0]$_DFFE_PP_  (.D(_00453_),
    .CK(clknet_leaf_40_clk),
    .Q(\samples_real[0][0] ),
    .QN(_06942_));
 DFF_X2 \samples_real[0][10]$_DFFE_PP_  (.D(_00454_),
    .CK(clknet_leaf_72_clk),
    .Q(\samples_real[0][10] ),
    .QN(_06941_));
 DFF_X2 \samples_real[0][11]$_DFFE_PP_  (.D(_00455_),
    .CK(clknet_leaf_71_clk),
    .Q(\samples_real[0][11] ),
    .QN(_06940_));
 DFF_X2 \samples_real[0][12]$_DFFE_PP_  (.D(_00456_),
    .CK(clknet_leaf_70_clk),
    .Q(\samples_real[0][12] ),
    .QN(_06939_));
 DFF_X2 \samples_real[0][13]$_DFFE_PP_  (.D(_00457_),
    .CK(clknet_leaf_69_clk),
    .Q(\samples_real[0][13] ),
    .QN(_06938_));
 DFF_X2 \samples_real[0][14]$_DFFE_PP_  (.D(_00458_),
    .CK(clknet_leaf_70_clk),
    .Q(\samples_real[0][14] ),
    .QN(_06937_));
 DFF_X2 \samples_real[0][15]$_DFFE_PP_  (.D(_00459_),
    .CK(clknet_leaf_37_clk),
    .Q(\samples_real[0][15] ),
    .QN(_06936_));
 DFF_X2 \samples_real[0][1]$_DFFE_PP_  (.D(_00460_),
    .CK(clknet_leaf_71_clk),
    .Q(\samples_real[0][1] ),
    .QN(_06935_));
 DFF_X2 \samples_real[0][2]$_DFFE_PP_  (.D(_00461_),
    .CK(clknet_leaf_38_clk),
    .Q(\samples_real[0][2] ),
    .QN(_06934_));
 DFF_X2 \samples_real[0][3]$_DFFE_PP_  (.D(_00462_),
    .CK(clknet_leaf_72_clk),
    .Q(\samples_real[0][3] ),
    .QN(_06933_));
 DFF_X2 \samples_real[0][4]$_DFFE_PP_  (.D(_00463_),
    .CK(clknet_leaf_38_clk),
    .Q(\samples_real[0][4] ),
    .QN(_06932_));
 DFF_X2 \samples_real[0][5]$_DFFE_PP_  (.D(_00464_),
    .CK(clknet_leaf_73_clk),
    .Q(\samples_real[0][5] ),
    .QN(_06931_));
 DFF_X2 \samples_real[0][6]$_DFFE_PP_  (.D(_00465_),
    .CK(clknet_leaf_38_clk),
    .Q(\samples_real[0][6] ),
    .QN(_06930_));
 DFF_X2 \samples_real[0][7]$_DFFE_PP_  (.D(_00466_),
    .CK(clknet_leaf_38_clk),
    .Q(\samples_real[0][7] ),
    .QN(_06929_));
 DFF_X2 \samples_real[0][8]$_DFFE_PP_  (.D(_00467_),
    .CK(clknet_leaf_73_clk),
    .Q(\samples_real[0][8] ),
    .QN(_06928_));
 DFF_X2 \samples_real[0][9]$_DFFE_PP_  (.D(_00468_),
    .CK(clknet_leaf_37_clk),
    .Q(\samples_real[0][9] ),
    .QN(_06927_));
 DFF_X1 \samples_real[1][0]$_DFFE_PP_  (.D(_00469_),
    .CK(clknet_leaf_50_clk),
    .Q(\samples_real[1][0] ),
    .QN(_06926_));
 DFF_X1 \samples_real[1][10]$_DFFE_PP_  (.D(_00470_),
    .CK(clknet_leaf_43_clk),
    .Q(\samples_real[1][10] ),
    .QN(_06925_));
 DFF_X1 \samples_real[1][11]$_DFFE_PP_  (.D(_00471_),
    .CK(clknet_leaf_51_clk),
    .Q(\samples_real[1][11] ),
    .QN(_06924_));
 DFF_X1 \samples_real[1][12]$_DFFE_PP_  (.D(_00472_),
    .CK(clknet_leaf_50_clk),
    .Q(\samples_real[1][12] ),
    .QN(_06923_));
 DFF_X2 \samples_real[1][13]$_DFFE_PP_  (.D(_00473_),
    .CK(clknet_leaf_52_clk),
    .Q(\samples_real[1][13] ),
    .QN(_06922_));
 DFF_X1 \samples_real[1][14]$_DFFE_PP_  (.D(_00474_),
    .CK(clknet_leaf_52_clk),
    .Q(\samples_real[1][14] ),
    .QN(_06921_));
 DFF_X1 \samples_real[1][15]$_DFFE_PP_  (.D(_00475_),
    .CK(clknet_leaf_33_clk),
    .Q(\samples_real[1][15] ),
    .QN(_06920_));
 DFF_X1 \samples_real[1][1]$_DFFE_PP_  (.D(_00476_),
    .CK(clknet_leaf_51_clk),
    .Q(\samples_real[1][1] ),
    .QN(_06919_));
 DFF_X2 \samples_real[1][2]$_DFFE_PP_  (.D(_00477_),
    .CK(clknet_leaf_42_clk),
    .Q(\samples_real[1][2] ),
    .QN(_06918_));
 DFF_X1 \samples_real[1][3]$_DFFE_PP_  (.D(_00478_),
    .CK(clknet_leaf_51_clk),
    .Q(\samples_real[1][3] ),
    .QN(_06917_));
 DFF_X1 \samples_real[1][4]$_DFFE_PP_  (.D(_00479_),
    .CK(clknet_leaf_47_clk),
    .Q(\samples_real[1][4] ),
    .QN(_06916_));
 DFF_X1 \samples_real[1][5]$_DFFE_PP_  (.D(_00480_),
    .CK(clknet_leaf_50_clk),
    .Q(\samples_real[1][5] ),
    .QN(_06915_));
 DFF_X1 \samples_real[1][6]$_DFFE_PP_  (.D(_00481_),
    .CK(clknet_leaf_44_clk),
    .Q(\samples_real[1][6] ),
    .QN(_06914_));
 DFF_X1 \samples_real[1][7]$_DFFE_PP_  (.D(_00482_),
    .CK(clknet_leaf_42_clk),
    .Q(\samples_real[1][7] ),
    .QN(_06913_));
 DFF_X1 \samples_real[1][8]$_DFFE_PP_  (.D(_00483_),
    .CK(clknet_leaf_44_clk),
    .Q(\samples_real[1][8] ),
    .QN(_06912_));
 DFF_X1 \samples_real[1][9]$_DFFE_PP_  (.D(_00484_),
    .CK(clknet_leaf_44_clk),
    .Q(\samples_real[1][9] ),
    .QN(_06911_));
 DFF_X1 \samples_real[2][0]$_DFFE_PP_  (.D(_00485_),
    .CK(clknet_leaf_41_clk),
    .Q(\samples_real[2][0] ),
    .QN(_06910_));
 DFF_X1 \samples_real[2][10]$_DFFE_PP_  (.D(_00486_),
    .CK(clknet_leaf_41_clk),
    .Q(\samples_real[2][10] ),
    .QN(_06909_));
 DFF_X1 \samples_real[2][11]$_DFFE_PP_  (.D(_00487_),
    .CK(clknet_leaf_52_clk),
    .Q(\samples_real[2][11] ),
    .QN(_06908_));
 DFF_X1 \samples_real[2][12]$_DFFE_PP_  (.D(_00488_),
    .CK(clknet_leaf_52_clk),
    .Q(\samples_real[2][12] ),
    .QN(_06907_));
 DFF_X1 \samples_real[2][13]$_DFFE_PP_  (.D(_00489_),
    .CK(clknet_leaf_52_clk),
    .Q(\samples_real[2][13] ),
    .QN(_06906_));
 DFF_X1 \samples_real[2][14]$_DFFE_PP_  (.D(_00490_),
    .CK(clknet_leaf_52_clk),
    .Q(\samples_real[2][14] ),
    .QN(_06905_));
 DFF_X1 \samples_real[2][15]$_DFFE_PP_  (.D(_00491_),
    .CK(clknet_leaf_32_clk),
    .Q(\samples_real[2][15] ),
    .QN(_06904_));
 DFF_X1 \samples_real[2][1]$_DFFE_PP_  (.D(_00492_),
    .CK(clknet_leaf_51_clk),
    .Q(\samples_real[2][1] ),
    .QN(_06903_));
 DFF_X1 \samples_real[2][2]$_DFFE_PP_  (.D(_00493_),
    .CK(clknet_leaf_42_clk),
    .Q(\samples_real[2][2] ),
    .QN(_06902_));
 DFF_X1 \samples_real[2][3]$_DFFE_PP_  (.D(_00494_),
    .CK(clknet_leaf_41_clk),
    .Q(\samples_real[2][3] ),
    .QN(_06901_));
 DFF_X1 \samples_real[2][4]$_DFFE_PP_  (.D(_00495_),
    .CK(clknet_leaf_41_clk),
    .Q(\samples_real[2][4] ),
    .QN(_06900_));
 DFF_X1 \samples_real[2][5]$_DFFE_PP_  (.D(_00496_),
    .CK(clknet_leaf_41_clk),
    .Q(\samples_real[2][5] ),
    .QN(_06899_));
 DFF_X1 \samples_real[2][6]$_DFFE_PP_  (.D(_00497_),
    .CK(clknet_leaf_33_clk),
    .Q(\samples_real[2][6] ),
    .QN(_06898_));
 DFF_X1 \samples_real[2][7]$_DFFE_PP_  (.D(_00498_),
    .CK(clknet_leaf_43_clk),
    .Q(\samples_real[2][7] ),
    .QN(_06897_));
 DFF_X2 \samples_real[2][8]$_DFFE_PP_  (.D(_00499_),
    .CK(clknet_leaf_43_clk),
    .Q(\samples_real[2][8] ),
    .QN(_06896_));
 DFF_X1 \samples_real[2][9]$_DFFE_PP_  (.D(_00500_),
    .CK(clknet_leaf_44_clk),
    .Q(\samples_real[2][9] ),
    .QN(_06895_));
 DFF_X1 \samples_real[3][0]$_DFFE_PP_  (.D(_00501_),
    .CK(clknet_leaf_47_clk),
    .Q(\samples_real[3][0] ),
    .QN(_06894_));
 DFF_X2 \samples_real[3][10]$_DFFE_PP_  (.D(_00502_),
    .CK(clknet_leaf_43_clk),
    .Q(\samples_real[3][10] ),
    .QN(_06893_));
 DFF_X2 \samples_real[3][11]$_DFFE_PP_  (.D(_00503_),
    .CK(clknet_leaf_53_clk),
    .Q(\samples_real[3][11] ),
    .QN(_06892_));
 DFF_X2 \samples_real[3][12]$_DFFE_PP_  (.D(_00504_),
    .CK(clknet_leaf_53_clk),
    .Q(\samples_real[3][12] ),
    .QN(_06891_));
 DFF_X1 \samples_real[3][13]$_DFFE_PP_  (.D(_00505_),
    .CK(clknet_leaf_53_clk),
    .Q(\samples_real[3][13] ),
    .QN(_06890_));
 DFF_X2 \samples_real[3][14]$_DFFE_PP_  (.D(_00506_),
    .CK(clknet_leaf_53_clk),
    .Q(\samples_real[3][14] ),
    .QN(_06889_));
 DFF_X2 \samples_real[3][15]$_DFFE_PP_  (.D(_00507_),
    .CK(clknet_leaf_42_clk),
    .Q(\samples_real[3][15] ),
    .QN(_06888_));
 DFF_X1 \samples_real[3][1]$_DFFE_PP_  (.D(_00508_),
    .CK(clknet_leaf_51_clk),
    .Q(\samples_real[3][1] ),
    .QN(_06887_));
 DFF_X1 \samples_real[3][2]$_DFFE_PP_  (.D(_00509_),
    .CK(clknet_leaf_42_clk),
    .Q(\samples_real[3][2] ),
    .QN(_06886_));
 DFF_X1 \samples_real[3][3]$_DFFE_PP_  (.D(_00510_),
    .CK(clknet_leaf_51_clk),
    .Q(\samples_real[3][3] ),
    .QN(_06885_));
 DFF_X1 \samples_real[3][4]$_DFFE_PP_  (.D(_00511_),
    .CK(clknet_leaf_41_clk),
    .Q(\samples_real[3][4] ),
    .QN(_06884_));
 DFF_X1 \samples_real[3][5]$_DFFE_PP_  (.D(_00512_),
    .CK(clknet_leaf_51_clk),
    .Q(\samples_real[3][5] ),
    .QN(_06883_));
 DFF_X1 \samples_real[3][6]$_DFFE_PP_  (.D(_00513_),
    .CK(clknet_leaf_43_clk),
    .Q(\samples_real[3][6] ),
    .QN(_06882_));
 DFF_X1 \samples_real[3][7]$_DFFE_PP_  (.D(_00514_),
    .CK(clknet_leaf_43_clk),
    .Q(\samples_real[3][7] ),
    .QN(_06881_));
 DFF_X1 \samples_real[3][8]$_DFFE_PP_  (.D(_00515_),
    .CK(clknet_leaf_43_clk),
    .Q(\samples_real[3][8] ),
    .QN(_06880_));
 DFF_X1 \samples_real[3][9]$_DFFE_PP_  (.D(_00516_),
    .CK(clknet_leaf_44_clk),
    .Q(\samples_real[3][9] ),
    .QN(_06879_));
 DFF_X2 \samples_real[4][0]$_DFFE_PP_  (.D(_00517_),
    .CK(clknet_leaf_53_clk),
    .Q(\samples_real[4][0] ),
    .QN(_06878_));
 DFF_X2 \samples_real[4][10]$_DFFE_PP_  (.D(_00518_),
    .CK(clknet_leaf_53_clk),
    .Q(\samples_real[4][10] ),
    .QN(_06877_));
 DFF_X1 \samples_real[4][11]$_DFFE_PP_  (.D(_00519_),
    .CK(clknet_leaf_63_clk),
    .Q(\samples_real[4][11] ),
    .QN(_06876_));
 DFF_X1 \samples_real[4][12]$_DFFE_PP_  (.D(_00520_),
    .CK(clknet_leaf_63_clk),
    .Q(\samples_real[4][12] ),
    .QN(_06875_));
 DFF_X1 \samples_real[4][13]$_DFFE_PP_  (.D(_00521_),
    .CK(clknet_leaf_52_clk),
    .Q(\samples_real[4][13] ),
    .QN(_06874_));
 DFF_X1 \samples_real[4][14]$_DFFE_PP_  (.D(_00522_),
    .CK(clknet_leaf_63_clk),
    .Q(\samples_real[4][14] ),
    .QN(_06873_));
 DFF_X2 \samples_real[4][15]$_DFFE_PP_  (.D(_00523_),
    .CK(clknet_leaf_39_clk),
    .Q(\samples_real[4][15] ),
    .QN(_06872_));
 DFF_X2 \samples_real[4][1]$_DFFE_PP_  (.D(_00524_),
    .CK(clknet_leaf_64_clk),
    .Q(\samples_real[4][1] ),
    .QN(_06871_));
 DFF_X2 \samples_real[4][2]$_DFFE_PP_  (.D(_00525_),
    .CK(clknet_leaf_39_clk),
    .Q(\samples_real[4][2] ),
    .QN(_06870_));
 DFF_X2 \samples_real[4][3]$_DFFE_PP_  (.D(_00526_),
    .CK(clknet_leaf_52_clk),
    .Q(\samples_real[4][3] ),
    .QN(_06869_));
 DFF_X2 \samples_real[4][4]$_DFFE_PP_  (.D(_00527_),
    .CK(clknet_leaf_64_clk),
    .Q(\samples_real[4][4] ),
    .QN(_06868_));
 DFF_X1 \samples_real[4][5]$_DFFE_PP_  (.D(_00528_),
    .CK(clknet_leaf_63_clk),
    .Q(\samples_real[4][5] ),
    .QN(_06867_));
 DFF_X2 \samples_real[4][6]$_DFFE_PP_  (.D(_00529_),
    .CK(clknet_leaf_41_clk),
    .Q(\samples_real[4][6] ),
    .QN(_06866_));
 DFF_X2 \samples_real[4][7]$_DFFE_PP_  (.D(_00530_),
    .CK(clknet_leaf_40_clk),
    .Q(\samples_real[4][7] ),
    .QN(_06865_));
 DFF_X2 \samples_real[4][8]$_DFFE_PP_  (.D(_00531_),
    .CK(clknet_leaf_39_clk),
    .Q(\samples_real[4][8] ),
    .QN(_06864_));
 DFF_X2 \samples_real[4][9]$_DFFE_PP_  (.D(_00532_),
    .CK(clknet_leaf_40_clk),
    .Q(\samples_real[4][9] ),
    .QN(_06863_));
 DFF_X2 \samples_real[5][0]$_DFFE_PP_  (.D(_00533_),
    .CK(clknet_leaf_70_clk),
    .Q(\samples_real[5][0] ),
    .QN(_06862_));
 DFF_X2 \samples_real[5][10]$_DFFE_PP_  (.D(_00534_),
    .CK(clknet_leaf_69_clk),
    .Q(\samples_real[5][10] ),
    .QN(_06861_));
 DFF_X1 \samples_real[5][11]$_DFFE_PP_  (.D(_00535_),
    .CK(clknet_leaf_65_clk),
    .Q(\samples_real[5][11] ),
    .QN(_06860_));
 DFF_X1 \samples_real[5][12]$_DFFE_PP_  (.D(_00536_),
    .CK(clknet_leaf_65_clk),
    .Q(\samples_real[5][12] ),
    .QN(_06859_));
 DFF_X2 \samples_real[5][13]$_DFFE_PP_  (.D(_00537_),
    .CK(clknet_leaf_69_clk),
    .Q(\samples_real[5][13] ),
    .QN(_06858_));
 DFF_X1 \samples_real[5][14]$_DFFE_PP_  (.D(_00538_),
    .CK(clknet_leaf_69_clk),
    .Q(\samples_real[5][14] ),
    .QN(_06857_));
 DFF_X2 \samples_real[5][15]$_DFFE_PP_  (.D(_00539_),
    .CK(clknet_leaf_38_clk),
    .Q(\samples_real[5][15] ),
    .QN(_06856_));
 DFF_X2 \samples_real[5][1]$_DFFE_PP_  (.D(_00540_),
    .CK(clknet_leaf_65_clk),
    .Q(\samples_real[5][1] ),
    .QN(_06855_));
 DFF_X2 \samples_real[5][2]$_DFFE_PP_  (.D(_00541_),
    .CK(clknet_leaf_39_clk),
    .Q(\samples_real[5][2] ),
    .QN(_06854_));
 DFF_X2 \samples_real[5][3]$_DFFE_PP_  (.D(_00542_),
    .CK(clknet_leaf_70_clk),
    .Q(\samples_real[5][3] ),
    .QN(_06853_));
 DFF_X2 \samples_real[5][4]$_DFFE_PP_  (.D(_00543_),
    .CK(clknet_leaf_70_clk),
    .Q(\samples_real[5][4] ),
    .QN(_06852_));
 DFF_X1 \samples_real[5][5]$_DFFE_PP_  (.D(_00544_),
    .CK(clknet_leaf_65_clk),
    .Q(\samples_real[5][5] ),
    .QN(_06851_));
 DFF_X2 \samples_real[5][6]$_DFFE_PP_  (.D(_00545_),
    .CK(clknet_leaf_71_clk),
    .Q(\samples_real[5][6] ),
    .QN(_06850_));
 DFF_X2 \samples_real[5][7]$_DFFE_PP_  (.D(_00546_),
    .CK(clknet_leaf_70_clk),
    .Q(\samples_real[5][7] ),
    .QN(_06849_));
 DFF_X2 \samples_real[5][8]$_DFFE_PP_  (.D(_00547_),
    .CK(clknet_leaf_40_clk),
    .Q(\samples_real[5][8] ),
    .QN(_06848_));
 DFF_X2 \samples_real[5][9]$_DFFE_PP_  (.D(_00548_),
    .CK(clknet_leaf_72_clk),
    .Q(\samples_real[5][9] ),
    .QN(_06847_));
 DFF_X2 \samples_real[6][0]$_DFFE_PP_  (.D(_00549_),
    .CK(clknet_leaf_68_clk),
    .Q(\samples_real[6][0] ),
    .QN(_06846_));
 DFF_X2 \samples_real[6][10]$_DFFE_PP_  (.D(_00550_),
    .CK(clknet_leaf_69_clk),
    .Q(\samples_real[6][10] ),
    .QN(_06845_));
 DFF_X2 \samples_real[6][11]$_DFFE_PP_  (.D(_00551_),
    .CK(clknet_leaf_67_clk),
    .Q(\samples_real[6][11] ),
    .QN(_06844_));
 DFF_X2 \samples_real[6][12]$_DFFE_PP_  (.D(_00552_),
    .CK(clknet_leaf_68_clk),
    .Q(\samples_real[6][12] ),
    .QN(_06843_));
 DFF_X2 \samples_real[6][13]$_DFFE_PP_  (.D(_00553_),
    .CK(clknet_leaf_69_clk),
    .Q(\samples_real[6][13] ),
    .QN(_06842_));
 DFF_X2 \samples_real[6][14]$_DFFE_PP_  (.D(_00554_),
    .CK(clknet_leaf_69_clk),
    .Q(\samples_real[6][14] ),
    .QN(_06841_));
 DFF_X2 \samples_real[6][15]$_DFFE_PP_  (.D(_00555_),
    .CK(clknet_leaf_38_clk),
    .Q(\samples_real[6][15] ),
    .QN(_06840_));
 DFF_X2 \samples_real[6][1]$_DFFE_PP_  (.D(_00556_),
    .CK(clknet_leaf_68_clk),
    .Q(\samples_real[6][1] ),
    .QN(_06839_));
 DFF_X2 \samples_real[6][2]$_DFFE_PP_  (.D(_00557_),
    .CK(clknet_leaf_38_clk),
    .Q(\samples_real[6][2] ),
    .QN(_06838_));
 DFF_X2 \samples_real[6][3]$_DFFE_PP_  (.D(_00558_),
    .CK(clknet_leaf_68_clk),
    .Q(\samples_real[6][3] ),
    .QN(_06837_));
 DFF_X2 \samples_real[6][4]$_DFFE_PP_  (.D(_00559_),
    .CK(clknet_leaf_69_clk),
    .Q(\samples_real[6][4] ),
    .QN(_06836_));
 DFF_X2 \samples_real[6][5]$_DFFE_PP_  (.D(_00560_),
    .CK(clknet_leaf_68_clk),
    .Q(\samples_real[6][5] ),
    .QN(_06835_));
 DFF_X2 \samples_real[6][6]$_DFFE_PP_  (.D(_00561_),
    .CK(clknet_leaf_73_clk),
    .Q(\samples_real[6][6] ),
    .QN(_06834_));
 DFF_X2 \samples_real[6][7]$_DFFE_PP_  (.D(_00562_),
    .CK(clknet_leaf_73_clk),
    .Q(\samples_real[6][7] ),
    .QN(_06833_));
 DFF_X2 \samples_real[6][8]$_DFFE_PP_  (.D(_00563_),
    .CK(clknet_leaf_72_clk),
    .Q(\samples_real[6][8] ),
    .QN(_06832_));
 DFF_X2 \samples_real[6][9]$_DFFE_PP_  (.D(_00564_),
    .CK(clknet_leaf_72_clk),
    .Q(\samples_real[6][9] ),
    .QN(_06831_));
 DFF_X2 \samples_real[7][0]$_DFFE_PP_  (.D(_00565_),
    .CK(clknet_leaf_70_clk),
    .Q(\samples_real[7][0] ),
    .QN(_06830_));
 DFF_X2 \samples_real[7][10]$_DFFE_PP_  (.D(_00566_),
    .CK(clknet_leaf_71_clk),
    .Q(\samples_real[7][10] ),
    .QN(_06829_));
 DFF_X2 \samples_real[7][11]$_DFFE_PP_  (.D(_00567_),
    .CK(clknet_leaf_66_clk),
    .Q(\samples_real[7][11] ),
    .QN(_06828_));
 DFF_X2 \samples_real[7][12]$_DFFE_PP_  (.D(_00568_),
    .CK(clknet_leaf_66_clk),
    .Q(\samples_real[7][12] ),
    .QN(_06827_));
 DFF_X2 \samples_real[7][13]$_DFFE_PP_  (.D(_00569_),
    .CK(clknet_leaf_71_clk),
    .Q(\samples_real[7][13] ),
    .QN(_06826_));
 DFF_X2 \samples_real[7][14]$_DFFE_PP_  (.D(_00570_),
    .CK(clknet_leaf_64_clk),
    .Q(\samples_real[7][14] ),
    .QN(_06825_));
 DFF_X2 \samples_real[7][15]$_DFFE_PP_  (.D(_00571_),
    .CK(clknet_leaf_39_clk),
    .Q(\samples_real[7][15] ),
    .QN(_06824_));
 DFF_X2 \samples_real[7][1]$_DFFE_PP_  (.D(_00572_),
    .CK(clknet_leaf_64_clk),
    .Q(\samples_real[7][1] ),
    .QN(_06823_));
 DFF_X2 \samples_real[7][2]$_DFFE_PP_  (.D(_00573_),
    .CK(clknet_leaf_39_clk),
    .Q(\samples_real[7][2] ),
    .QN(_06822_));
 DFF_X1 \samples_real[7][3]$_DFFE_PP_  (.D(_00574_),
    .CK(clknet_leaf_64_clk),
    .Q(\samples_real[7][3] ),
    .QN(_06821_));
 DFF_X1 \samples_real[7][4]$_DFFE_PP_  (.D(_00575_),
    .CK(clknet_leaf_64_clk),
    .Q(\samples_real[7][4] ),
    .QN(_06820_));
 DFF_X1 \samples_real[7][5]$_DFFE_PP_  (.D(_00576_),
    .CK(clknet_leaf_66_clk),
    .Q(\samples_real[7][5] ),
    .QN(_06819_));
 DFF_X2 \samples_real[7][6]$_DFFE_PP_  (.D(_00577_),
    .CK(clknet_leaf_71_clk),
    .Q(\samples_real[7][6] ),
    .QN(_06818_));
 DFF_X2 \samples_real[7][7]$_DFFE_PP_  (.D(_00578_),
    .CK(clknet_leaf_71_clk),
    .Q(\samples_real[7][7] ),
    .QN(_06817_));
 DFF_X2 \samples_real[7][8]$_DFFE_PP_  (.D(_00579_),
    .CK(clknet_leaf_40_clk),
    .Q(\samples_real[7][8] ),
    .QN(_06816_));
 DFF_X2 \samples_real[7][9]$_DFFE_PP_  (.D(_00580_),
    .CK(clknet_leaf_72_clk),
    .Q(\samples_real[7][9] ),
    .QN(_06815_));
 DFF_X2 \stage[0]$_SDFFE_PN0P_  (.D(_00581_),
    .CK(clknet_leaf_78_clk),
    .Q(\stage[0] ),
    .QN(_09361_));
 DFF_X2 \stage[1]$_SDFFE_PN0P_  (.D(_00582_),
    .CK(clknet_leaf_78_clk),
    .Q(\stage[1] ),
    .QN(_09362_));
 DFF_X2 \stage[2]$_SDFFE_PN0P_  (.D(_00583_),
    .CK(clknet_leaf_78_clk),
    .Q(\stage[2] ),
    .QN(_09340_));
 DFF_X1 \state[0]$_DFF_P_  (.D(_00010_),
    .CK(clknet_leaf_1_clk),
    .Q(\state[0] ),
    .QN(_07346_));
 DFF_X1 \state[1]$_DFF_P_  (.D(_00011_),
    .CK(clknet_leaf_79_clk),
    .Q(\state[1] ),
    .QN(_00031_));
 DFF_X1 \state[2]$_DFF_P_  (.D(_00012_),
    .CK(clknet_leaf_79_clk),
    .Q(\state[2] ),
    .QN(_00020_));
 DFF_X1 \state[3]$_DFF_P_  (.D(_00009_),
    .CK(clknet_leaf_79_clk),
    .Q(\state[3] ),
    .QN(_00041_));
 DFF_X2 \temp_imag[0]$_DFFE_PP_  (.D(_00584_),
    .CK(clknet_leaf_1_clk),
    .Q(\temp_imag[0] ),
    .QN(_07347_));
 DFF_X2 \temp_real[0]$_DFFE_PP_  (.D(_00585_),
    .CK(clknet_leaf_75_clk),
    .Q(\temp_real[0] ),
    .QN(_07355_));
 DFF_X1 \twiddle_idx[0]$_DFFE_PP_  (.D(_00006_),
    .CK(clknet_leaf_75_clk),
    .Q(\twiddle_idx[0] ),
    .QN(_06814_));
 DFF_X1 \twiddle_idx[1]$_DFFE_PP_  (.D(_00019_),
    .CK(clknet_leaf_75_clk),
    .Q(\twiddle_idx[1] ),
    .QN(_06813_));
 NOR4_X4 clone1 (.A1(_03748_),
    .A2(_03723_),
    .A3(_03736_),
    .A4(_03680_),
    .ZN(net1));
 NAND3_X4 clone2 (.A1(_02196_),
    .A2(_02259_),
    .A3(_02232_),
    .ZN(net2));
 BUF_X4 clone14 (.A(_03990_),
    .Z(net14));
 NOR3_X4 clone15 (.A1(_02116_),
    .A2(_02097_),
    .A3(_02120_),
    .ZN(net15));
 BUF_X4 clone17 (.A(_02278_),
    .Z(net17));
 BUF_X4 clone18 (.A(_02641_),
    .Z(net18));
 BUF_X2 clone19 (.A(_02334_),
    .Z(net19));
 NAND2_X2 clone20 (.A1(net21),
    .A2(_03501_),
    .ZN(net20));
 AND3_X1 clone21 (.A1(net403),
    .A2(_03412_),
    .A3(_03473_),
    .ZN(net21));
 BUF_X4 clone23 (.A(_03789_),
    .Z(net23));
 BUF_X4 clone24 (.A(_04723_),
    .Z(net24));
 BUF_X4 clone25 (.A(_01300_),
    .Z(net25));
 BUF_X4 clone26 (.A(_04356_),
    .Z(net26));
 NAND4_X4 clone27 (.A1(_02697_),
    .A2(_02685_),
    .A3(net380),
    .A4(_02731_),
    .ZN(net27));
 BUF_X4 clone28 (.A(_02016_),
    .Z(net28));
 BUF_X4 clone29 (.A(_02132_),
    .Z(net29));
 BUF_X2 clone31 (.A(_09309_),
    .Z(net31));
 BUF_X4 clone32 (.A(_03351_),
    .Z(net32));
 BUF_X8 clone34 (.A(net411),
    .Z(net34));
 BUF_X4 clone35 (.A(_02523_),
    .Z(net35));
 BUF_X4 clone36 (.A(_01308_),
    .Z(net36));
 NAND2_X4 clone37 (.A1(net429),
    .A2(_04521_),
    .ZN(net37));
 BUF_X4 clone38 (.A(_03502_),
    .Z(net38));
 BUF_X4 clone39 (.A(_03112_),
    .Z(net39));
 BUF_X4 clone40 (.A(_04134_),
    .Z(net40));
 BUF_X4 clone41 (.A(_03051_),
    .Z(net41));
 NAND2_X4 clone42 (.A1(_01082_),
    .A2(_01081_),
    .ZN(net42));
 BUF_X1 split43 (.A(_08828_),
    .Z(net43));
 BUF_X4 clone44 (.A(_04724_),
    .Z(net44));
 BUF_X4 clone51 (.A(_00004_),
    .Z(net51));
 BUF_X4 clone53 (.A(_04869_),
    .Z(net53));
 BUF_X1 split61 (.A(_00001_),
    .Z(net61));
 BUF_X16 clone93 (.A(_06119_),
    .Z(net93));
 BUF_X8 clone101 (.A(_06146_),
    .Z(net101));
 BUF_X16 clone104 (.A(_06173_),
    .Z(net104));
 BUF_X16 clone107 (.A(_06200_),
    .Z(net107));
 BUF_X16 clone130 (.A(net458),
    .Z(net130));
 BUF_X16 clone131 (.A(_05761_),
    .Z(net131));
 MUX2_X2 clone138 (.A(_05358_),
    .B(_05341_),
    .S(_05418_),
    .Z(net138));
 BUF_X4 clone139 (.A(_05421_),
    .Z(net139));
 BUF_X4 clone140 (.A(_05424_),
    .Z(net140));
 BUF_X2 clone143 (.A(_05789_),
    .Z(net143));
 BUF_X4 clone144 (.A(net534),
    .Z(net144));
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Right_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Right_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Right_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Right_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Right_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Right_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Right_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Right_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Right_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Right_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Right_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Right_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Right_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Right_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Right_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Right_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Right_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Right_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Right_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Right_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Right_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Right_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Right_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Right_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Right_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Right_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Left_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Left_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Left_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Left_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Left_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Left_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Left_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Left_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Left_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Left_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Left_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Left_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Left_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Left_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Left_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Left_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Left_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Left_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Left_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Left_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Left_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Left_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Left_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Left_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Left_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Left_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Left_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Left_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Left_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Left_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Left_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Left_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Left_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Left_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Left_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Left_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Left_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Left_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Left_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Left_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Left_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Left_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Left_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Left_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Left_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Left_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Left_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Left_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Left_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Left_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Left_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Left_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Left_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Left_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Left_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Left_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Left_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Left_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Left_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Left_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Left_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Left_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Left_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Left_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Left_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Left_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Left_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Left_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Left_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Left_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Left_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Left_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Left_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Left_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Left_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Left_265 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_266 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_267 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_268 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_269 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_270 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_271 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_272 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_273 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_274 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_275 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_276 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_277 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_278 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_279 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_280 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_281 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_282 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_283 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_284 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_285 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_286 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_287 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_288 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_289 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_290 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_291 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_292 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_293 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_294 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_295 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_296 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_297 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_298 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_299 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_300 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_301 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_302 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_303 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_304 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_305 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_306 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_307 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_308 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_309 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_310 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_311 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_312 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_313 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_314 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_315 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_316 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_317 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_318 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_319 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_320 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_321 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_322 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_323 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_324 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_325 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_326 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_327 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_328 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_329 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_330 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_331 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_332 ();
 BUF_X2 input1 (.A(data_in_imag[0]),
    .Z(net45));
 CLKBUF_X2 input2 (.A(data_in_imag[10]),
    .Z(net46));
 CLKBUF_X2 input3 (.A(data_in_imag[11]),
    .Z(net47));
 CLKBUF_X2 input4 (.A(data_in_imag[12]),
    .Z(net48));
 CLKBUF_X2 input5 (.A(data_in_imag[13]),
    .Z(net49));
 BUF_X2 input6 (.A(data_in_imag[14]),
    .Z(net50));
 BUF_X1 input7 (.A(data_in_imag[15]),
    .Z(net54));
 BUF_X2 input8 (.A(data_in_imag[1]),
    .Z(net55));
 BUF_X2 input9 (.A(data_in_imag[2]),
    .Z(net62));
 BUF_X2 input10 (.A(data_in_imag[3]),
    .Z(net63));
 BUF_X2 input11 (.A(data_in_imag[4]),
    .Z(net64));
 BUF_X2 input12 (.A(data_in_imag[5]),
    .Z(net65));
 BUF_X2 input13 (.A(data_in_imag[6]),
    .Z(net66));
 BUF_X2 input14 (.A(data_in_imag[7]),
    .Z(net67));
 BUF_X2 input15 (.A(data_in_imag[8]),
    .Z(net68));
 CLKBUF_X2 input16 (.A(data_in_imag[9]),
    .Z(net69));
 BUF_X2 input17 (.A(data_in_real[0]),
    .Z(net70));
 BUF_X2 input18 (.A(data_in_real[10]),
    .Z(net71));
 BUF_X2 input19 (.A(data_in_real[11]),
    .Z(net72));
 BUF_X2 input20 (.A(data_in_real[12]),
    .Z(net73));
 BUF_X2 input21 (.A(data_in_real[13]),
    .Z(net74));
 BUF_X2 input22 (.A(data_in_real[14]),
    .Z(net75));
 CLKBUF_X2 input23 (.A(data_in_real[15]),
    .Z(net76));
 BUF_X2 input24 (.A(data_in_real[1]),
    .Z(net77));
 BUF_X2 input25 (.A(data_in_real[2]),
    .Z(net78));
 BUF_X2 input26 (.A(data_in_real[3]),
    .Z(net79));
 BUF_X2 input27 (.A(data_in_real[4]),
    .Z(net80));
 BUF_X2 input28 (.A(data_in_real[5]),
    .Z(net81));
 BUF_X2 input29 (.A(data_in_real[6]),
    .Z(net82));
 BUF_X2 input30 (.A(data_in_real[7]),
    .Z(net83));
 BUF_X2 input31 (.A(data_in_real[8]),
    .Z(net84));
 BUF_X2 input32 (.A(data_in_real[9]),
    .Z(net85));
 BUF_X2 input33 (.A(data_valid_in),
    .Z(net86));
 BUF_X2 input34 (.A(start),
    .Z(net87));
 BUF_X1 output35 (.A(net88),
    .Z(busy));
 BUF_X1 output36 (.A(net89),
    .Z(data_out_imag[0]));
 BUF_X1 output37 (.A(net90),
    .Z(data_out_imag[100]));
 BUF_X1 output38 (.A(net91),
    .Z(data_out_imag[101]));
 BUF_X1 output39 (.A(net92),
    .Z(data_out_imag[102]));
 BUF_X1 output40 (.A(net95),
    .Z(data_out_imag[103]));
 BUF_X1 output41 (.A(net96),
    .Z(data_out_imag[104]));
 BUF_X1 output42 (.A(net99),
    .Z(data_out_imag[105]));
 BUF_X1 output43 (.A(net100),
    .Z(data_out_imag[106]));
 BUF_X1 output44 (.A(net102),
    .Z(data_out_imag[107]));
 BUF_X1 output45 (.A(net103),
    .Z(data_out_imag[108]));
 BUF_X1 output46 (.A(net105),
    .Z(data_out_imag[109]));
 BUF_X1 output47 (.A(net106),
    .Z(data_out_imag[10]));
 BUF_X1 output48 (.A(net108),
    .Z(data_out_imag[110]));
 BUF_X1 output49 (.A(net109),
    .Z(data_out_imag[111]));
 BUF_X1 output50 (.A(net110),
    .Z(data_out_imag[112]));
 BUF_X1 output51 (.A(net111),
    .Z(data_out_imag[113]));
 BUF_X1 output52 (.A(net112),
    .Z(data_out_imag[114]));
 BUF_X1 output53 (.A(net113),
    .Z(data_out_imag[115]));
 BUF_X1 output54 (.A(net114),
    .Z(data_out_imag[116]));
 BUF_X1 output55 (.A(net115),
    .Z(data_out_imag[117]));
 BUF_X1 output56 (.A(net116),
    .Z(data_out_imag[118]));
 BUF_X1 output57 (.A(net117),
    .Z(data_out_imag[119]));
 BUF_X1 output58 (.A(net118),
    .Z(data_out_imag[11]));
 BUF_X1 output59 (.A(net119),
    .Z(data_out_imag[120]));
 BUF_X1 output60 (.A(net120),
    .Z(data_out_imag[121]));
 BUF_X1 output61 (.A(net121),
    .Z(data_out_imag[122]));
 BUF_X1 output62 (.A(net122),
    .Z(data_out_imag[123]));
 BUF_X1 output63 (.A(net123),
    .Z(data_out_imag[124]));
 BUF_X1 output64 (.A(net124),
    .Z(data_out_imag[125]));
 BUF_X1 output65 (.A(net126),
    .Z(data_out_imag[126]));
 BUF_X1 output66 (.A(net127),
    .Z(data_out_imag[127]));
 BUF_X1 output67 (.A(net128),
    .Z(data_out_imag[12]));
 BUF_X1 output68 (.A(net134),
    .Z(data_out_imag[13]));
 BUF_X1 output69 (.A(net135),
    .Z(data_out_imag[14]));
 BUF_X1 output70 (.A(net136),
    .Z(data_out_imag[15]));
 BUF_X1 output71 (.A(net141),
    .Z(data_out_imag[16]));
 BUF_X1 output72 (.A(net142),
    .Z(data_out_imag[17]));
 BUF_X1 output73 (.A(net145),
    .Z(data_out_imag[18]));
 BUF_X1 output74 (.A(net146),
    .Z(data_out_imag[19]));
 BUF_X1 output75 (.A(net147),
    .Z(data_out_imag[1]));
 BUF_X1 output76 (.A(net148),
    .Z(data_out_imag[20]));
 BUF_X1 output77 (.A(net150),
    .Z(data_out_imag[21]));
 BUF_X1 output78 (.A(net155),
    .Z(data_out_imag[22]));
 BUF_X1 output79 (.A(net157),
    .Z(data_out_imag[23]));
 BUF_X1 output80 (.A(net159),
    .Z(data_out_imag[24]));
 BUF_X1 output81 (.A(net160),
    .Z(data_out_imag[25]));
 BUF_X1 output82 (.A(net161),
    .Z(data_out_imag[26]));
 BUF_X1 output83 (.A(net162),
    .Z(data_out_imag[27]));
 BUF_X1 output84 (.A(net163),
    .Z(data_out_imag[28]));
 BUF_X1 output85 (.A(net164),
    .Z(data_out_imag[29]));
 BUF_X1 output86 (.A(net165),
    .Z(data_out_imag[2]));
 BUF_X1 output87 (.A(net166),
    .Z(data_out_imag[30]));
 BUF_X1 output88 (.A(net167),
    .Z(data_out_imag[31]));
 BUF_X1 output89 (.A(net168),
    .Z(data_out_imag[32]));
 BUF_X1 output90 (.A(net169),
    .Z(data_out_imag[33]));
 BUF_X1 output91 (.A(net170),
    .Z(data_out_imag[34]));
 BUF_X1 output92 (.A(net171),
    .Z(data_out_imag[35]));
 BUF_X1 output93 (.A(net172),
    .Z(data_out_imag[36]));
 BUF_X1 output94 (.A(net173),
    .Z(data_out_imag[37]));
 BUF_X1 output95 (.A(net174),
    .Z(data_out_imag[38]));
 BUF_X1 output96 (.A(net175),
    .Z(data_out_imag[39]));
 BUF_X1 output97 (.A(net176),
    .Z(data_out_imag[3]));
 BUF_X1 output98 (.A(net177),
    .Z(data_out_imag[40]));
 BUF_X1 output99 (.A(net178),
    .Z(data_out_imag[41]));
 BUF_X1 output100 (.A(net179),
    .Z(data_out_imag[42]));
 BUF_X1 output101 (.A(net180),
    .Z(data_out_imag[43]));
 BUF_X1 output102 (.A(net181),
    .Z(data_out_imag[44]));
 BUF_X1 output103 (.A(net182),
    .Z(data_out_imag[45]));
 BUF_X1 output104 (.A(net183),
    .Z(data_out_imag[46]));
 BUF_X1 output105 (.A(net184),
    .Z(data_out_imag[47]));
 BUF_X1 output106 (.A(net185),
    .Z(data_out_imag[48]));
 BUF_X1 output107 (.A(net186),
    .Z(data_out_imag[49]));
 BUF_X1 output108 (.A(net187),
    .Z(data_out_imag[4]));
 BUF_X1 output109 (.A(net188),
    .Z(data_out_imag[50]));
 BUF_X1 output110 (.A(net189),
    .Z(data_out_imag[51]));
 BUF_X1 output111 (.A(net190),
    .Z(data_out_imag[52]));
 BUF_X1 output112 (.A(net191),
    .Z(data_out_imag[53]));
 BUF_X1 output113 (.A(net192),
    .Z(data_out_imag[54]));
 BUF_X1 output114 (.A(net193),
    .Z(data_out_imag[55]));
 BUF_X1 output115 (.A(net194),
    .Z(data_out_imag[56]));
 BUF_X1 output116 (.A(net195),
    .Z(data_out_imag[57]));
 BUF_X1 output117 (.A(net196),
    .Z(data_out_imag[58]));
 BUF_X1 output118 (.A(net197),
    .Z(data_out_imag[59]));
 BUF_X1 output119 (.A(net198),
    .Z(data_out_imag[5]));
 BUF_X1 output120 (.A(net199),
    .Z(data_out_imag[60]));
 BUF_X1 output121 (.A(net200),
    .Z(data_out_imag[61]));
 BUF_X1 output122 (.A(net201),
    .Z(data_out_imag[62]));
 BUF_X1 output123 (.A(net202),
    .Z(data_out_imag[63]));
 BUF_X1 output124 (.A(net203),
    .Z(data_out_imag[64]));
 BUF_X1 output125 (.A(net204),
    .Z(data_out_imag[65]));
 BUF_X1 output126 (.A(net205),
    .Z(data_out_imag[66]));
 BUF_X1 output127 (.A(net206),
    .Z(data_out_imag[67]));
 BUF_X1 output128 (.A(net207),
    .Z(data_out_imag[68]));
 BUF_X1 output129 (.A(net208),
    .Z(data_out_imag[69]));
 BUF_X1 output130 (.A(net209),
    .Z(data_out_imag[6]));
 BUF_X1 output131 (.A(net210),
    .Z(data_out_imag[70]));
 BUF_X1 output132 (.A(net211),
    .Z(data_out_imag[71]));
 BUF_X1 output133 (.A(net212),
    .Z(data_out_imag[72]));
 BUF_X1 output134 (.A(net213),
    .Z(data_out_imag[73]));
 BUF_X1 output135 (.A(net214),
    .Z(data_out_imag[74]));
 BUF_X1 output136 (.A(net215),
    .Z(data_out_imag[75]));
 BUF_X1 output137 (.A(net216),
    .Z(data_out_imag[76]));
 BUF_X1 output138 (.A(net217),
    .Z(data_out_imag[77]));
 BUF_X1 output139 (.A(net218),
    .Z(data_out_imag[78]));
 BUF_X1 output140 (.A(net219),
    .Z(data_out_imag[79]));
 BUF_X1 output141 (.A(net220),
    .Z(data_out_imag[7]));
 BUF_X1 output142 (.A(net221),
    .Z(data_out_imag[80]));
 BUF_X1 output143 (.A(net222),
    .Z(data_out_imag[81]));
 BUF_X1 output144 (.A(net223),
    .Z(data_out_imag[82]));
 BUF_X1 output145 (.A(net224),
    .Z(data_out_imag[83]));
 BUF_X1 output146 (.A(net225),
    .Z(data_out_imag[84]));
 BUF_X1 output147 (.A(net226),
    .Z(data_out_imag[85]));
 BUF_X1 output148 (.A(net227),
    .Z(data_out_imag[86]));
 BUF_X1 output149 (.A(net228),
    .Z(data_out_imag[87]));
 BUF_X1 output150 (.A(net229),
    .Z(data_out_imag[88]));
 BUF_X1 output151 (.A(net230),
    .Z(data_out_imag[89]));
 BUF_X1 output152 (.A(net231),
    .Z(data_out_imag[8]));
 BUF_X1 output153 (.A(net232),
    .Z(data_out_imag[90]));
 BUF_X1 output154 (.A(net233),
    .Z(data_out_imag[91]));
 BUF_X1 output155 (.A(net234),
    .Z(data_out_imag[92]));
 BUF_X1 output156 (.A(net235),
    .Z(data_out_imag[93]));
 BUF_X1 output157 (.A(net236),
    .Z(data_out_imag[94]));
 BUF_X1 output158 (.A(net237),
    .Z(data_out_imag[95]));
 BUF_X1 output159 (.A(net238),
    .Z(data_out_imag[96]));
 BUF_X1 output160 (.A(net239),
    .Z(data_out_imag[97]));
 BUF_X1 output161 (.A(net240),
    .Z(data_out_imag[98]));
 BUF_X1 output162 (.A(net241),
    .Z(data_out_imag[99]));
 BUF_X1 output163 (.A(net242),
    .Z(data_out_imag[9]));
 BUF_X1 output164 (.A(net243),
    .Z(data_out_real[0]));
 BUF_X1 output165 (.A(net244),
    .Z(data_out_real[100]));
 BUF_X1 output166 (.A(net245),
    .Z(data_out_real[101]));
 BUF_X1 output167 (.A(net246),
    .Z(data_out_real[102]));
 BUF_X1 output168 (.A(net247),
    .Z(data_out_real[103]));
 BUF_X1 output169 (.A(net248),
    .Z(data_out_real[104]));
 BUF_X1 output170 (.A(net249),
    .Z(data_out_real[105]));
 BUF_X1 output171 (.A(net250),
    .Z(data_out_real[106]));
 BUF_X1 output172 (.A(net251),
    .Z(data_out_real[107]));
 BUF_X1 output173 (.A(net252),
    .Z(data_out_real[108]));
 BUF_X1 output174 (.A(net253),
    .Z(data_out_real[109]));
 BUF_X1 output175 (.A(net254),
    .Z(data_out_real[10]));
 BUF_X1 output176 (.A(net255),
    .Z(data_out_real[110]));
 BUF_X1 output177 (.A(net256),
    .Z(data_out_real[111]));
 BUF_X1 output178 (.A(net257),
    .Z(data_out_real[112]));
 BUF_X1 output179 (.A(net258),
    .Z(data_out_real[113]));
 BUF_X1 output180 (.A(net259),
    .Z(data_out_real[114]));
 BUF_X1 output181 (.A(net260),
    .Z(data_out_real[115]));
 BUF_X1 output182 (.A(net261),
    .Z(data_out_real[116]));
 BUF_X1 output183 (.A(net262),
    .Z(data_out_real[117]));
 BUF_X1 output184 (.A(net263),
    .Z(data_out_real[118]));
 BUF_X1 output185 (.A(net264),
    .Z(data_out_real[119]));
 BUF_X1 output186 (.A(net265),
    .Z(data_out_real[11]));
 BUF_X1 output187 (.A(net266),
    .Z(data_out_real[120]));
 BUF_X1 output188 (.A(net267),
    .Z(data_out_real[121]));
 BUF_X1 output189 (.A(net268),
    .Z(data_out_real[122]));
 BUF_X1 output190 (.A(net269),
    .Z(data_out_real[123]));
 BUF_X1 output191 (.A(net270),
    .Z(data_out_real[124]));
 BUF_X1 output192 (.A(net271),
    .Z(data_out_real[125]));
 BUF_X1 output193 (.A(net272),
    .Z(data_out_real[126]));
 BUF_X1 output194 (.A(net273),
    .Z(data_out_real[127]));
 BUF_X1 output195 (.A(net274),
    .Z(data_out_real[12]));
 BUF_X1 output196 (.A(net275),
    .Z(data_out_real[13]));
 BUF_X1 output197 (.A(net276),
    .Z(data_out_real[14]));
 BUF_X1 output198 (.A(net277),
    .Z(data_out_real[15]));
 BUF_X1 output199 (.A(net278),
    .Z(data_out_real[16]));
 BUF_X1 output200 (.A(net279),
    .Z(data_out_real[17]));
 BUF_X1 output201 (.A(net280),
    .Z(data_out_real[18]));
 BUF_X1 output202 (.A(net281),
    .Z(data_out_real[19]));
 BUF_X1 output203 (.A(net282),
    .Z(data_out_real[1]));
 BUF_X1 output204 (.A(net283),
    .Z(data_out_real[20]));
 BUF_X1 output205 (.A(net284),
    .Z(data_out_real[21]));
 BUF_X1 output206 (.A(net285),
    .Z(data_out_real[22]));
 BUF_X1 output207 (.A(net286),
    .Z(data_out_real[23]));
 BUF_X1 output208 (.A(net287),
    .Z(data_out_real[24]));
 BUF_X1 output209 (.A(net288),
    .Z(data_out_real[25]));
 BUF_X1 output210 (.A(net289),
    .Z(data_out_real[26]));
 BUF_X1 output211 (.A(net290),
    .Z(data_out_real[27]));
 BUF_X1 output212 (.A(net291),
    .Z(data_out_real[28]));
 BUF_X1 output213 (.A(net292),
    .Z(data_out_real[29]));
 BUF_X1 output214 (.A(net293),
    .Z(data_out_real[2]));
 BUF_X1 output215 (.A(net294),
    .Z(data_out_real[30]));
 BUF_X1 output216 (.A(net295),
    .Z(data_out_real[31]));
 BUF_X1 output217 (.A(net296),
    .Z(data_out_real[32]));
 BUF_X1 output218 (.A(net297),
    .Z(data_out_real[33]));
 BUF_X1 output219 (.A(net298),
    .Z(data_out_real[34]));
 BUF_X1 output220 (.A(net299),
    .Z(data_out_real[35]));
 BUF_X1 output221 (.A(net300),
    .Z(data_out_real[36]));
 BUF_X1 output222 (.A(net301),
    .Z(data_out_real[37]));
 BUF_X1 output223 (.A(net302),
    .Z(data_out_real[38]));
 BUF_X1 output224 (.A(net303),
    .Z(data_out_real[39]));
 BUF_X1 output225 (.A(net304),
    .Z(data_out_real[3]));
 BUF_X1 output226 (.A(net305),
    .Z(data_out_real[40]));
 BUF_X1 output227 (.A(net306),
    .Z(data_out_real[41]));
 BUF_X1 output228 (.A(net307),
    .Z(data_out_real[42]));
 BUF_X1 output229 (.A(net308),
    .Z(data_out_real[43]));
 BUF_X1 output230 (.A(net309),
    .Z(data_out_real[44]));
 BUF_X1 output231 (.A(net310),
    .Z(data_out_real[45]));
 BUF_X1 output232 (.A(net311),
    .Z(data_out_real[46]));
 BUF_X1 output233 (.A(net312),
    .Z(data_out_real[47]));
 BUF_X1 output234 (.A(net313),
    .Z(data_out_real[48]));
 BUF_X1 output235 (.A(net314),
    .Z(data_out_real[49]));
 BUF_X1 output236 (.A(net315),
    .Z(data_out_real[4]));
 BUF_X1 output237 (.A(net316),
    .Z(data_out_real[50]));
 BUF_X1 output238 (.A(net317),
    .Z(data_out_real[51]));
 BUF_X1 output239 (.A(net318),
    .Z(data_out_real[52]));
 BUF_X1 output240 (.A(net319),
    .Z(data_out_real[53]));
 BUF_X1 output241 (.A(net320),
    .Z(data_out_real[54]));
 BUF_X1 output242 (.A(net321),
    .Z(data_out_real[55]));
 BUF_X1 output243 (.A(net322),
    .Z(data_out_real[56]));
 BUF_X1 output244 (.A(net323),
    .Z(data_out_real[57]));
 BUF_X1 output245 (.A(net324),
    .Z(data_out_real[58]));
 BUF_X1 output246 (.A(net325),
    .Z(data_out_real[59]));
 BUF_X1 output247 (.A(net326),
    .Z(data_out_real[5]));
 BUF_X1 output248 (.A(net327),
    .Z(data_out_real[60]));
 BUF_X1 output249 (.A(net328),
    .Z(data_out_real[61]));
 BUF_X1 output250 (.A(net329),
    .Z(data_out_real[62]));
 BUF_X1 output251 (.A(net330),
    .Z(data_out_real[63]));
 BUF_X1 output252 (.A(net331),
    .Z(data_out_real[64]));
 BUF_X1 output253 (.A(net332),
    .Z(data_out_real[65]));
 BUF_X1 output254 (.A(net333),
    .Z(data_out_real[66]));
 BUF_X1 output255 (.A(net334),
    .Z(data_out_real[67]));
 BUF_X1 output256 (.A(net335),
    .Z(data_out_real[68]));
 BUF_X1 output257 (.A(net336),
    .Z(data_out_real[69]));
 BUF_X1 output258 (.A(net337),
    .Z(data_out_real[6]));
 BUF_X1 output259 (.A(net338),
    .Z(data_out_real[70]));
 BUF_X1 output260 (.A(net339),
    .Z(data_out_real[71]));
 BUF_X1 output261 (.A(net340),
    .Z(data_out_real[72]));
 BUF_X1 output262 (.A(net341),
    .Z(data_out_real[73]));
 BUF_X1 output263 (.A(net342),
    .Z(data_out_real[74]));
 BUF_X1 output264 (.A(net343),
    .Z(data_out_real[75]));
 BUF_X1 output265 (.A(net344),
    .Z(data_out_real[76]));
 BUF_X1 output266 (.A(net345),
    .Z(data_out_real[77]));
 BUF_X1 output267 (.A(net346),
    .Z(data_out_real[78]));
 BUF_X1 output268 (.A(net347),
    .Z(data_out_real[79]));
 BUF_X1 output269 (.A(net348),
    .Z(data_out_real[7]));
 BUF_X1 output270 (.A(net349),
    .Z(data_out_real[80]));
 BUF_X1 output271 (.A(net350),
    .Z(data_out_real[81]));
 BUF_X1 output272 (.A(net351),
    .Z(data_out_real[82]));
 BUF_X1 output273 (.A(net352),
    .Z(data_out_real[83]));
 BUF_X1 output274 (.A(net353),
    .Z(data_out_real[84]));
 BUF_X1 output275 (.A(net354),
    .Z(data_out_real[85]));
 BUF_X1 output276 (.A(net355),
    .Z(data_out_real[86]));
 BUF_X1 output277 (.A(net356),
    .Z(data_out_real[87]));
 BUF_X1 output278 (.A(net357),
    .Z(data_out_real[88]));
 BUF_X1 output279 (.A(net358),
    .Z(data_out_real[89]));
 BUF_X1 output280 (.A(net359),
    .Z(data_out_real[8]));
 BUF_X1 output281 (.A(net360),
    .Z(data_out_real[90]));
 BUF_X1 output282 (.A(net361),
    .Z(data_out_real[91]));
 BUF_X1 output283 (.A(net362),
    .Z(data_out_real[92]));
 BUF_X1 output284 (.A(net363),
    .Z(data_out_real[93]));
 BUF_X1 output285 (.A(net364),
    .Z(data_out_real[94]));
 BUF_X1 output286 (.A(net365),
    .Z(data_out_real[95]));
 BUF_X1 output287 (.A(net366),
    .Z(data_out_real[96]));
 BUF_X1 output288 (.A(net367),
    .Z(data_out_real[97]));
 BUF_X1 output289 (.A(net368),
    .Z(data_out_real[98]));
 BUF_X1 output290 (.A(net369),
    .Z(data_out_real[99]));
 BUF_X1 output291 (.A(net370),
    .Z(data_out_real[9]));
 BUF_X1 output292 (.A(net371),
    .Z(data_ready));
 BUF_X1 output293 (.A(net372),
    .Z(data_valid_out));
 BUF_X2 max_cap294 (.A(_04439_),
    .Z(net373));
 BUF_X2 max_cap295 (.A(_04410_),
    .Z(net374));
 BUF_X2 max_cap296 (.A(_04046_),
    .Z(net375));
 CLKBUF_X3 wire297 (.A(_03637_),
    .Z(net376));
 CLKBUF_X2 max_cap298 (.A(_03341_),
    .Z(net377));
 BUF_X2 max_cap299 (.A(_02987_),
    .Z(net378));
 BUF_X1 max_cap300 (.A(net380),
    .Z(net379));
 BUF_X1 max_cap301 (.A(_02709_),
    .Z(net380));
 BUF_X2 max_cap302 (.A(net382),
    .Z(net381));
 BUF_X2 max_cap303 (.A(_02004_),
    .Z(net382));
 BUF_X4 max_cap304 (.A(_01108_),
    .Z(net383));
 LOGIC0_X1 _17624__305 (.Z(net384));
 LOGIC0_X1 _17633__306 (.Z(net385));
 LOGIC0_X1 _17646__307 (.Z(net386));
 LOGIC0_X1 _17660__308 (.Z(net387));
 LOGIC0_X1 _17670__309 (.Z(net388));
 LOGIC0_X1 _17686__310 (.Z(net389));
 LOGIC0_X1 _17702__311 (.Z(net390));
 LOGIC0_X1 _17710__312 (.Z(net391));
 LOGIC0_X1 _17724__313 (.Z(net392));
 LOGIC0_X1 _17742__314 (.Z(net393));
 LOGIC0_X1 _17758__315 (.Z(net394));
 LOGIC0_X1 _17766__316 (.Z(net395));
 LOGIC0_X1 _17783__317 (.Z(net396));
 LOGIC0_X1 _17797__318 (.Z(net397));
 CLKBUF_X3 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_1_clk));
 CLKBUF_X3 clkbuf_leaf_2_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_2_clk));
 CLKBUF_X3 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_3_clk));
 CLKBUF_X3 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_4_clk));
 CLKBUF_X3 clkbuf_leaf_5_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_5_clk));
 CLKBUF_X3 clkbuf_leaf_6_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_6_clk));
 CLKBUF_X3 clkbuf_leaf_7_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_7_clk));
 CLKBUF_X3 clkbuf_leaf_8_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_8_clk));
 CLKBUF_X3 clkbuf_leaf_9_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_9_clk));
 CLKBUF_X3 clkbuf_leaf_10_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_10_clk));
 CLKBUF_X3 clkbuf_leaf_11_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_11_clk));
 CLKBUF_X3 clkbuf_leaf_12_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_12_clk));
 CLKBUF_X3 clkbuf_leaf_13_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_13_clk));
 CLKBUF_X3 clkbuf_leaf_14_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_14_clk));
 CLKBUF_X3 clkbuf_leaf_15_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_15_clk));
 CLKBUF_X3 clkbuf_leaf_16_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_16_clk));
 CLKBUF_X3 clkbuf_leaf_17_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_17_clk));
 CLKBUF_X3 clkbuf_leaf_18_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_18_clk));
 CLKBUF_X3 clkbuf_leaf_19_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_19_clk));
 CLKBUF_X3 clkbuf_leaf_20_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_20_clk));
 CLKBUF_X3 clkbuf_leaf_21_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_21_clk));
 CLKBUF_X3 clkbuf_leaf_22_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_22_clk));
 CLKBUF_X3 clkbuf_leaf_23_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_23_clk));
 CLKBUF_X3 clkbuf_leaf_24_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_24_clk));
 CLKBUF_X3 clkbuf_leaf_25_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_25_clk));
 CLKBUF_X3 clkbuf_leaf_26_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_26_clk));
 CLKBUF_X3 clkbuf_leaf_27_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_27_clk));
 CLKBUF_X3 clkbuf_leaf_28_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_28_clk));
 CLKBUF_X3 clkbuf_leaf_29_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_29_clk));
 CLKBUF_X3 clkbuf_leaf_30_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_30_clk));
 CLKBUF_X3 clkbuf_leaf_31_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_31_clk));
 CLKBUF_X3 clkbuf_leaf_32_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_32_clk));
 CLKBUF_X3 clkbuf_leaf_33_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_33_clk));
 CLKBUF_X3 clkbuf_leaf_34_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_34_clk));
 CLKBUF_X3 clkbuf_leaf_35_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_35_clk));
 CLKBUF_X3 clkbuf_leaf_36_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_36_clk));
 CLKBUF_X3 clkbuf_leaf_37_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_37_clk));
 CLKBUF_X3 clkbuf_leaf_38_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_38_clk));
 CLKBUF_X3 clkbuf_leaf_39_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_39_clk));
 CLKBUF_X3 clkbuf_leaf_40_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_40_clk));
 CLKBUF_X3 clkbuf_leaf_41_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_41_clk));
 CLKBUF_X3 clkbuf_leaf_42_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_42_clk));
 CLKBUF_X3 clkbuf_leaf_43_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_43_clk));
 CLKBUF_X3 clkbuf_leaf_44_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_44_clk));
 CLKBUF_X3 clkbuf_leaf_45_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_45_clk));
 CLKBUF_X3 clkbuf_leaf_46_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_46_clk));
 CLKBUF_X3 clkbuf_leaf_47_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_47_clk));
 CLKBUF_X3 clkbuf_leaf_48_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_48_clk));
 CLKBUF_X3 clkbuf_leaf_49_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_49_clk));
 CLKBUF_X3 clkbuf_leaf_50_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_50_clk));
 CLKBUF_X3 clkbuf_leaf_51_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_51_clk));
 CLKBUF_X3 clkbuf_leaf_52_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_52_clk));
 CLKBUF_X3 clkbuf_leaf_53_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_53_clk));
 CLKBUF_X3 clkbuf_leaf_54_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_54_clk));
 CLKBUF_X3 clkbuf_leaf_55_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_55_clk));
 CLKBUF_X3 clkbuf_leaf_56_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_56_clk));
 CLKBUF_X3 clkbuf_leaf_57_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_57_clk));
 CLKBUF_X3 clkbuf_leaf_58_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_58_clk));
 CLKBUF_X3 clkbuf_leaf_59_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_59_clk));
 CLKBUF_X3 clkbuf_leaf_60_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_60_clk));
 CLKBUF_X3 clkbuf_leaf_61_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_61_clk));
 CLKBUF_X3 clkbuf_leaf_62_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_62_clk));
 CLKBUF_X3 clkbuf_leaf_63_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_63_clk));
 CLKBUF_X3 clkbuf_leaf_64_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_64_clk));
 CLKBUF_X3 clkbuf_leaf_65_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_65_clk));
 CLKBUF_X3 clkbuf_leaf_66_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_66_clk));
 CLKBUF_X3 clkbuf_leaf_67_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_67_clk));
 CLKBUF_X3 clkbuf_leaf_68_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_68_clk));
 CLKBUF_X3 clkbuf_leaf_69_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_69_clk));
 CLKBUF_X3 clkbuf_leaf_70_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_70_clk));
 CLKBUF_X3 clkbuf_leaf_71_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_71_clk));
 CLKBUF_X3 clkbuf_leaf_72_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_72_clk));
 CLKBUF_X3 clkbuf_leaf_73_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_73_clk));
 CLKBUF_X3 clkbuf_leaf_74_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_74_clk));
 CLKBUF_X3 clkbuf_leaf_75_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_75_clk));
 CLKBUF_X3 clkbuf_leaf_76_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_76_clk));
 CLKBUF_X3 clkbuf_leaf_77_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_77_clk));
 CLKBUF_X3 clkbuf_leaf_78_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_78_clk));
 CLKBUF_X3 clkbuf_leaf_79_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_79_clk));
 CLKBUF_X3 clkbuf_leaf_80_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_80_clk));
 CLKBUF_X3 clkbuf_leaf_81_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_81_clk));
 CLKBUF_X3 clkbuf_leaf_82_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_82_clk));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_0__leaf_clk));
 CLKBUF_X3 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_1__leaf_clk));
 CLKBUF_X3 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_2__leaf_clk));
 CLKBUF_X3 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_3__leaf_clk));
 CLKBUF_X3 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_4__leaf_clk));
 CLKBUF_X3 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_5__leaf_clk));
 CLKBUF_X3 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_6__leaf_clk));
 CLKBUF_X3 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_7__leaf_clk));
 INV_X4 clkload0 (.A(clknet_3_0__leaf_clk));
 INV_X2 clkload1 (.A(clknet_3_1__leaf_clk));
 INV_X4 clkload2 (.A(clknet_3_2__leaf_clk));
 INV_X4 clkload3 (.A(clknet_3_4__leaf_clk));
 INV_X2 clkload4 (.A(clknet_3_5__leaf_clk));
 CLKBUF_X3 clkload5 (.A(clknet_3_7__leaf_clk));
 CLKBUF_X1 clkload6 (.A(clknet_leaf_0_clk));
 INV_X1 clkload7 (.A(clknet_leaf_1_clk));
 CLKBUF_X1 clkload8 (.A(clknet_leaf_2_clk));
 CLKBUF_X1 clkload9 (.A(clknet_leaf_8_clk));
 CLKBUF_X1 clkload10 (.A(clknet_leaf_80_clk));
 CLKBUF_X1 clkload11 (.A(clknet_leaf_81_clk));
 INV_X2 clkload12 (.A(clknet_leaf_3_clk));
 CLKBUF_X1 clkload13 (.A(clknet_leaf_4_clk));
 CLKBUF_X1 clkload14 (.A(clknet_leaf_5_clk));
 INV_X1 clkload15 (.A(clknet_leaf_6_clk));
 CLKBUF_X1 clkload16 (.A(clknet_leaf_7_clk));
 CLKBUF_X1 clkload17 (.A(clknet_leaf_10_clk));
 CLKBUF_X1 clkload18 (.A(clknet_leaf_12_clk));
 INV_X1 clkload19 (.A(clknet_leaf_13_clk));
 INV_X1 clkload20 (.A(clknet_leaf_37_clk));
 CLKBUF_X1 clkload21 (.A(clknet_leaf_14_clk));
 CLKBUF_X1 clkload22 (.A(clknet_leaf_15_clk));
 INV_X2 clkload23 (.A(clknet_leaf_24_clk));
 CLKBUF_X1 clkload24 (.A(clknet_leaf_34_clk));
 INV_X1 clkload25 (.A(clknet_leaf_35_clk));
 INV_X1 clkload26 (.A(clknet_leaf_36_clk));
 INV_X1 clkload27 (.A(clknet_leaf_19_clk));
 CLKBUF_X1 clkload28 (.A(clknet_leaf_20_clk));
 CLKBUF_X1 clkload29 (.A(clknet_leaf_21_clk));
 CLKBUF_X1 clkload30 (.A(clknet_leaf_22_clk));
 INV_X1 clkload31 (.A(clknet_leaf_25_clk));
 CLKBUF_X1 clkload32 (.A(clknet_leaf_26_clk));
 CLKBUF_X1 clkload33 (.A(clknet_leaf_27_clk));
 CLKBUF_X1 clkload34 (.A(clknet_leaf_28_clk));
 INV_X1 clkload35 (.A(clknet_leaf_29_clk));
 CLKBUF_X1 clkload36 (.A(clknet_leaf_30_clk));
 CLKBUF_X1 clkload37 (.A(clknet_leaf_31_clk));
 INV_X1 clkload38 (.A(clknet_leaf_33_clk));
 INV_X1 clkload39 (.A(clknet_leaf_72_clk));
 INV_X2 clkload40 (.A(clknet_leaf_73_clk));
 INV_X2 clkload41 (.A(clknet_leaf_74_clk));
 INV_X2 clkload42 (.A(clknet_leaf_75_clk));
 INV_X2 clkload43 (.A(clknet_leaf_76_clk));
 CLKBUF_X1 clkload44 (.A(clknet_leaf_77_clk));
 INV_X2 clkload45 (.A(clknet_leaf_78_clk));
 CLKBUF_X1 clkload46 (.A(clknet_leaf_38_clk));
 INV_X1 clkload47 (.A(clknet_leaf_39_clk));
 INV_X2 clkload48 (.A(clknet_leaf_40_clk));
 CLKBUF_X1 clkload49 (.A(clknet_leaf_65_clk));
 INV_X1 clkload50 (.A(clknet_leaf_66_clk));
 CLKBUF_X1 clkload51 (.A(clknet_leaf_67_clk));
 CLKBUF_X1 clkload52 (.A(clknet_leaf_68_clk));
 CLKBUF_X1 clkload53 (.A(clknet_leaf_70_clk));
 CLKBUF_X1 clkload54 (.A(clknet_leaf_71_clk));
 CLKBUF_X1 clkload55 (.A(clknet_leaf_52_clk));
 CLKBUF_X1 clkload56 (.A(clknet_leaf_53_clk));
 CLKBUF_X1 clkload57 (.A(clknet_leaf_54_clk));
 CLKBUF_X1 clkload58 (.A(clknet_leaf_55_clk));
 CLKBUF_X1 clkload59 (.A(clknet_leaf_57_clk));
 CLKBUF_X1 clkload60 (.A(clknet_leaf_58_clk));
 CLKBUF_X1 clkload61 (.A(clknet_leaf_60_clk));
 CLKBUF_X1 clkload62 (.A(clknet_leaf_61_clk));
 INV_X1 clkload63 (.A(clknet_leaf_62_clk));
 CLKBUF_X1 clkload64 (.A(clknet_leaf_63_clk));
 INV_X1 clkload65 (.A(clknet_leaf_64_clk));
 CLKBUF_X1 clkload66 (.A(clknet_leaf_32_clk));
 CLKBUF_X1 clkload67 (.A(clknet_leaf_41_clk));
 INV_X2 clkload68 (.A(clknet_leaf_42_clk));
 CLKBUF_X1 clkload69 (.A(clknet_leaf_43_clk));
 CLKBUF_X1 clkload70 (.A(clknet_leaf_44_clk));
 CLKBUF_X1 clkload71 (.A(clknet_leaf_46_clk));
 INV_X1 clkload72 (.A(clknet_leaf_47_clk));
 CLKBUF_X1 clkload73 (.A(clknet_leaf_48_clk));
 CLKBUF_X1 clkload74 (.A(clknet_leaf_49_clk));
 CLKBUF_X1 clkload75 (.A(clknet_leaf_50_clk));
 CLKBUF_X1 clkload76 (.A(clknet_leaf_51_clk));
 BUF_X1 rebuffer1 (.A(_04356_),
    .Z(net399));
 BUF_X1 rebuffer2 (.A(net399),
    .Z(net400));
 BUF_X1 rebuffer3 (.A(net399),
    .Z(net401));
 NAND3_X2 clone43 (.A1(net403),
    .A2(_03412_),
    .A3(_03473_),
    .ZN(net402));
 OAI22_X2 clone45 (.A1(_03351_),
    .A2(_03430_),
    .B1(_03432_),
    .B2(_03445_),
    .ZN(net403));
 BUF_X1 rebuffer46 (.A(_04247_),
    .Z(net404));
 BUF_X1 rebuffer47 (.A(_04248_),
    .Z(net405));
 BUF_X1 rebuffer48 (.A(_04248_),
    .Z(net406));
 BUF_X1 rebuffer49 (.A(_04096_),
    .Z(net407));
 BUF_X4 clone50 (.A(_04070_),
    .Z(net408));
 BUF_X1 rebuffer51 (.A(_09264_),
    .Z(net409));
 BUF_X1 rebuffer52 (.A(_04567_),
    .Z(net410));
 BUF_X1 rebuffer53 (.A(_04567_),
    .Z(net411));
 BUF_X1 rebuffer54 (.A(net414),
    .Z(net412));
 BUF_X1 rebuffer55 (.A(_04566_),
    .Z(net413));
 BUF_X1 rebuffer57 (.A(net416),
    .Z(net415));
 BUF_X1 rebuffer58 (.A(net417),
    .Z(net416));
 BUF_X1 rebuffer59 (.A(net418),
    .Z(net417));
 BUF_X1 rebuffer60 (.A(net419),
    .Z(net418));
 BUF_X1 rebuffer61 (.A(net420),
    .Z(net419));
 BUF_X1 rebuffer62 (.A(net421),
    .Z(net420));
 BUF_X1 rebuffer63 (.A(net422),
    .Z(net421));
 BUF_X4 rebuffer64 (.A(_04565_),
    .Z(net422));
 BUF_X1 rebuffer65 (.A(_04568_),
    .Z(net423));
 BUF_X4 clone66 (.A(_03053_),
    .Z(net424));
 BUF_X8 clone67 (.A(_02927_),
    .Z(net425));
 BUF_X1 rebuffer71 (.A(_04568_),
    .Z(net429));
 BUF_X1 rebuffer86 (.A(_08702_),
    .Z(net444));
 BUF_X1 rebuffer87 (.A(_08702_),
    .Z(net445));
 BUF_X1 rebuffer88 (.A(_08707_),
    .Z(net446));
 BUF_X1 rebuffer89 (.A(_08707_),
    .Z(net447));
 BUF_X1 rebuffer90 (.A(net474),
    .Z(net448));
 BUF_X1 rebuffer91 (.A(_05893_),
    .Z(net449));
 BUF_X1 rebuffer92 (.A(_05891_),
    .Z(net450));
 BUF_X2 rebuffer93 (.A(_05889_),
    .Z(net451));
 BUF_X2 rebuffer94 (.A(_00001_),
    .Z(net452));
 BUF_X16 rebuffer95 (.A(net485),
    .Z(net453));
 BUF_X1 rebuffer96 (.A(_05877_),
    .Z(net454));
 BUF_X1 rebuffer97 (.A(_05871_),
    .Z(net455));
 BUF_X1 rebuffer98 (.A(_05906_),
    .Z(net456));
 BUF_X1 rebuffer99 (.A(_07358_),
    .Z(net457));
 BUF_X16 rebuffer100 (.A(_00873_),
    .Z(net458));
 BUF_X1 rebuffer101 (.A(_05900_),
    .Z(net459));
 BUF_X2 rebuffer116 (.A(_08707_),
    .Z(net474));
 BUF_X1 rebuffer117 (.A(net458),
    .Z(net475));
 BUF_X1 rebuffer118 (.A(net130),
    .Z(net476));
 BUF_X1 rebuffer119 (.A(net130),
    .Z(net477));
 BUF_X1 rebuffer120 (.A(_05856_),
    .Z(net478));
 BUF_X4 rebuffer123 (.A(_08637_),
    .Z(net481));
 BUF_X16 clone124 (.A(_06065_),
    .Z(net482));
 BUF_X8 clone126 (.A(_06092_),
    .Z(net483));
 BUF_X16 clone141 (.A(_05936_),
    .Z(net491));
 BUF_X2 rebuffer143 (.A(_08626_),
    .Z(net493));
 BUF_X1 rebuffer144 (.A(net493),
    .Z(net494));
 BUF_X1 rebuffer145 (.A(_08626_),
    .Z(net495));
 BUF_X1 rebuffer146 (.A(_05418_),
    .Z(net496));
 BUF_X4 rebuffer147 (.A(_05419_),
    .Z(net497));
 BUF_X1 rebuffer148 (.A(_05394_),
    .Z(net498));
 BUF_X4 rebuffer149 (.A(_05390_),
    .Z(net499));
 BUF_X1 rebuffer150 (.A(_07350_),
    .Z(net500));
 BUF_X1 rebuffer151 (.A(_05382_),
    .Z(net501));
 BUF_X1 rebuffer152 (.A(_05388_),
    .Z(net502));
 BUF_X1 rebuffer153 (.A(_05375_),
    .Z(net503));
 BUF_X4 rebuffer154 (.A(_05392_),
    .Z(net504));
 BUF_X1 rebuffer155 (.A(net508),
    .Z(net505));
 BUF_X1 rebuffer156 (.A(_05373_),
    .Z(net506));
 BUF_X1 rebuffer157 (.A(_05386_),
    .Z(net507));
 BUF_X2 rebuffer158 (.A(_05384_),
    .Z(net508));
 BUF_X4 rebuffer159 (.A(_05377_),
    .Z(net509));
 BUF_X1 rebuffer160 (.A(_05371_),
    .Z(net510));
 BUF_X1 rebuffer162 (.A(_05414_),
    .Z(net512));
 BUF_X1 rebuffer164 (.A(_06198_),
    .Z(net514));
 BUF_X2 rebuffer165 (.A(_06225_),
    .Z(net515));
 BUF_X16 clone166 (.A(_06227_),
    .Z(net516));
 BUF_X2 rebuffer167 (.A(_06144_),
    .Z(net517));
 BUF_X2 rebuffer168 (.A(net487),
    .Z(net518));
 BUF_X1 rebuffer129 (.A(_05338_),
    .Z(net520));
 BUF_X2 max_cap1 (.A(_04046_),
    .Z(net426));
 NOR2_X2 clone47 (.A1(_03504_),
    .A2(_03505_),
    .ZN(net428));
 BUF_X4 rebuffer73 (.A(_04882_),
    .Z(net437));
 BUF_X1 rebuffer74 (.A(_04962_),
    .Z(net438));
 BUF_X2 rebuffer79 (.A(_05926_),
    .Z(net443));
 BUF_X1 rebuffer80 (.A(net443),
    .Z(net460));
 BUF_X4 rebuffer81 (.A(_05930_),
    .Z(net461));
 BUF_X1 rebuffer82 (.A(_05921_),
    .Z(net462));
 BUF_X1 rebuffer83 (.A(_05886_),
    .Z(net463));
 BUF_X1 rebuffer84 (.A(_05901_),
    .Z(net464));
 AND2_X2 clone106 (.A1(_05859_),
    .A2(_05298_),
    .ZN(net470));
 BUF_X8 rebuffer113 (.A(_05929_),
    .Z(net485));
 BUF_X8 rebuffer114 (.A(_06065_),
    .Z(net486));
 BUF_X4 rebuffer115 (.A(_06171_),
    .Z(net487));
 BUF_X4 rebuffer121 (.A(net534),
    .Z(net488));
 BUF_X1 rebuffer122 (.A(_05367_),
    .Z(net489));
 BUF_X16 rebuffer126 (.A(_00931_),
    .Z(net511));
 BUF_X4 rebuffer127 (.A(_05577_),
    .Z(net513));
 BUF_X1 rebuffer130 (.A(_08629_),
    .Z(net521));
 BUF_X1 rebuffer131 (.A(_08619_),
    .Z(net522));
 BUF_X8 rebuffer133 (.A(_06092_),
    .Z(net524));
 BUF_X4 rebuffer135 (.A(_05342_),
    .Z(net526));
 BUF_X1 rebuffer136 (.A(_05723_),
    .Z(net527));
 BUF_X4 rebuffer137 (.A(_05468_),
    .Z(net528));
 BUF_X2 rebuffer138 (.A(_05475_),
    .Z(net529));
 BUF_X4 rebuffer139 (.A(_05431_),
    .Z(net530));
 BUF_X8 rebuffer140 (.A(_05508_),
    .Z(net531));
 BUF_X4 rebuffer163 (.A(_05577_),
    .Z(net534));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X32 FILLER_0_129 ();
 FILLCELL_X32 FILLER_0_161 ();
 FILLCELL_X32 FILLER_0_193 ();
 FILLCELL_X32 FILLER_0_225 ();
 FILLCELL_X1 FILLER_0_263 ();
 FILLCELL_X16 FILLER_0_267 ();
 FILLCELL_X2 FILLER_0_286 ();
 FILLCELL_X1 FILLER_0_288 ();
 FILLCELL_X32 FILLER_0_295 ();
 FILLCELL_X16 FILLER_0_327 ();
 FILLCELL_X4 FILLER_0_343 ();
 FILLCELL_X4 FILLER_0_354 ();
 FILLCELL_X1 FILLER_0_358 ();
 FILLCELL_X32 FILLER_0_369 ();
 FILLCELL_X16 FILLER_0_401 ();
 FILLCELL_X8 FILLER_0_417 ();
 FILLCELL_X2 FILLER_0_425 ();
 FILLCELL_X1 FILLER_0_427 ();
 FILLCELL_X32 FILLER_0_434 ();
 FILLCELL_X32 FILLER_0_466 ();
 FILLCELL_X32 FILLER_0_498 ();
 FILLCELL_X32 FILLER_0_530 ();
 FILLCELL_X32 FILLER_0_562 ();
 FILLCELL_X32 FILLER_0_594 ();
 FILLCELL_X4 FILLER_0_626 ();
 FILLCELL_X1 FILLER_0_630 ();
 FILLCELL_X16 FILLER_0_632 ();
 FILLCELL_X8 FILLER_0_648 ();
 FILLCELL_X2 FILLER_0_656 ();
 FILLCELL_X1 FILLER_0_658 ();
 FILLCELL_X32 FILLER_0_663 ();
 FILLCELL_X32 FILLER_0_695 ();
 FILLCELL_X32 FILLER_0_727 ();
 FILLCELL_X32 FILLER_0_759 ();
 FILLCELL_X32 FILLER_0_791 ();
 FILLCELL_X32 FILLER_0_823 ();
 FILLCELL_X32 FILLER_0_855 ();
 FILLCELL_X32 FILLER_0_887 ();
 FILLCELL_X32 FILLER_0_919 ();
 FILLCELL_X16 FILLER_0_951 ();
 FILLCELL_X8 FILLER_0_967 ();
 FILLCELL_X4 FILLER_0_975 ();
 FILLCELL_X2 FILLER_0_979 ();
 FILLCELL_X1 FILLER_0_981 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X16 FILLER_1_257 ();
 FILLCELL_X1 FILLER_1_273 ();
 FILLCELL_X8 FILLER_1_313 ();
 FILLCELL_X2 FILLER_1_349 ();
 FILLCELL_X1 FILLER_1_358 ();
 FILLCELL_X8 FILLER_1_384 ();
 FILLCELL_X2 FILLER_1_392 ();
 FILLCELL_X1 FILLER_1_394 ();
 FILLCELL_X2 FILLER_1_397 ();
 FILLCELL_X2 FILLER_1_409 ();
 FILLCELL_X32 FILLER_1_420 ();
 FILLCELL_X32 FILLER_1_452 ();
 FILLCELL_X32 FILLER_1_484 ();
 FILLCELL_X16 FILLER_1_516 ();
 FILLCELL_X8 FILLER_1_532 ();
 FILLCELL_X2 FILLER_1_540 ();
 FILLCELL_X1 FILLER_1_542 ();
 FILLCELL_X32 FILLER_1_549 ();
 FILLCELL_X1 FILLER_1_581 ();
 FILLCELL_X1 FILLER_1_599 ();
 FILLCELL_X16 FILLER_1_607 ();
 FILLCELL_X4 FILLER_1_623 ();
 FILLCELL_X4 FILLER_1_641 ();
 FILLCELL_X2 FILLER_1_648 ();
 FILLCELL_X1 FILLER_1_650 ();
 FILLCELL_X2 FILLER_1_659 ();
 FILLCELL_X1 FILLER_1_661 ();
 FILLCELL_X1 FILLER_1_667 ();
 FILLCELL_X2 FILLER_1_681 ();
 FILLCELL_X1 FILLER_1_683 ();
 FILLCELL_X4 FILLER_1_693 ();
 FILLCELL_X8 FILLER_1_700 ();
 FILLCELL_X4 FILLER_1_708 ();
 FILLCELL_X2 FILLER_1_726 ();
 FILLCELL_X1 FILLER_1_728 ();
 FILLCELL_X4 FILLER_1_745 ();
 FILLCELL_X1 FILLER_1_749 ();
 FILLCELL_X4 FILLER_1_763 ();
 FILLCELL_X1 FILLER_1_767 ();
 FILLCELL_X1 FILLER_1_774 ();
 FILLCELL_X32 FILLER_1_788 ();
 FILLCELL_X32 FILLER_1_820 ();
 FILLCELL_X32 FILLER_1_852 ();
 FILLCELL_X32 FILLER_1_884 ();
 FILLCELL_X32 FILLER_1_916 ();
 FILLCELL_X32 FILLER_1_948 ();
 FILLCELL_X2 FILLER_1_980 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X16 FILLER_2_257 ();
 FILLCELL_X8 FILLER_2_273 ();
 FILLCELL_X4 FILLER_2_281 ();
 FILLCELL_X1 FILLER_2_285 ();
 FILLCELL_X1 FILLER_2_310 ();
 FILLCELL_X4 FILLER_2_314 ();
 FILLCELL_X1 FILLER_2_318 ();
 FILLCELL_X1 FILLER_2_353 ();
 FILLCELL_X2 FILLER_2_363 ();
 FILLCELL_X1 FILLER_2_365 ();
 FILLCELL_X1 FILLER_2_378 ();
 FILLCELL_X2 FILLER_2_389 ();
 FILLCELL_X8 FILLER_2_395 ();
 FILLCELL_X4 FILLER_2_403 ();
 FILLCELL_X2 FILLER_2_407 ();
 FILLCELL_X1 FILLER_2_412 ();
 FILLCELL_X32 FILLER_2_433 ();
 FILLCELL_X32 FILLER_2_465 ();
 FILLCELL_X8 FILLER_2_510 ();
 FILLCELL_X4 FILLER_2_518 ();
 FILLCELL_X1 FILLER_2_522 ();
 FILLCELL_X8 FILLER_2_525 ();
 FILLCELL_X4 FILLER_2_533 ();
 FILLCELL_X4 FILLER_2_544 ();
 FILLCELL_X2 FILLER_2_586 ();
 FILLCELL_X1 FILLER_2_588 ();
 FILLCELL_X1 FILLER_2_598 ();
 FILLCELL_X1 FILLER_2_603 ();
 FILLCELL_X2 FILLER_2_611 ();
 FILLCELL_X8 FILLER_2_623 ();
 FILLCELL_X2 FILLER_2_632 ();
 FILLCELL_X1 FILLER_2_634 ();
 FILLCELL_X1 FILLER_2_662 ();
 FILLCELL_X1 FILLER_2_699 ();
 FILLCELL_X1 FILLER_2_704 ();
 FILLCELL_X1 FILLER_2_707 ();
 FILLCELL_X4 FILLER_2_712 ();
 FILLCELL_X2 FILLER_2_716 ();
 FILLCELL_X2 FILLER_2_738 ();
 FILLCELL_X1 FILLER_2_740 ();
 FILLCELL_X32 FILLER_2_789 ();
 FILLCELL_X32 FILLER_2_821 ();
 FILLCELL_X32 FILLER_2_853 ();
 FILLCELL_X32 FILLER_2_885 ();
 FILLCELL_X32 FILLER_2_917 ();
 FILLCELL_X32 FILLER_2_949 ();
 FILLCELL_X1 FILLER_2_981 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X16 FILLER_3_161 ();
 FILLCELL_X8 FILLER_3_177 ();
 FILLCELL_X4 FILLER_3_185 ();
 FILLCELL_X2 FILLER_3_189 ();
 FILLCELL_X32 FILLER_3_200 ();
 FILLCELL_X16 FILLER_3_232 ();
 FILLCELL_X8 FILLER_3_248 ();
 FILLCELL_X4 FILLER_3_256 ();
 FILLCELL_X2 FILLER_3_260 ();
 FILLCELL_X2 FILLER_3_276 ();
 FILLCELL_X2 FILLER_3_284 ();
 FILLCELL_X4 FILLER_3_318 ();
 FILLCELL_X2 FILLER_3_322 ();
 FILLCELL_X1 FILLER_3_324 ();
 FILLCELL_X4 FILLER_3_327 ();
 FILLCELL_X2 FILLER_3_353 ();
 FILLCELL_X4 FILLER_3_399 ();
 FILLCELL_X1 FILLER_3_403 ();
 FILLCELL_X32 FILLER_3_430 ();
 FILLCELL_X32 FILLER_3_462 ();
 FILLCELL_X4 FILLER_3_494 ();
 FILLCELL_X1 FILLER_3_498 ();
 FILLCELL_X2 FILLER_3_506 ();
 FILLCELL_X1 FILLER_3_517 ();
 FILLCELL_X1 FILLER_3_541 ();
 FILLCELL_X1 FILLER_3_557 ();
 FILLCELL_X1 FILLER_3_569 ();
 FILLCELL_X1 FILLER_3_581 ();
 FILLCELL_X2 FILLER_3_587 ();
 FILLCELL_X1 FILLER_3_589 ();
 FILLCELL_X1 FILLER_3_600 ();
 FILLCELL_X1 FILLER_3_607 ();
 FILLCELL_X8 FILLER_3_612 ();
 FILLCELL_X4 FILLER_3_620 ();
 FILLCELL_X4 FILLER_3_630 ();
 FILLCELL_X1 FILLER_3_659 ();
 FILLCELL_X1 FILLER_3_664 ();
 FILLCELL_X4 FILLER_3_673 ();
 FILLCELL_X2 FILLER_3_677 ();
 FILLCELL_X1 FILLER_3_679 ();
 FILLCELL_X4 FILLER_3_690 ();
 FILLCELL_X4 FILLER_3_715 ();
 FILLCELL_X2 FILLER_3_723 ();
 FILLCELL_X1 FILLER_3_739 ();
 FILLCELL_X4 FILLER_3_744 ();
 FILLCELL_X2 FILLER_3_768 ();
 FILLCELL_X1 FILLER_3_770 ();
 FILLCELL_X32 FILLER_3_795 ();
 FILLCELL_X32 FILLER_3_827 ();
 FILLCELL_X32 FILLER_3_859 ();
 FILLCELL_X32 FILLER_3_891 ();
 FILLCELL_X32 FILLER_3_923 ();
 FILLCELL_X16 FILLER_3_955 ();
 FILLCELL_X8 FILLER_3_971 ();
 FILLCELL_X2 FILLER_3_979 ();
 FILLCELL_X1 FILLER_3_981 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X4 FILLER_4_65 ();
 FILLCELL_X2 FILLER_4_69 ();
 FILLCELL_X16 FILLER_4_77 ();
 FILLCELL_X8 FILLER_4_93 ();
 FILLCELL_X4 FILLER_4_101 ();
 FILLCELL_X1 FILLER_4_105 ();
 FILLCELL_X8 FILLER_4_115 ();
 FILLCELL_X1 FILLER_4_123 ();
 FILLCELL_X8 FILLER_4_132 ();
 FILLCELL_X4 FILLER_4_140 ();
 FILLCELL_X2 FILLER_4_144 ();
 FILLCELL_X4 FILLER_4_149 ();
 FILLCELL_X2 FILLER_4_153 ();
 FILLCELL_X8 FILLER_4_169 ();
 FILLCELL_X4 FILLER_4_177 ();
 FILLCELL_X4 FILLER_4_210 ();
 FILLCELL_X2 FILLER_4_217 ();
 FILLCELL_X16 FILLER_4_224 ();
 FILLCELL_X8 FILLER_4_240 ();
 FILLCELL_X4 FILLER_4_248 ();
 FILLCELL_X2 FILLER_4_252 ();
 FILLCELL_X4 FILLER_4_283 ();
 FILLCELL_X1 FILLER_4_287 ();
 FILLCELL_X8 FILLER_4_311 ();
 FILLCELL_X4 FILLER_4_319 ();
 FILLCELL_X1 FILLER_4_323 ();
 FILLCELL_X8 FILLER_4_338 ();
 FILLCELL_X1 FILLER_4_346 ();
 FILLCELL_X8 FILLER_4_356 ();
 FILLCELL_X2 FILLER_4_364 ();
 FILLCELL_X16 FILLER_4_375 ();
 FILLCELL_X4 FILLER_4_391 ();
 FILLCELL_X2 FILLER_4_395 ();
 FILLCELL_X2 FILLER_4_415 ();
 FILLCELL_X1 FILLER_4_417 ();
 FILLCELL_X32 FILLER_4_428 ();
 FILLCELL_X8 FILLER_4_460 ();
 FILLCELL_X2 FILLER_4_468 ();
 FILLCELL_X1 FILLER_4_470 ();
 FILLCELL_X8 FILLER_4_473 ();
 FILLCELL_X4 FILLER_4_493 ();
 FILLCELL_X1 FILLER_4_497 ();
 FILLCELL_X2 FILLER_4_508 ();
 FILLCELL_X1 FILLER_4_510 ();
 FILLCELL_X2 FILLER_4_517 ();
 FILLCELL_X8 FILLER_4_525 ();
 FILLCELL_X4 FILLER_4_533 ();
 FILLCELL_X1 FILLER_4_537 ();
 FILLCELL_X8 FILLER_4_563 ();
 FILLCELL_X2 FILLER_4_571 ();
 FILLCELL_X16 FILLER_4_600 ();
 FILLCELL_X8 FILLER_4_616 ();
 FILLCELL_X4 FILLER_4_624 ();
 FILLCELL_X2 FILLER_4_628 ();
 FILLCELL_X1 FILLER_4_630 ();
 FILLCELL_X2 FILLER_4_652 ();
 FILLCELL_X1 FILLER_4_654 ();
 FILLCELL_X32 FILLER_4_677 ();
 FILLCELL_X4 FILLER_4_709 ();
 FILLCELL_X2 FILLER_4_713 ();
 FILLCELL_X4 FILLER_4_728 ();
 FILLCELL_X2 FILLER_4_732 ();
 FILLCELL_X1 FILLER_4_734 ();
 FILLCELL_X1 FILLER_4_754 ();
 FILLCELL_X8 FILLER_4_761 ();
 FILLCELL_X4 FILLER_4_769 ();
 FILLCELL_X2 FILLER_4_780 ();
 FILLCELL_X32 FILLER_4_792 ();
 FILLCELL_X32 FILLER_4_824 ();
 FILLCELL_X32 FILLER_4_856 ();
 FILLCELL_X32 FILLER_4_888 ();
 FILLCELL_X32 FILLER_4_920 ();
 FILLCELL_X16 FILLER_4_952 ();
 FILLCELL_X8 FILLER_4_968 ();
 FILLCELL_X4 FILLER_4_976 ();
 FILLCELL_X2 FILLER_4_980 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X16 FILLER_5_33 ();
 FILLCELL_X8 FILLER_5_49 ();
 FILLCELL_X2 FILLER_5_57 ();
 FILLCELL_X4 FILLER_5_63 ();
 FILLCELL_X2 FILLER_5_67 ();
 FILLCELL_X1 FILLER_5_91 ();
 FILLCELL_X1 FILLER_5_101 ();
 FILLCELL_X8 FILLER_5_109 ();
 FILLCELL_X2 FILLER_5_117 ();
 FILLCELL_X2 FILLER_5_129 ();
 FILLCELL_X1 FILLER_5_135 ();
 FILLCELL_X4 FILLER_5_182 ();
 FILLCELL_X2 FILLER_5_194 ();
 FILLCELL_X2 FILLER_5_214 ();
 FILLCELL_X1 FILLER_5_216 ();
 FILLCELL_X32 FILLER_5_221 ();
 FILLCELL_X4 FILLER_5_253 ();
 FILLCELL_X2 FILLER_5_257 ();
 FILLCELL_X1 FILLER_5_259 ();
 FILLCELL_X2 FILLER_5_266 ();
 FILLCELL_X8 FILLER_5_284 ();
 FILLCELL_X2 FILLER_5_292 ();
 FILLCELL_X1 FILLER_5_294 ();
 FILLCELL_X2 FILLER_5_305 ();
 FILLCELL_X1 FILLER_5_307 ();
 FILLCELL_X4 FILLER_5_321 ();
 FILLCELL_X16 FILLER_5_332 ();
 FILLCELL_X8 FILLER_5_348 ();
 FILLCELL_X4 FILLER_5_356 ();
 FILLCELL_X8 FILLER_5_378 ();
 FILLCELL_X2 FILLER_5_386 ();
 FILLCELL_X1 FILLER_5_388 ();
 FILLCELL_X2 FILLER_5_392 ();
 FILLCELL_X8 FILLER_5_397 ();
 FILLCELL_X1 FILLER_5_405 ();
 FILLCELL_X16 FILLER_5_411 ();
 FILLCELL_X8 FILLER_5_427 ();
 FILLCELL_X4 FILLER_5_435 ();
 FILLCELL_X2 FILLER_5_439 ();
 FILLCELL_X4 FILLER_5_443 ();
 FILLCELL_X2 FILLER_5_447 ();
 FILLCELL_X1 FILLER_5_459 ();
 FILLCELL_X8 FILLER_5_483 ();
 FILLCELL_X4 FILLER_5_491 ();
 FILLCELL_X1 FILLER_5_495 ();
 FILLCELL_X1 FILLER_5_500 ();
 FILLCELL_X1 FILLER_5_505 ();
 FILLCELL_X16 FILLER_5_528 ();
 FILLCELL_X8 FILLER_5_544 ();
 FILLCELL_X1 FILLER_5_552 ();
 FILLCELL_X16 FILLER_5_563 ();
 FILLCELL_X4 FILLER_5_579 ();
 FILLCELL_X1 FILLER_5_583 ();
 FILLCELL_X8 FILLER_5_599 ();
 FILLCELL_X4 FILLER_5_607 ();
 FILLCELL_X2 FILLER_5_611 ();
 FILLCELL_X1 FILLER_5_621 ();
 FILLCELL_X2 FILLER_5_626 ();
 FILLCELL_X1 FILLER_5_628 ();
 FILLCELL_X4 FILLER_5_633 ();
 FILLCELL_X1 FILLER_5_637 ();
 FILLCELL_X2 FILLER_5_644 ();
 FILLCELL_X1 FILLER_5_650 ();
 FILLCELL_X2 FILLER_5_662 ();
 FILLCELL_X2 FILLER_5_671 ();
 FILLCELL_X1 FILLER_5_673 ();
 FILLCELL_X4 FILLER_5_682 ();
 FILLCELL_X2 FILLER_5_686 ();
 FILLCELL_X1 FILLER_5_688 ();
 FILLCELL_X2 FILLER_5_702 ();
 FILLCELL_X8 FILLER_5_717 ();
 FILLCELL_X4 FILLER_5_725 ();
 FILLCELL_X1 FILLER_5_729 ();
 FILLCELL_X4 FILLER_5_748 ();
 FILLCELL_X1 FILLER_5_752 ();
 FILLCELL_X4 FILLER_5_758 ();
 FILLCELL_X2 FILLER_5_762 ();
 FILLCELL_X1 FILLER_5_764 ();
 FILLCELL_X32 FILLER_5_792 ();
 FILLCELL_X32 FILLER_5_824 ();
 FILLCELL_X32 FILLER_5_856 ();
 FILLCELL_X32 FILLER_5_888 ();
 FILLCELL_X32 FILLER_5_920 ();
 FILLCELL_X16 FILLER_5_952 ();
 FILLCELL_X8 FILLER_5_968 ();
 FILLCELL_X4 FILLER_5_976 ();
 FILLCELL_X2 FILLER_5_980 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X16 FILLER_6_33 ();
 FILLCELL_X4 FILLER_6_49 ();
 FILLCELL_X2 FILLER_6_53 ();
 FILLCELL_X2 FILLER_6_86 ();
 FILLCELL_X1 FILLER_6_124 ();
 FILLCELL_X8 FILLER_6_134 ();
 FILLCELL_X2 FILLER_6_142 ();
 FILLCELL_X1 FILLER_6_144 ();
 FILLCELL_X1 FILLER_6_180 ();
 FILLCELL_X1 FILLER_6_194 ();
 FILLCELL_X1 FILLER_6_200 ();
 FILLCELL_X1 FILLER_6_210 ();
 FILLCELL_X8 FILLER_6_218 ();
 FILLCELL_X1 FILLER_6_226 ();
 FILLCELL_X4 FILLER_6_232 ();
 FILLCELL_X2 FILLER_6_236 ();
 FILLCELL_X8 FILLER_6_245 ();
 FILLCELL_X4 FILLER_6_253 ();
 FILLCELL_X2 FILLER_6_257 ();
 FILLCELL_X1 FILLER_6_259 ();
 FILLCELL_X2 FILLER_6_266 ();
 FILLCELL_X1 FILLER_6_270 ();
 FILLCELL_X8 FILLER_6_276 ();
 FILLCELL_X2 FILLER_6_284 ();
 FILLCELL_X2 FILLER_6_300 ();
 FILLCELL_X8 FILLER_6_322 ();
 FILLCELL_X2 FILLER_6_330 ();
 FILLCELL_X1 FILLER_6_332 ();
 FILLCELL_X8 FILLER_6_338 ();
 FILLCELL_X4 FILLER_6_346 ();
 FILLCELL_X1 FILLER_6_350 ();
 FILLCELL_X8 FILLER_6_374 ();
 FILLCELL_X2 FILLER_6_382 ();
 FILLCELL_X1 FILLER_6_384 ();
 FILLCELL_X2 FILLER_6_388 ();
 FILLCELL_X8 FILLER_6_402 ();
 FILLCELL_X4 FILLER_6_410 ();
 FILLCELL_X16 FILLER_6_424 ();
 FILLCELL_X8 FILLER_6_440 ();
 FILLCELL_X1 FILLER_6_448 ();
 FILLCELL_X16 FILLER_6_471 ();
 FILLCELL_X8 FILLER_6_487 ();
 FILLCELL_X4 FILLER_6_495 ();
 FILLCELL_X2 FILLER_6_499 ();
 FILLCELL_X1 FILLER_6_501 ();
 FILLCELL_X2 FILLER_6_509 ();
 FILLCELL_X1 FILLER_6_511 ();
 FILLCELL_X16 FILLER_6_525 ();
 FILLCELL_X8 FILLER_6_541 ();
 FILLCELL_X4 FILLER_6_549 ();
 FILLCELL_X1 FILLER_6_553 ();
 FILLCELL_X2 FILLER_6_574 ();
 FILLCELL_X1 FILLER_6_576 ();
 FILLCELL_X1 FILLER_6_598 ();
 FILLCELL_X2 FILLER_6_617 ();
 FILLCELL_X2 FILLER_6_646 ();
 FILLCELL_X1 FILLER_6_648 ();
 FILLCELL_X8 FILLER_6_667 ();
 FILLCELL_X2 FILLER_6_675 ();
 FILLCELL_X4 FILLER_6_707 ();
 FILLCELL_X1 FILLER_6_711 ();
 FILLCELL_X2 FILLER_6_715 ();
 FILLCELL_X1 FILLER_6_717 ();
 FILLCELL_X1 FILLER_6_721 ();
 FILLCELL_X4 FILLER_6_725 ();
 FILLCELL_X2 FILLER_6_729 ();
 FILLCELL_X1 FILLER_6_731 ();
 FILLCELL_X2 FILLER_6_758 ();
 FILLCELL_X8 FILLER_6_777 ();
 FILLCELL_X1 FILLER_6_785 ();
 FILLCELL_X32 FILLER_6_795 ();
 FILLCELL_X32 FILLER_6_827 ();
 FILLCELL_X32 FILLER_6_859 ();
 FILLCELL_X32 FILLER_6_891 ();
 FILLCELL_X32 FILLER_6_923 ();
 FILLCELL_X16 FILLER_6_955 ();
 FILLCELL_X8 FILLER_6_971 ();
 FILLCELL_X2 FILLER_6_979 ();
 FILLCELL_X1 FILLER_6_981 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X16 FILLER_7_33 ();
 FILLCELL_X4 FILLER_7_49 ();
 FILLCELL_X2 FILLER_7_53 ();
 FILLCELL_X2 FILLER_7_92 ();
 FILLCELL_X2 FILLER_7_149 ();
 FILLCELL_X1 FILLER_7_151 ();
 FILLCELL_X8 FILLER_7_161 ();
 FILLCELL_X4 FILLER_7_169 ();
 FILLCELL_X4 FILLER_7_186 ();
 FILLCELL_X2 FILLER_7_190 ();
 FILLCELL_X1 FILLER_7_192 ();
 FILLCELL_X8 FILLER_7_206 ();
 FILLCELL_X4 FILLER_7_214 ();
 FILLCELL_X2 FILLER_7_218 ();
 FILLCELL_X1 FILLER_7_220 ();
 FILLCELL_X8 FILLER_7_252 ();
 FILLCELL_X4 FILLER_7_260 ();
 FILLCELL_X1 FILLER_7_264 ();
 FILLCELL_X2 FILLER_7_300 ();
 FILLCELL_X16 FILLER_7_315 ();
 FILLCELL_X8 FILLER_7_331 ();
 FILLCELL_X4 FILLER_7_339 ();
 FILLCELL_X2 FILLER_7_371 ();
 FILLCELL_X2 FILLER_7_400 ();
 FILLCELL_X1 FILLER_7_411 ();
 FILLCELL_X4 FILLER_7_419 ();
 FILLCELL_X4 FILLER_7_427 ();
 FILLCELL_X1 FILLER_7_431 ();
 FILLCELL_X8 FILLER_7_468 ();
 FILLCELL_X4 FILLER_7_476 ();
 FILLCELL_X4 FILLER_7_489 ();
 FILLCELL_X1 FILLER_7_493 ();
 FILLCELL_X32 FILLER_7_518 ();
 FILLCELL_X32 FILLER_7_550 ();
 FILLCELL_X2 FILLER_7_582 ();
 FILLCELL_X1 FILLER_7_584 ();
 FILLCELL_X2 FILLER_7_589 ();
 FILLCELL_X1 FILLER_7_591 ();
 FILLCELL_X2 FILLER_7_594 ();
 FILLCELL_X4 FILLER_7_612 ();
 FILLCELL_X2 FILLER_7_620 ();
 FILLCELL_X1 FILLER_7_622 ();
 FILLCELL_X8 FILLER_7_643 ();
 FILLCELL_X1 FILLER_7_651 ();
 FILLCELL_X8 FILLER_7_664 ();
 FILLCELL_X2 FILLER_7_672 ();
 FILLCELL_X4 FILLER_7_685 ();
 FILLCELL_X8 FILLER_7_696 ();
 FILLCELL_X4 FILLER_7_704 ();
 FILLCELL_X1 FILLER_7_718 ();
 FILLCELL_X2 FILLER_7_725 ();
 FILLCELL_X1 FILLER_7_747 ();
 FILLCELL_X1 FILLER_7_768 ();
 FILLCELL_X4 FILLER_7_772 ();
 FILLCELL_X2 FILLER_7_776 ();
 FILLCELL_X1 FILLER_7_778 ();
 FILLCELL_X32 FILLER_7_792 ();
 FILLCELL_X32 FILLER_7_824 ();
 FILLCELL_X32 FILLER_7_856 ();
 FILLCELL_X32 FILLER_7_888 ();
 FILLCELL_X32 FILLER_7_920 ();
 FILLCELL_X16 FILLER_7_952 ();
 FILLCELL_X8 FILLER_7_968 ();
 FILLCELL_X4 FILLER_7_976 ();
 FILLCELL_X2 FILLER_7_980 ();
 FILLCELL_X8 FILLER_8_1 ();
 FILLCELL_X4 FILLER_8_9 ();
 FILLCELL_X2 FILLER_8_13 ();
 FILLCELL_X1 FILLER_8_15 ();
 FILLCELL_X8 FILLER_8_23 ();
 FILLCELL_X1 FILLER_8_31 ();
 FILLCELL_X1 FILLER_8_50 ();
 FILLCELL_X2 FILLER_8_55 ();
 FILLCELL_X2 FILLER_8_62 ();
 FILLCELL_X2 FILLER_8_69 ();
 FILLCELL_X1 FILLER_8_71 ();
 FILLCELL_X2 FILLER_8_83 ();
 FILLCELL_X4 FILLER_8_90 ();
 FILLCELL_X2 FILLER_8_94 ();
 FILLCELL_X1 FILLER_8_96 ();
 FILLCELL_X4 FILLER_8_138 ();
 FILLCELL_X2 FILLER_8_142 ();
 FILLCELL_X1 FILLER_8_144 ();
 FILLCELL_X1 FILLER_8_154 ();
 FILLCELL_X1 FILLER_8_179 ();
 FILLCELL_X16 FILLER_8_187 ();
 FILLCELL_X1 FILLER_8_248 ();
 FILLCELL_X4 FILLER_8_256 ();
 FILLCELL_X8 FILLER_8_270 ();
 FILLCELL_X2 FILLER_8_278 ();
 FILLCELL_X1 FILLER_8_280 ();
 FILLCELL_X16 FILLER_8_308 ();
 FILLCELL_X2 FILLER_8_324 ();
 FILLCELL_X1 FILLER_8_326 ();
 FILLCELL_X2 FILLER_8_336 ();
 FILLCELL_X1 FILLER_8_360 ();
 FILLCELL_X1 FILLER_8_381 ();
 FILLCELL_X2 FILLER_8_391 ();
 FILLCELL_X1 FILLER_8_403 ();
 FILLCELL_X1 FILLER_8_416 ();
 FILLCELL_X2 FILLER_8_420 ();
 FILLCELL_X32 FILLER_8_438 ();
 FILLCELL_X16 FILLER_8_470 ();
 FILLCELL_X8 FILLER_8_486 ();
 FILLCELL_X2 FILLER_8_494 ();
 FILLCELL_X16 FILLER_8_518 ();
 FILLCELL_X8 FILLER_8_534 ();
 FILLCELL_X4 FILLER_8_542 ();
 FILLCELL_X2 FILLER_8_546 ();
 FILLCELL_X4 FILLER_8_555 ();
 FILLCELL_X2 FILLER_8_559 ();
 FILLCELL_X4 FILLER_8_573 ();
 FILLCELL_X2 FILLER_8_577 ();
 FILLCELL_X2 FILLER_8_582 ();
 FILLCELL_X4 FILLER_8_597 ();
 FILLCELL_X2 FILLER_8_601 ();
 FILLCELL_X1 FILLER_8_603 ();
 FILLCELL_X16 FILLER_8_613 ();
 FILLCELL_X2 FILLER_8_629 ();
 FILLCELL_X8 FILLER_8_632 ();
 FILLCELL_X4 FILLER_8_640 ();
 FILLCELL_X2 FILLER_8_644 ();
 FILLCELL_X2 FILLER_8_658 ();
 FILLCELL_X8 FILLER_8_665 ();
 FILLCELL_X4 FILLER_8_677 ();
 FILLCELL_X8 FILLER_8_684 ();
 FILLCELL_X4 FILLER_8_692 ();
 FILLCELL_X1 FILLER_8_700 ();
 FILLCELL_X4 FILLER_8_712 ();
 FILLCELL_X2 FILLER_8_716 ();
 FILLCELL_X1 FILLER_8_718 ();
 FILLCELL_X1 FILLER_8_736 ();
 FILLCELL_X32 FILLER_8_791 ();
 FILLCELL_X32 FILLER_8_823 ();
 FILLCELL_X32 FILLER_8_855 ();
 FILLCELL_X32 FILLER_8_887 ();
 FILLCELL_X32 FILLER_8_919 ();
 FILLCELL_X16 FILLER_8_951 ();
 FILLCELL_X8 FILLER_8_967 ();
 FILLCELL_X4 FILLER_8_975 ();
 FILLCELL_X2 FILLER_8_979 ();
 FILLCELL_X1 FILLER_8_981 ();
 FILLCELL_X8 FILLER_9_1 ();
 FILLCELL_X1 FILLER_9_9 ();
 FILLCELL_X1 FILLER_9_13 ();
 FILLCELL_X2 FILLER_9_46 ();
 FILLCELL_X2 FILLER_9_57 ();
 FILLCELL_X4 FILLER_9_76 ();
 FILLCELL_X2 FILLER_9_85 ();
 FILLCELL_X1 FILLER_9_117 ();
 FILLCELL_X16 FILLER_9_131 ();
 FILLCELL_X8 FILLER_9_147 ();
 FILLCELL_X4 FILLER_9_155 ();
 FILLCELL_X1 FILLER_9_159 ();
 FILLCELL_X4 FILLER_9_162 ();
 FILLCELL_X4 FILLER_9_170 ();
 FILLCELL_X1 FILLER_9_174 ();
 FILLCELL_X1 FILLER_9_178 ();
 FILLCELL_X4 FILLER_9_195 ();
 FILLCELL_X2 FILLER_9_199 ();
 FILLCELL_X4 FILLER_9_205 ();
 FILLCELL_X1 FILLER_9_223 ();
 FILLCELL_X16 FILLER_9_231 ();
 FILLCELL_X4 FILLER_9_247 ();
 FILLCELL_X2 FILLER_9_251 ();
 FILLCELL_X1 FILLER_9_253 ();
 FILLCELL_X32 FILLER_9_256 ();
 FILLCELL_X4 FILLER_9_288 ();
 FILLCELL_X1 FILLER_9_292 ();
 FILLCELL_X2 FILLER_9_307 ();
 FILLCELL_X4 FILLER_9_316 ();
 FILLCELL_X2 FILLER_9_333 ();
 FILLCELL_X1 FILLER_9_348 ();
 FILLCELL_X1 FILLER_9_356 ();
 FILLCELL_X1 FILLER_9_361 ();
 FILLCELL_X2 FILLER_9_375 ();
 FILLCELL_X1 FILLER_9_384 ();
 FILLCELL_X1 FILLER_9_390 ();
 FILLCELL_X2 FILLER_9_402 ();
 FILLCELL_X1 FILLER_9_417 ();
 FILLCELL_X2 FILLER_9_424 ();
 FILLCELL_X2 FILLER_9_431 ();
 FILLCELL_X8 FILLER_9_446 ();
 FILLCELL_X2 FILLER_9_454 ();
 FILLCELL_X1 FILLER_9_456 ();
 FILLCELL_X4 FILLER_9_473 ();
 FILLCELL_X1 FILLER_9_477 ();
 FILLCELL_X4 FILLER_9_482 ();
 FILLCELL_X2 FILLER_9_486 ();
 FILLCELL_X1 FILLER_9_488 ();
 FILLCELL_X1 FILLER_9_495 ();
 FILLCELL_X16 FILLER_9_509 ();
 FILLCELL_X8 FILLER_9_525 ();
 FILLCELL_X4 FILLER_9_550 ();
 FILLCELL_X4 FILLER_9_598 ();
 FILLCELL_X1 FILLER_9_602 ();
 FILLCELL_X16 FILLER_9_618 ();
 FILLCELL_X1 FILLER_9_634 ();
 FILLCELL_X1 FILLER_9_657 ();
 FILLCELL_X1 FILLER_9_660 ();
 FILLCELL_X2 FILLER_9_671 ();
 FILLCELL_X4 FILLER_9_680 ();
 FILLCELL_X2 FILLER_9_706 ();
 FILLCELL_X1 FILLER_9_708 ();
 FILLCELL_X1 FILLER_9_734 ();
 FILLCELL_X8 FILLER_9_740 ();
 FILLCELL_X2 FILLER_9_776 ();
 FILLCELL_X1 FILLER_9_796 ();
 FILLCELL_X32 FILLER_9_815 ();
 FILLCELL_X32 FILLER_9_847 ();
 FILLCELL_X32 FILLER_9_879 ();
 FILLCELL_X32 FILLER_9_911 ();
 FILLCELL_X32 FILLER_9_943 ();
 FILLCELL_X4 FILLER_9_975 ();
 FILLCELL_X2 FILLER_9_979 ();
 FILLCELL_X1 FILLER_9_981 ();
 FILLCELL_X8 FILLER_10_1 ();
 FILLCELL_X1 FILLER_10_9 ();
 FILLCELL_X4 FILLER_10_21 ();
 FILLCELL_X2 FILLER_10_25 ();
 FILLCELL_X4 FILLER_10_38 ();
 FILLCELL_X2 FILLER_10_42 ();
 FILLCELL_X1 FILLER_10_44 ();
 FILLCELL_X2 FILLER_10_64 ();
 FILLCELL_X4 FILLER_10_69 ();
 FILLCELL_X1 FILLER_10_119 ();
 FILLCELL_X4 FILLER_10_140 ();
 FILLCELL_X1 FILLER_10_144 ();
 FILLCELL_X1 FILLER_10_189 ();
 FILLCELL_X8 FILLER_10_195 ();
 FILLCELL_X4 FILLER_10_219 ();
 FILLCELL_X2 FILLER_10_223 ();
 FILLCELL_X4 FILLER_10_229 ();
 FILLCELL_X2 FILLER_10_233 ();
 FILLCELL_X1 FILLER_10_263 ();
 FILLCELL_X16 FILLER_10_271 ();
 FILLCELL_X4 FILLER_10_287 ();
 FILLCELL_X1 FILLER_10_291 ();
 FILLCELL_X4 FILLER_10_312 ();
 FILLCELL_X4 FILLER_10_325 ();
 FILLCELL_X2 FILLER_10_329 ();
 FILLCELL_X2 FILLER_10_334 ();
 FILLCELL_X2 FILLER_10_345 ();
 FILLCELL_X1 FILLER_10_347 ();
 FILLCELL_X2 FILLER_10_351 ();
 FILLCELL_X1 FILLER_10_353 ();
 FILLCELL_X1 FILLER_10_357 ();
 FILLCELL_X4 FILLER_10_365 ();
 FILLCELL_X4 FILLER_10_406 ();
 FILLCELL_X2 FILLER_10_413 ();
 FILLCELL_X1 FILLER_10_415 ();
 FILLCELL_X16 FILLER_10_439 ();
 FILLCELL_X4 FILLER_10_474 ();
 FILLCELL_X1 FILLER_10_478 ();
 FILLCELL_X2 FILLER_10_486 ();
 FILLCELL_X2 FILLER_10_491 ();
 FILLCELL_X16 FILLER_10_505 ();
 FILLCELL_X1 FILLER_10_528 ();
 FILLCELL_X2 FILLER_10_541 ();
 FILLCELL_X1 FILLER_10_543 ();
 FILLCELL_X1 FILLER_10_591 ();
 FILLCELL_X2 FILLER_10_618 ();
 FILLCELL_X1 FILLER_10_630 ();
 FILLCELL_X4 FILLER_10_632 ();
 FILLCELL_X2 FILLER_10_640 ();
 FILLCELL_X1 FILLER_10_646 ();
 FILLCELL_X2 FILLER_10_655 ();
 FILLCELL_X2 FILLER_10_660 ();
 FILLCELL_X1 FILLER_10_679 ();
 FILLCELL_X4 FILLER_10_686 ();
 FILLCELL_X1 FILLER_10_690 ();
 FILLCELL_X16 FILLER_10_710 ();
 FILLCELL_X2 FILLER_10_726 ();
 FILLCELL_X1 FILLER_10_731 ();
 FILLCELL_X8 FILLER_10_734 ();
 FILLCELL_X4 FILLER_10_742 ();
 FILLCELL_X1 FILLER_10_746 ();
 FILLCELL_X8 FILLER_10_767 ();
 FILLCELL_X4 FILLER_10_775 ();
 FILLCELL_X1 FILLER_10_779 ();
 FILLCELL_X4 FILLER_10_790 ();
 FILLCELL_X1 FILLER_10_794 ();
 FILLCELL_X2 FILLER_10_804 ();
 FILLCELL_X1 FILLER_10_806 ();
 FILLCELL_X2 FILLER_10_811 ();
 FILLCELL_X32 FILLER_10_818 ();
 FILLCELL_X32 FILLER_10_850 ();
 FILLCELL_X32 FILLER_10_882 ();
 FILLCELL_X32 FILLER_10_914 ();
 FILLCELL_X32 FILLER_10_946 ();
 FILLCELL_X4 FILLER_10_978 ();
 FILLCELL_X8 FILLER_11_1 ();
 FILLCELL_X2 FILLER_11_9 ();
 FILLCELL_X4 FILLER_11_35 ();
 FILLCELL_X16 FILLER_11_43 ();
 FILLCELL_X8 FILLER_11_59 ();
 FILLCELL_X8 FILLER_11_90 ();
 FILLCELL_X4 FILLER_11_98 ();
 FILLCELL_X4 FILLER_11_119 ();
 FILLCELL_X1 FILLER_11_123 ();
 FILLCELL_X1 FILLER_11_147 ();
 FILLCELL_X1 FILLER_11_190 ();
 FILLCELL_X1 FILLER_11_253 ();
 FILLCELL_X8 FILLER_11_283 ();
 FILLCELL_X2 FILLER_11_291 ();
 FILLCELL_X1 FILLER_11_293 ();
 FILLCELL_X4 FILLER_11_345 ();
 FILLCELL_X1 FILLER_11_349 ();
 FILLCELL_X4 FILLER_11_376 ();
 FILLCELL_X2 FILLER_11_380 ();
 FILLCELL_X1 FILLER_11_382 ();
 FILLCELL_X32 FILLER_11_393 ();
 FILLCELL_X16 FILLER_11_425 ();
 FILLCELL_X8 FILLER_11_441 ();
 FILLCELL_X2 FILLER_11_449 ();
 FILLCELL_X1 FILLER_11_451 ();
 FILLCELL_X4 FILLER_11_462 ();
 FILLCELL_X2 FILLER_11_466 ();
 FILLCELL_X1 FILLER_11_477 ();
 FILLCELL_X2 FILLER_11_488 ();
 FILLCELL_X1 FILLER_11_490 ();
 FILLCELL_X8 FILLER_11_512 ();
 FILLCELL_X1 FILLER_11_520 ();
 FILLCELL_X1 FILLER_11_526 ();
 FILLCELL_X1 FILLER_11_537 ();
 FILLCELL_X1 FILLER_11_547 ();
 FILLCELL_X1 FILLER_11_564 ();
 FILLCELL_X2 FILLER_11_578 ();
 FILLCELL_X2 FILLER_11_590 ();
 FILLCELL_X1 FILLER_11_592 ();
 FILLCELL_X2 FILLER_11_603 ();
 FILLCELL_X1 FILLER_11_621 ();
 FILLCELL_X8 FILLER_11_638 ();
 FILLCELL_X1 FILLER_11_646 ();
 FILLCELL_X32 FILLER_11_654 ();
 FILLCELL_X1 FILLER_11_686 ();
 FILLCELL_X8 FILLER_11_690 ();
 FILLCELL_X4 FILLER_11_698 ();
 FILLCELL_X4 FILLER_11_705 ();
 FILLCELL_X2 FILLER_11_709 ();
 FILLCELL_X1 FILLER_11_717 ();
 FILLCELL_X4 FILLER_11_742 ();
 FILLCELL_X1 FILLER_11_746 ();
 FILLCELL_X2 FILLER_11_756 ();
 FILLCELL_X1 FILLER_11_758 ();
 FILLCELL_X4 FILLER_11_769 ();
 FILLCELL_X2 FILLER_11_773 ();
 FILLCELL_X32 FILLER_11_830 ();
 FILLCELL_X32 FILLER_11_862 ();
 FILLCELL_X32 FILLER_11_894 ();
 FILLCELL_X32 FILLER_11_926 ();
 FILLCELL_X16 FILLER_11_958 ();
 FILLCELL_X8 FILLER_11_974 ();
 FILLCELL_X8 FILLER_12_1 ();
 FILLCELL_X4 FILLER_12_9 ();
 FILLCELL_X1 FILLER_12_13 ();
 FILLCELL_X32 FILLER_12_26 ();
 FILLCELL_X16 FILLER_12_58 ();
 FILLCELL_X4 FILLER_12_74 ();
 FILLCELL_X2 FILLER_12_78 ();
 FILLCELL_X16 FILLER_12_89 ();
 FILLCELL_X8 FILLER_12_105 ();
 FILLCELL_X4 FILLER_12_113 ();
 FILLCELL_X1 FILLER_12_117 ();
 FILLCELL_X4 FILLER_12_138 ();
 FILLCELL_X1 FILLER_12_142 ();
 FILLCELL_X1 FILLER_12_176 ();
 FILLCELL_X1 FILLER_12_182 ();
 FILLCELL_X1 FILLER_12_194 ();
 FILLCELL_X1 FILLER_12_198 ();
 FILLCELL_X4 FILLER_12_208 ();
 FILLCELL_X2 FILLER_12_219 ();
 FILLCELL_X1 FILLER_12_280 ();
 FILLCELL_X2 FILLER_12_323 ();
 FILLCELL_X4 FILLER_12_375 ();
 FILLCELL_X2 FILLER_12_379 ();
 FILLCELL_X1 FILLER_12_381 ();
 FILLCELL_X16 FILLER_12_386 ();
 FILLCELL_X4 FILLER_12_402 ();
 FILLCELL_X8 FILLER_12_412 ();
 FILLCELL_X4 FILLER_12_420 ();
 FILLCELL_X16 FILLER_12_435 ();
 FILLCELL_X2 FILLER_12_451 ();
 FILLCELL_X1 FILLER_12_456 ();
 FILLCELL_X32 FILLER_12_460 ();
 FILLCELL_X8 FILLER_12_492 ();
 FILLCELL_X2 FILLER_12_534 ();
 FILLCELL_X1 FILLER_12_547 ();
 FILLCELL_X1 FILLER_12_554 ();
 FILLCELL_X16 FILLER_12_567 ();
 FILLCELL_X8 FILLER_12_583 ();
 FILLCELL_X2 FILLER_12_591 ();
 FILLCELL_X4 FILLER_12_598 ();
 FILLCELL_X1 FILLER_12_602 ();
 FILLCELL_X2 FILLER_12_628 ();
 FILLCELL_X1 FILLER_12_630 ();
 FILLCELL_X8 FILLER_12_632 ();
 FILLCELL_X4 FILLER_12_640 ();
 FILLCELL_X2 FILLER_12_644 ();
 FILLCELL_X1 FILLER_12_646 ();
 FILLCELL_X16 FILLER_12_656 ();
 FILLCELL_X2 FILLER_12_672 ();
 FILLCELL_X1 FILLER_12_674 ();
 FILLCELL_X4 FILLER_12_692 ();
 FILLCELL_X1 FILLER_12_696 ();
 FILLCELL_X1 FILLER_12_714 ();
 FILLCELL_X1 FILLER_12_720 ();
 FILLCELL_X2 FILLER_12_744 ();
 FILLCELL_X1 FILLER_12_746 ();
 FILLCELL_X1 FILLER_12_772 ();
 FILLCELL_X1 FILLER_12_821 ();
 FILLCELL_X4 FILLER_12_829 ();
 FILLCELL_X2 FILLER_12_841 ();
 FILLCELL_X1 FILLER_12_843 ();
 FILLCELL_X32 FILLER_12_851 ();
 FILLCELL_X32 FILLER_12_883 ();
 FILLCELL_X32 FILLER_12_915 ();
 FILLCELL_X32 FILLER_12_947 ();
 FILLCELL_X2 FILLER_12_979 ();
 FILLCELL_X1 FILLER_12_981 ();
 FILLCELL_X8 FILLER_13_1 ();
 FILLCELL_X1 FILLER_13_9 ();
 FILLCELL_X1 FILLER_13_17 ();
 FILLCELL_X1 FILLER_13_27 ();
 FILLCELL_X2 FILLER_13_31 ();
 FILLCELL_X2 FILLER_13_38 ();
 FILLCELL_X2 FILLER_13_57 ();
 FILLCELL_X2 FILLER_13_65 ();
 FILLCELL_X1 FILLER_13_67 ();
 FILLCELL_X32 FILLER_13_91 ();
 FILLCELL_X1 FILLER_13_123 ();
 FILLCELL_X16 FILLER_13_127 ();
 FILLCELL_X4 FILLER_13_143 ();
 FILLCELL_X1 FILLER_13_147 ();
 FILLCELL_X2 FILLER_13_158 ();
 FILLCELL_X1 FILLER_13_160 ();
 FILLCELL_X8 FILLER_13_170 ();
 FILLCELL_X4 FILLER_13_178 ();
 FILLCELL_X2 FILLER_13_182 ();
 FILLCELL_X1 FILLER_13_184 ();
 FILLCELL_X2 FILLER_13_198 ();
 FILLCELL_X1 FILLER_13_207 ();
 FILLCELL_X2 FILLER_13_237 ();
 FILLCELL_X1 FILLER_13_239 ();
 FILLCELL_X1 FILLER_13_245 ();
 FILLCELL_X2 FILLER_13_250 ();
 FILLCELL_X1 FILLER_13_252 ();
 FILLCELL_X4 FILLER_13_255 ();
 FILLCELL_X2 FILLER_13_259 ();
 FILLCELL_X2 FILLER_13_270 ();
 FILLCELL_X1 FILLER_13_272 ();
 FILLCELL_X4 FILLER_13_279 ();
 FILLCELL_X2 FILLER_13_283 ();
 FILLCELL_X1 FILLER_13_326 ();
 FILLCELL_X8 FILLER_13_331 ();
 FILLCELL_X1 FILLER_13_339 ();
 FILLCELL_X8 FILLER_13_358 ();
 FILLCELL_X8 FILLER_13_370 ();
 FILLCELL_X2 FILLER_13_378 ();
 FILLCELL_X1 FILLER_13_380 ();
 FILLCELL_X2 FILLER_13_394 ();
 FILLCELL_X1 FILLER_13_396 ();
 FILLCELL_X8 FILLER_13_427 ();
 FILLCELL_X4 FILLER_13_435 ();
 FILLCELL_X2 FILLER_13_439 ();
 FILLCELL_X1 FILLER_13_441 ();
 FILLCELL_X8 FILLER_13_452 ();
 FILLCELL_X2 FILLER_13_460 ();
 FILLCELL_X8 FILLER_13_468 ();
 FILLCELL_X4 FILLER_13_476 ();
 FILLCELL_X2 FILLER_13_480 ();
 FILLCELL_X4 FILLER_13_499 ();
 FILLCELL_X2 FILLER_13_503 ();
 FILLCELL_X1 FILLER_13_505 ();
 FILLCELL_X32 FILLER_13_511 ();
 FILLCELL_X32 FILLER_13_543 ();
 FILLCELL_X16 FILLER_13_575 ();
 FILLCELL_X8 FILLER_13_591 ();
 FILLCELL_X4 FILLER_13_606 ();
 FILLCELL_X4 FILLER_13_618 ();
 FILLCELL_X1 FILLER_13_622 ();
 FILLCELL_X4 FILLER_13_633 ();
 FILLCELL_X2 FILLER_13_637 ();
 FILLCELL_X1 FILLER_13_639 ();
 FILLCELL_X2 FILLER_13_647 ();
 FILLCELL_X4 FILLER_13_662 ();
 FILLCELL_X1 FILLER_13_666 ();
 FILLCELL_X1 FILLER_13_671 ();
 FILLCELL_X1 FILLER_13_677 ();
 FILLCELL_X1 FILLER_13_711 ();
 FILLCELL_X1 FILLER_13_746 ();
 FILLCELL_X8 FILLER_13_766 ();
 FILLCELL_X1 FILLER_13_774 ();
 FILLCELL_X1 FILLER_13_780 ();
 FILLCELL_X2 FILLER_13_790 ();
 FILLCELL_X1 FILLER_13_792 ();
 FILLCELL_X8 FILLER_13_797 ();
 FILLCELL_X1 FILLER_13_805 ();
 FILLCELL_X4 FILLER_13_829 ();
 FILLCELL_X1 FILLER_13_833 ();
 FILLCELL_X32 FILLER_13_852 ();
 FILLCELL_X32 FILLER_13_884 ();
 FILLCELL_X32 FILLER_13_916 ();
 FILLCELL_X32 FILLER_13_948 ();
 FILLCELL_X2 FILLER_13_980 ();
 FILLCELL_X8 FILLER_14_1 ();
 FILLCELL_X2 FILLER_14_9 ();
 FILLCELL_X2 FILLER_14_58 ();
 FILLCELL_X32 FILLER_14_69 ();
 FILLCELL_X16 FILLER_14_101 ();
 FILLCELL_X2 FILLER_14_117 ();
 FILLCELL_X1 FILLER_14_119 ();
 FILLCELL_X2 FILLER_14_129 ();
 FILLCELL_X1 FILLER_14_131 ();
 FILLCELL_X8 FILLER_14_150 ();
 FILLCELL_X4 FILLER_14_158 ();
 FILLCELL_X1 FILLER_14_162 ();
 FILLCELL_X2 FILLER_14_169 ();
 FILLCELL_X8 FILLER_14_178 ();
 FILLCELL_X4 FILLER_14_186 ();
 FILLCELL_X2 FILLER_14_190 ();
 FILLCELL_X1 FILLER_14_192 ();
 FILLCELL_X8 FILLER_14_209 ();
 FILLCELL_X2 FILLER_14_217 ();
 FILLCELL_X4 FILLER_14_235 ();
 FILLCELL_X1 FILLER_14_250 ();
 FILLCELL_X8 FILLER_14_273 ();
 FILLCELL_X4 FILLER_14_281 ();
 FILLCELL_X2 FILLER_14_285 ();
 FILLCELL_X32 FILLER_14_343 ();
 FILLCELL_X1 FILLER_14_375 ();
 FILLCELL_X2 FILLER_14_403 ();
 FILLCELL_X8 FILLER_14_421 ();
 FILLCELL_X2 FILLER_14_429 ();
 FILLCELL_X1 FILLER_14_431 ();
 FILLCELL_X8 FILLER_14_451 ();
 FILLCELL_X1 FILLER_14_459 ();
 FILLCELL_X4 FILLER_14_492 ();
 FILLCELL_X1 FILLER_14_496 ();
 FILLCELL_X32 FILLER_14_507 ();
 FILLCELL_X8 FILLER_14_539 ();
 FILLCELL_X4 FILLER_14_547 ();
 FILLCELL_X2 FILLER_14_567 ();
 FILLCELL_X1 FILLER_14_569 ();
 FILLCELL_X4 FILLER_14_578 ();
 FILLCELL_X8 FILLER_14_586 ();
 FILLCELL_X1 FILLER_14_600 ();
 FILLCELL_X1 FILLER_14_632 ();
 FILLCELL_X1 FILLER_14_648 ();
 FILLCELL_X1 FILLER_14_651 ();
 FILLCELL_X1 FILLER_14_665 ();
 FILLCELL_X2 FILLER_14_669 ();
 FILLCELL_X2 FILLER_14_675 ();
 FILLCELL_X1 FILLER_14_722 ();
 FILLCELL_X2 FILLER_14_730 ();
 FILLCELL_X1 FILLER_14_732 ();
 FILLCELL_X1 FILLER_14_778 ();
 FILLCELL_X1 FILLER_14_782 ();
 FILLCELL_X1 FILLER_14_790 ();
 FILLCELL_X8 FILLER_14_798 ();
 FILLCELL_X4 FILLER_14_806 ();
 FILLCELL_X2 FILLER_14_810 ();
 FILLCELL_X2 FILLER_14_818 ();
 FILLCELL_X1 FILLER_14_820 ();
 FILLCELL_X4 FILLER_14_823 ();
 FILLCELL_X32 FILLER_14_853 ();
 FILLCELL_X32 FILLER_14_885 ();
 FILLCELL_X32 FILLER_14_917 ();
 FILLCELL_X32 FILLER_14_949 ();
 FILLCELL_X1 FILLER_14_981 ();
 FILLCELL_X8 FILLER_15_1 ();
 FILLCELL_X4 FILLER_15_9 ();
 FILLCELL_X2 FILLER_15_13 ();
 FILLCELL_X16 FILLER_15_52 ();
 FILLCELL_X2 FILLER_15_68 ();
 FILLCELL_X16 FILLER_15_82 ();
 FILLCELL_X4 FILLER_15_98 ();
 FILLCELL_X4 FILLER_15_123 ();
 FILLCELL_X4 FILLER_15_130 ();
 FILLCELL_X1 FILLER_15_134 ();
 FILLCELL_X1 FILLER_15_139 ();
 FILLCELL_X2 FILLER_15_152 ();
 FILLCELL_X1 FILLER_15_177 ();
 FILLCELL_X4 FILLER_15_194 ();
 FILLCELL_X2 FILLER_15_198 ();
 FILLCELL_X2 FILLER_15_228 ();
 FILLCELL_X1 FILLER_15_230 ();
 FILLCELL_X4 FILLER_15_250 ();
 FILLCELL_X1 FILLER_15_254 ();
 FILLCELL_X16 FILLER_15_268 ();
 FILLCELL_X4 FILLER_15_284 ();
 FILLCELL_X2 FILLER_15_288 ();
 FILLCELL_X16 FILLER_15_325 ();
 FILLCELL_X2 FILLER_15_341 ();
 FILLCELL_X8 FILLER_15_348 ();
 FILLCELL_X4 FILLER_15_373 ();
 FILLCELL_X4 FILLER_15_384 ();
 FILLCELL_X16 FILLER_15_408 ();
 FILLCELL_X2 FILLER_15_424 ();
 FILLCELL_X8 FILLER_15_438 ();
 FILLCELL_X1 FILLER_15_446 ();
 FILLCELL_X2 FILLER_15_469 ();
 FILLCELL_X1 FILLER_15_471 ();
 FILLCELL_X4 FILLER_15_477 ();
 FILLCELL_X16 FILLER_15_484 ();
 FILLCELL_X8 FILLER_15_500 ();
 FILLCELL_X4 FILLER_15_508 ();
 FILLCELL_X2 FILLER_15_512 ();
 FILLCELL_X1 FILLER_15_514 ();
 FILLCELL_X8 FILLER_15_518 ();
 FILLCELL_X1 FILLER_15_526 ();
 FILLCELL_X1 FILLER_15_532 ();
 FILLCELL_X8 FILLER_15_540 ();
 FILLCELL_X2 FILLER_15_548 ();
 FILLCELL_X4 FILLER_15_563 ();
 FILLCELL_X2 FILLER_15_598 ();
 FILLCELL_X8 FILLER_15_616 ();
 FILLCELL_X2 FILLER_15_624 ();
 FILLCELL_X8 FILLER_15_630 ();
 FILLCELL_X4 FILLER_15_638 ();
 FILLCELL_X1 FILLER_15_642 ();
 FILLCELL_X8 FILLER_15_652 ();
 FILLCELL_X2 FILLER_15_660 ();
 FILLCELL_X2 FILLER_15_680 ();
 FILLCELL_X2 FILLER_15_703 ();
 FILLCELL_X1 FILLER_15_728 ();
 FILLCELL_X1 FILLER_15_746 ();
 FILLCELL_X4 FILLER_15_751 ();
 FILLCELL_X1 FILLER_15_761 ();
 FILLCELL_X2 FILLER_15_768 ();
 FILLCELL_X1 FILLER_15_779 ();
 FILLCELL_X2 FILLER_15_787 ();
 FILLCELL_X16 FILLER_15_803 ();
 FILLCELL_X1 FILLER_15_819 ();
 FILLCELL_X2 FILLER_15_824 ();
 FILLCELL_X1 FILLER_15_826 ();
 FILLCELL_X1 FILLER_15_841 ();
 FILLCELL_X32 FILLER_15_844 ();
 FILLCELL_X32 FILLER_15_876 ();
 FILLCELL_X32 FILLER_15_908 ();
 FILLCELL_X32 FILLER_15_940 ();
 FILLCELL_X8 FILLER_15_972 ();
 FILLCELL_X2 FILLER_15_980 ();
 FILLCELL_X8 FILLER_16_1 ();
 FILLCELL_X2 FILLER_16_9 ();
 FILLCELL_X16 FILLER_16_36 ();
 FILLCELL_X8 FILLER_16_52 ();
 FILLCELL_X4 FILLER_16_60 ();
 FILLCELL_X2 FILLER_16_70 ();
 FILLCELL_X1 FILLER_16_85 ();
 FILLCELL_X1 FILLER_16_105 ();
 FILLCELL_X2 FILLER_16_128 ();
 FILLCELL_X1 FILLER_16_134 ();
 FILLCELL_X16 FILLER_16_143 ();
 FILLCELL_X4 FILLER_16_159 ();
 FILLCELL_X1 FILLER_16_163 ();
 FILLCELL_X16 FILLER_16_187 ();
 FILLCELL_X4 FILLER_16_203 ();
 FILLCELL_X2 FILLER_16_207 ();
 FILLCELL_X1 FILLER_16_234 ();
 FILLCELL_X2 FILLER_16_242 ();
 FILLCELL_X2 FILLER_16_250 ();
 FILLCELL_X1 FILLER_16_263 ();
 FILLCELL_X16 FILLER_16_274 ();
 FILLCELL_X1 FILLER_16_290 ();
 FILLCELL_X1 FILLER_16_306 ();
 FILLCELL_X1 FILLER_16_309 ();
 FILLCELL_X16 FILLER_16_313 ();
 FILLCELL_X4 FILLER_16_329 ();
 FILLCELL_X1 FILLER_16_333 ();
 FILLCELL_X32 FILLER_16_341 ();
 FILLCELL_X2 FILLER_16_373 ();
 FILLCELL_X1 FILLER_16_375 ();
 FILLCELL_X2 FILLER_16_414 ();
 FILLCELL_X1 FILLER_16_416 ();
 FILLCELL_X1 FILLER_16_421 ();
 FILLCELL_X1 FILLER_16_426 ();
 FILLCELL_X1 FILLER_16_431 ();
 FILLCELL_X1 FILLER_16_451 ();
 FILLCELL_X2 FILLER_16_454 ();
 FILLCELL_X2 FILLER_16_481 ();
 FILLCELL_X16 FILLER_16_487 ();
 FILLCELL_X8 FILLER_16_503 ();
 FILLCELL_X2 FILLER_16_511 ();
 FILLCELL_X1 FILLER_16_513 ();
 FILLCELL_X4 FILLER_16_527 ();
 FILLCELL_X2 FILLER_16_560 ();
 FILLCELL_X1 FILLER_16_562 ();
 FILLCELL_X32 FILLER_16_586 ();
 FILLCELL_X8 FILLER_16_618 ();
 FILLCELL_X4 FILLER_16_626 ();
 FILLCELL_X1 FILLER_16_630 ();
 FILLCELL_X32 FILLER_16_632 ();
 FILLCELL_X16 FILLER_16_664 ();
 FILLCELL_X2 FILLER_16_680 ();
 FILLCELL_X2 FILLER_16_686 ();
 FILLCELL_X1 FILLER_16_688 ();
 FILLCELL_X1 FILLER_16_703 ();
 FILLCELL_X4 FILLER_16_717 ();
 FILLCELL_X1 FILLER_16_724 ();
 FILLCELL_X2 FILLER_16_728 ();
 FILLCELL_X1 FILLER_16_730 ();
 FILLCELL_X16 FILLER_16_749 ();
 FILLCELL_X4 FILLER_16_765 ();
 FILLCELL_X1 FILLER_16_769 ();
 FILLCELL_X2 FILLER_16_784 ();
 FILLCELL_X16 FILLER_16_791 ();
 FILLCELL_X8 FILLER_16_807 ();
 FILLCELL_X4 FILLER_16_815 ();
 FILLCELL_X2 FILLER_16_819 ();
 FILLCELL_X1 FILLER_16_830 ();
 FILLCELL_X1 FILLER_16_833 ();
 FILLCELL_X32 FILLER_16_849 ();
 FILLCELL_X32 FILLER_16_881 ();
 FILLCELL_X32 FILLER_16_913 ();
 FILLCELL_X32 FILLER_16_945 ();
 FILLCELL_X4 FILLER_16_977 ();
 FILLCELL_X1 FILLER_16_981 ();
 FILLCELL_X16 FILLER_17_1 ();
 FILLCELL_X8 FILLER_17_17 ();
 FILLCELL_X2 FILLER_17_25 ();
 FILLCELL_X1 FILLER_17_34 ();
 FILLCELL_X4 FILLER_17_53 ();
 FILLCELL_X2 FILLER_17_57 ();
 FILLCELL_X1 FILLER_17_59 ();
 FILLCELL_X2 FILLER_17_67 ();
 FILLCELL_X1 FILLER_17_78 ();
 FILLCELL_X4 FILLER_17_81 ();
 FILLCELL_X1 FILLER_17_91 ();
 FILLCELL_X2 FILLER_17_111 ();
 FILLCELL_X4 FILLER_17_123 ();
 FILLCELL_X2 FILLER_17_127 ();
 FILLCELL_X1 FILLER_17_129 ();
 FILLCELL_X16 FILLER_17_142 ();
 FILLCELL_X1 FILLER_17_158 ();
 FILLCELL_X16 FILLER_17_168 ();
 FILLCELL_X4 FILLER_17_184 ();
 FILLCELL_X16 FILLER_17_190 ();
 FILLCELL_X8 FILLER_17_206 ();
 FILLCELL_X2 FILLER_17_214 ();
 FILLCELL_X1 FILLER_17_219 ();
 FILLCELL_X4 FILLER_17_239 ();
 FILLCELL_X2 FILLER_17_243 ();
 FILLCELL_X4 FILLER_17_268 ();
 FILLCELL_X1 FILLER_17_281 ();
 FILLCELL_X2 FILLER_17_287 ();
 FILLCELL_X1 FILLER_17_289 ();
 FILLCELL_X16 FILLER_17_306 ();
 FILLCELL_X4 FILLER_17_322 ();
 FILLCELL_X2 FILLER_17_326 ();
 FILLCELL_X1 FILLER_17_328 ();
 FILLCELL_X4 FILLER_17_341 ();
 FILLCELL_X1 FILLER_17_345 ();
 FILLCELL_X16 FILLER_17_353 ();
 FILLCELL_X8 FILLER_17_369 ();
 FILLCELL_X2 FILLER_17_377 ();
 FILLCELL_X4 FILLER_17_416 ();
 FILLCELL_X2 FILLER_17_420 ();
 FILLCELL_X16 FILLER_17_438 ();
 FILLCELL_X8 FILLER_17_454 ();
 FILLCELL_X4 FILLER_17_462 ();
 FILLCELL_X8 FILLER_17_470 ();
 FILLCELL_X1 FILLER_17_478 ();
 FILLCELL_X8 FILLER_17_500 ();
 FILLCELL_X8 FILLER_17_535 ();
 FILLCELL_X2 FILLER_17_543 ();
 FILLCELL_X1 FILLER_17_545 ();
 FILLCELL_X1 FILLER_17_550 ();
 FILLCELL_X32 FILLER_17_555 ();
 FILLCELL_X32 FILLER_17_587 ();
 FILLCELL_X16 FILLER_17_619 ();
 FILLCELL_X4 FILLER_17_635 ();
 FILLCELL_X2 FILLER_17_639 ();
 FILLCELL_X1 FILLER_17_641 ();
 FILLCELL_X1 FILLER_17_646 ();
 FILLCELL_X16 FILLER_17_653 ();
 FILLCELL_X2 FILLER_17_669 ();
 FILLCELL_X1 FILLER_17_671 ();
 FILLCELL_X16 FILLER_17_676 ();
 FILLCELL_X1 FILLER_17_692 ();
 FILLCELL_X1 FILLER_17_712 ();
 FILLCELL_X4 FILLER_17_718 ();
 FILLCELL_X2 FILLER_17_732 ();
 FILLCELL_X1 FILLER_17_734 ();
 FILLCELL_X32 FILLER_17_740 ();
 FILLCELL_X2 FILLER_17_772 ();
 FILLCELL_X1 FILLER_17_781 ();
 FILLCELL_X2 FILLER_17_798 ();
 FILLCELL_X1 FILLER_17_800 ();
 FILLCELL_X4 FILLER_17_820 ();
 FILLCELL_X2 FILLER_17_832 ();
 FILLCELL_X32 FILLER_17_846 ();
 FILLCELL_X32 FILLER_17_878 ();
 FILLCELL_X32 FILLER_17_910 ();
 FILLCELL_X32 FILLER_17_942 ();
 FILLCELL_X8 FILLER_17_974 ();
 FILLCELL_X8 FILLER_18_1 ();
 FILLCELL_X8 FILLER_18_19 ();
 FILLCELL_X1 FILLER_18_27 ();
 FILLCELL_X16 FILLER_18_38 ();
 FILLCELL_X8 FILLER_18_54 ();
 FILLCELL_X1 FILLER_18_62 ();
 FILLCELL_X8 FILLER_18_72 ();
 FILLCELL_X4 FILLER_18_80 ();
 FILLCELL_X1 FILLER_18_84 ();
 FILLCELL_X2 FILLER_18_92 ();
 FILLCELL_X4 FILLER_18_118 ();
 FILLCELL_X1 FILLER_18_122 ();
 FILLCELL_X8 FILLER_18_130 ();
 FILLCELL_X4 FILLER_18_138 ();
 FILLCELL_X2 FILLER_18_142 ();
 FILLCELL_X2 FILLER_18_165 ();
 FILLCELL_X1 FILLER_18_167 ();
 FILLCELL_X16 FILLER_18_194 ();
 FILLCELL_X2 FILLER_18_210 ();
 FILLCELL_X2 FILLER_18_236 ();
 FILLCELL_X8 FILLER_18_275 ();
 FILLCELL_X2 FILLER_18_283 ();
 FILLCELL_X1 FILLER_18_285 ();
 FILLCELL_X2 FILLER_18_292 ();
 FILLCELL_X1 FILLER_18_294 ();
 FILLCELL_X32 FILLER_18_302 ();
 FILLCELL_X8 FILLER_18_334 ();
 FILLCELL_X2 FILLER_18_342 ();
 FILLCELL_X1 FILLER_18_344 ();
 FILLCELL_X16 FILLER_18_363 ();
 FILLCELL_X4 FILLER_18_379 ();
 FILLCELL_X1 FILLER_18_383 ();
 FILLCELL_X1 FILLER_18_391 ();
 FILLCELL_X1 FILLER_18_402 ();
 FILLCELL_X1 FILLER_18_406 ();
 FILLCELL_X8 FILLER_18_412 ();
 FILLCELL_X2 FILLER_18_420 ();
 FILLCELL_X1 FILLER_18_422 ();
 FILLCELL_X16 FILLER_18_433 ();
 FILLCELL_X8 FILLER_18_449 ();
 FILLCELL_X2 FILLER_18_457 ();
 FILLCELL_X2 FILLER_18_476 ();
 FILLCELL_X1 FILLER_18_478 ();
 FILLCELL_X16 FILLER_18_486 ();
 FILLCELL_X8 FILLER_18_502 ();
 FILLCELL_X4 FILLER_18_510 ();
 FILLCELL_X2 FILLER_18_514 ();
 FILLCELL_X1 FILLER_18_516 ();
 FILLCELL_X2 FILLER_18_521 ();
 FILLCELL_X8 FILLER_18_533 ();
 FILLCELL_X4 FILLER_18_541 ();
 FILLCELL_X2 FILLER_18_545 ();
 FILLCELL_X1 FILLER_18_547 ();
 FILLCELL_X2 FILLER_18_565 ();
 FILLCELL_X8 FILLER_18_577 ();
 FILLCELL_X2 FILLER_18_585 ();
 FILLCELL_X1 FILLER_18_587 ();
 FILLCELL_X8 FILLER_18_605 ();
 FILLCELL_X1 FILLER_18_613 ();
 FILLCELL_X1 FILLER_18_621 ();
 FILLCELL_X2 FILLER_18_629 ();
 FILLCELL_X1 FILLER_18_640 ();
 FILLCELL_X4 FILLER_18_664 ();
 FILLCELL_X2 FILLER_18_672 ();
 FILLCELL_X16 FILLER_18_700 ();
 FILLCELL_X2 FILLER_18_716 ();
 FILLCELL_X16 FILLER_18_727 ();
 FILLCELL_X4 FILLER_18_743 ();
 FILLCELL_X4 FILLER_18_754 ();
 FILLCELL_X1 FILLER_18_774 ();
 FILLCELL_X4 FILLER_18_782 ();
 FILLCELL_X2 FILLER_18_786 ();
 FILLCELL_X4 FILLER_18_793 ();
 FILLCELL_X1 FILLER_18_797 ();
 FILLCELL_X8 FILLER_18_814 ();
 FILLCELL_X4 FILLER_18_831 ();
 FILLCELL_X1 FILLER_18_835 ();
 FILLCELL_X32 FILLER_18_842 ();
 FILLCELL_X32 FILLER_18_874 ();
 FILLCELL_X32 FILLER_18_906 ();
 FILLCELL_X32 FILLER_18_938 ();
 FILLCELL_X8 FILLER_18_970 ();
 FILLCELL_X4 FILLER_18_978 ();
 FILLCELL_X4 FILLER_19_1 ();
 FILLCELL_X2 FILLER_19_5 ();
 FILLCELL_X1 FILLER_19_13 ();
 FILLCELL_X1 FILLER_19_23 ();
 FILLCELL_X1 FILLER_19_31 ();
 FILLCELL_X1 FILLER_19_35 ();
 FILLCELL_X8 FILLER_19_40 ();
 FILLCELL_X4 FILLER_19_48 ();
 FILLCELL_X1 FILLER_19_52 ();
 FILLCELL_X8 FILLER_19_58 ();
 FILLCELL_X2 FILLER_19_66 ();
 FILLCELL_X32 FILLER_19_78 ();
 FILLCELL_X16 FILLER_19_110 ();
 FILLCELL_X8 FILLER_19_126 ();
 FILLCELL_X4 FILLER_19_134 ();
 FILLCELL_X2 FILLER_19_138 ();
 FILLCELL_X2 FILLER_19_159 ();
 FILLCELL_X1 FILLER_19_161 ();
 FILLCELL_X2 FILLER_19_182 ();
 FILLCELL_X32 FILLER_19_207 ();
 FILLCELL_X4 FILLER_19_239 ();
 FILLCELL_X16 FILLER_19_265 ();
 FILLCELL_X8 FILLER_19_281 ();
 FILLCELL_X2 FILLER_19_289 ();
 FILLCELL_X1 FILLER_19_291 ();
 FILLCELL_X16 FILLER_19_328 ();
 FILLCELL_X4 FILLER_19_344 ();
 FILLCELL_X2 FILLER_19_348 ();
 FILLCELL_X4 FILLER_19_367 ();
 FILLCELL_X4 FILLER_19_380 ();
 FILLCELL_X8 FILLER_19_397 ();
 FILLCELL_X4 FILLER_19_424 ();
 FILLCELL_X2 FILLER_19_428 ();
 FILLCELL_X2 FILLER_19_461 ();
 FILLCELL_X1 FILLER_19_463 ();
 FILLCELL_X8 FILLER_19_467 ();
 FILLCELL_X4 FILLER_19_475 ();
 FILLCELL_X32 FILLER_19_488 ();
 FILLCELL_X8 FILLER_19_520 ();
 FILLCELL_X4 FILLER_19_528 ();
 FILLCELL_X1 FILLER_19_596 ();
 FILLCELL_X1 FILLER_19_620 ();
 FILLCELL_X2 FILLER_19_707 ();
 FILLCELL_X1 FILLER_19_709 ();
 FILLCELL_X4 FILLER_19_733 ();
 FILLCELL_X2 FILLER_19_759 ();
 FILLCELL_X1 FILLER_19_761 ();
 FILLCELL_X2 FILLER_19_784 ();
 FILLCELL_X8 FILLER_19_790 ();
 FILLCELL_X4 FILLER_19_798 ();
 FILLCELL_X2 FILLER_19_802 ();
 FILLCELL_X1 FILLER_19_804 ();
 FILLCELL_X4 FILLER_19_823 ();
 FILLCELL_X32 FILLER_19_845 ();
 FILLCELL_X32 FILLER_19_877 ();
 FILLCELL_X32 FILLER_19_909 ();
 FILLCELL_X32 FILLER_19_941 ();
 FILLCELL_X8 FILLER_19_973 ();
 FILLCELL_X1 FILLER_19_981 ();
 FILLCELL_X8 FILLER_20_1 ();
 FILLCELL_X2 FILLER_20_9 ();
 FILLCELL_X1 FILLER_20_11 ();
 FILLCELL_X2 FILLER_20_30 ();
 FILLCELL_X8 FILLER_20_38 ();
 FILLCELL_X2 FILLER_20_46 ();
 FILLCELL_X2 FILLER_20_64 ();
 FILLCELL_X4 FILLER_20_87 ();
 FILLCELL_X1 FILLER_20_91 ();
 FILLCELL_X2 FILLER_20_102 ();
 FILLCELL_X8 FILLER_20_114 ();
 FILLCELL_X4 FILLER_20_122 ();
 FILLCELL_X1 FILLER_20_126 ();
 FILLCELL_X16 FILLER_20_134 ();
 FILLCELL_X4 FILLER_20_150 ();
 FILLCELL_X32 FILLER_20_199 ();
 FILLCELL_X16 FILLER_20_231 ();
 FILLCELL_X1 FILLER_20_247 ();
 FILLCELL_X2 FILLER_20_253 ();
 FILLCELL_X4 FILLER_20_257 ();
 FILLCELL_X2 FILLER_20_261 ();
 FILLCELL_X1 FILLER_20_263 ();
 FILLCELL_X4 FILLER_20_274 ();
 FILLCELL_X8 FILLER_20_280 ();
 FILLCELL_X1 FILLER_20_288 ();
 FILLCELL_X1 FILLER_20_301 ();
 FILLCELL_X1 FILLER_20_306 ();
 FILLCELL_X8 FILLER_20_326 ();
 FILLCELL_X2 FILLER_20_339 ();
 FILLCELL_X8 FILLER_20_344 ();
 FILLCELL_X1 FILLER_20_359 ();
 FILLCELL_X16 FILLER_20_376 ();
 FILLCELL_X8 FILLER_20_392 ();
 FILLCELL_X4 FILLER_20_400 ();
 FILLCELL_X1 FILLER_20_404 ();
 FILLCELL_X4 FILLER_20_425 ();
 FILLCELL_X1 FILLER_20_429 ();
 FILLCELL_X4 FILLER_20_433 ();
 FILLCELL_X1 FILLER_20_437 ();
 FILLCELL_X16 FILLER_20_441 ();
 FILLCELL_X8 FILLER_20_457 ();
 FILLCELL_X2 FILLER_20_465 ();
 FILLCELL_X4 FILLER_20_474 ();
 FILLCELL_X4 FILLER_20_505 ();
 FILLCELL_X2 FILLER_20_516 ();
 FILLCELL_X1 FILLER_20_543 ();
 FILLCELL_X4 FILLER_20_550 ();
 FILLCELL_X2 FILLER_20_554 ();
 FILLCELL_X4 FILLER_20_563 ();
 FILLCELL_X2 FILLER_20_567 ();
 FILLCELL_X4 FILLER_20_578 ();
 FILLCELL_X1 FILLER_20_582 ();
 FILLCELL_X4 FILLER_20_589 ();
 FILLCELL_X16 FILLER_20_606 ();
 FILLCELL_X2 FILLER_20_622 ();
 FILLCELL_X4 FILLER_20_627 ();
 FILLCELL_X1 FILLER_20_632 ();
 FILLCELL_X2 FILLER_20_653 ();
 FILLCELL_X8 FILLER_20_668 ();
 FILLCELL_X4 FILLER_20_686 ();
 FILLCELL_X2 FILLER_20_690 ();
 FILLCELL_X8 FILLER_20_695 ();
 FILLCELL_X4 FILLER_20_703 ();
 FILLCELL_X1 FILLER_20_749 ();
 FILLCELL_X1 FILLER_20_764 ();
 FILLCELL_X1 FILLER_20_773 ();
 FILLCELL_X16 FILLER_20_781 ();
 FILLCELL_X4 FILLER_20_797 ();
 FILLCELL_X4 FILLER_20_817 ();
 FILLCELL_X2 FILLER_20_821 ();
 FILLCELL_X1 FILLER_20_823 ();
 FILLCELL_X32 FILLER_20_833 ();
 FILLCELL_X32 FILLER_20_865 ();
 FILLCELL_X32 FILLER_20_897 ();
 FILLCELL_X32 FILLER_20_929 ();
 FILLCELL_X16 FILLER_20_961 ();
 FILLCELL_X4 FILLER_20_977 ();
 FILLCELL_X1 FILLER_20_981 ();
 FILLCELL_X8 FILLER_21_1 ();
 FILLCELL_X2 FILLER_21_9 ();
 FILLCELL_X2 FILLER_21_14 ();
 FILLCELL_X16 FILLER_21_22 ();
 FILLCELL_X8 FILLER_21_38 ();
 FILLCELL_X4 FILLER_21_46 ();
 FILLCELL_X1 FILLER_21_50 ();
 FILLCELL_X2 FILLER_21_68 ();
 FILLCELL_X2 FILLER_21_112 ();
 FILLCELL_X1 FILLER_21_114 ();
 FILLCELL_X1 FILLER_21_119 ();
 FILLCELL_X32 FILLER_21_130 ();
 FILLCELL_X32 FILLER_21_162 ();
 FILLCELL_X16 FILLER_21_194 ();
 FILLCELL_X8 FILLER_21_210 ();
 FILLCELL_X2 FILLER_21_218 ();
 FILLCELL_X1 FILLER_21_220 ();
 FILLCELL_X1 FILLER_21_228 ();
 FILLCELL_X8 FILLER_21_250 ();
 FILLCELL_X4 FILLER_21_258 ();
 FILLCELL_X2 FILLER_21_262 ();
 FILLCELL_X2 FILLER_21_267 ();
 FILLCELL_X8 FILLER_21_290 ();
 FILLCELL_X16 FILLER_21_322 ();
 FILLCELL_X1 FILLER_21_338 ();
 FILLCELL_X1 FILLER_21_350 ();
 FILLCELL_X4 FILLER_21_364 ();
 FILLCELL_X1 FILLER_21_378 ();
 FILLCELL_X1 FILLER_21_386 ();
 FILLCELL_X4 FILLER_21_392 ();
 FILLCELL_X2 FILLER_21_396 ();
 FILLCELL_X1 FILLER_21_398 ();
 FILLCELL_X2 FILLER_21_423 ();
 FILLCELL_X1 FILLER_21_440 ();
 FILLCELL_X8 FILLER_21_450 ();
 FILLCELL_X4 FILLER_21_458 ();
 FILLCELL_X2 FILLER_21_462 ();
 FILLCELL_X1 FILLER_21_464 ();
 FILLCELL_X2 FILLER_21_482 ();
 FILLCELL_X8 FILLER_21_486 ();
 FILLCELL_X2 FILLER_21_494 ();
 FILLCELL_X4 FILLER_21_533 ();
 FILLCELL_X2 FILLER_21_537 ();
 FILLCELL_X1 FILLER_21_539 ();
 FILLCELL_X8 FILLER_21_548 ();
 FILLCELL_X4 FILLER_21_556 ();
 FILLCELL_X2 FILLER_21_560 ();
 FILLCELL_X32 FILLER_21_566 ();
 FILLCELL_X8 FILLER_21_598 ();
 FILLCELL_X8 FILLER_21_608 ();
 FILLCELL_X4 FILLER_21_616 ();
 FILLCELL_X16 FILLER_21_622 ();
 FILLCELL_X8 FILLER_21_638 ();
 FILLCELL_X2 FILLER_21_646 ();
 FILLCELL_X2 FILLER_21_650 ();
 FILLCELL_X1 FILLER_21_652 ();
 FILLCELL_X2 FILLER_21_659 ();
 FILLCELL_X1 FILLER_21_661 ();
 FILLCELL_X8 FILLER_21_669 ();
 FILLCELL_X8 FILLER_21_686 ();
 FILLCELL_X2 FILLER_21_694 ();
 FILLCELL_X1 FILLER_21_696 ();
 FILLCELL_X4 FILLER_21_755 ();
 FILLCELL_X4 FILLER_21_806 ();
 FILLCELL_X2 FILLER_21_810 ();
 FILLCELL_X32 FILLER_21_837 ();
 FILLCELL_X32 FILLER_21_869 ();
 FILLCELL_X32 FILLER_21_901 ();
 FILLCELL_X32 FILLER_21_933 ();
 FILLCELL_X16 FILLER_21_965 ();
 FILLCELL_X1 FILLER_21_981 ();
 FILLCELL_X16 FILLER_22_1 ();
 FILLCELL_X2 FILLER_22_17 ();
 FILLCELL_X1 FILLER_22_19 ();
 FILLCELL_X4 FILLER_22_25 ();
 FILLCELL_X1 FILLER_22_29 ();
 FILLCELL_X2 FILLER_22_42 ();
 FILLCELL_X1 FILLER_22_44 ();
 FILLCELL_X8 FILLER_22_67 ();
 FILLCELL_X1 FILLER_22_75 ();
 FILLCELL_X8 FILLER_22_83 ();
 FILLCELL_X2 FILLER_22_91 ();
 FILLCELL_X2 FILLER_22_99 ();
 FILLCELL_X8 FILLER_22_128 ();
 FILLCELL_X4 FILLER_22_136 ();
 FILLCELL_X2 FILLER_22_140 ();
 FILLCELL_X32 FILLER_22_152 ();
 FILLCELL_X16 FILLER_22_184 ();
 FILLCELL_X2 FILLER_22_200 ();
 FILLCELL_X1 FILLER_22_209 ();
 FILLCELL_X1 FILLER_22_212 ();
 FILLCELL_X2 FILLER_22_223 ();
 FILLCELL_X16 FILLER_22_241 ();
 FILLCELL_X1 FILLER_22_269 ();
 FILLCELL_X16 FILLER_22_287 ();
 FILLCELL_X16 FILLER_22_323 ();
 FILLCELL_X2 FILLER_22_415 ();
 FILLCELL_X1 FILLER_22_426 ();
 FILLCELL_X4 FILLER_22_437 ();
 FILLCELL_X2 FILLER_22_441 ();
 FILLCELL_X32 FILLER_22_453 ();
 FILLCELL_X4 FILLER_22_485 ();
 FILLCELL_X1 FILLER_22_489 ();
 FILLCELL_X2 FILLER_22_493 ();
 FILLCELL_X1 FILLER_22_495 ();
 FILLCELL_X32 FILLER_22_513 ();
 FILLCELL_X1 FILLER_22_545 ();
 FILLCELL_X8 FILLER_22_549 ();
 FILLCELL_X4 FILLER_22_583 ();
 FILLCELL_X2 FILLER_22_587 ();
 FILLCELL_X1 FILLER_22_606 ();
 FILLCELL_X2 FILLER_22_629 ();
 FILLCELL_X16 FILLER_22_632 ();
 FILLCELL_X4 FILLER_22_648 ();
 FILLCELL_X8 FILLER_22_662 ();
 FILLCELL_X1 FILLER_22_711 ();
 FILLCELL_X2 FILLER_22_715 ();
 FILLCELL_X4 FILLER_22_738 ();
 FILLCELL_X2 FILLER_22_742 ();
 FILLCELL_X8 FILLER_22_748 ();
 FILLCELL_X4 FILLER_22_756 ();
 FILLCELL_X4 FILLER_22_778 ();
 FILLCELL_X2 FILLER_22_782 ();
 FILLCELL_X1 FILLER_22_784 ();
 FILLCELL_X1 FILLER_22_821 ();
 FILLCELL_X1 FILLER_22_831 ();
 FILLCELL_X32 FILLER_22_839 ();
 FILLCELL_X32 FILLER_22_871 ();
 FILLCELL_X32 FILLER_22_903 ();
 FILLCELL_X32 FILLER_22_935 ();
 FILLCELL_X8 FILLER_22_967 ();
 FILLCELL_X4 FILLER_22_975 ();
 FILLCELL_X2 FILLER_22_979 ();
 FILLCELL_X1 FILLER_22_981 ();
 FILLCELL_X8 FILLER_23_1 ();
 FILLCELL_X4 FILLER_23_9 ();
 FILLCELL_X2 FILLER_23_22 ();
 FILLCELL_X8 FILLER_23_48 ();
 FILLCELL_X16 FILLER_23_61 ();
 FILLCELL_X8 FILLER_23_77 ();
 FILLCELL_X4 FILLER_23_85 ();
 FILLCELL_X1 FILLER_23_89 ();
 FILLCELL_X8 FILLER_23_97 ();
 FILLCELL_X2 FILLER_23_105 ();
 FILLCELL_X4 FILLER_23_114 ();
 FILLCELL_X4 FILLER_23_122 ();
 FILLCELL_X2 FILLER_23_132 ();
 FILLCELL_X1 FILLER_23_144 ();
 FILLCELL_X1 FILLER_23_151 ();
 FILLCELL_X2 FILLER_23_158 ();
 FILLCELL_X4 FILLER_23_166 ();
 FILLCELL_X16 FILLER_23_180 ();
 FILLCELL_X1 FILLER_23_196 ();
 FILLCELL_X1 FILLER_23_226 ();
 FILLCELL_X4 FILLER_23_234 ();
 FILLCELL_X8 FILLER_23_240 ();
 FILLCELL_X1 FILLER_23_248 ();
 FILLCELL_X4 FILLER_23_256 ();
 FILLCELL_X2 FILLER_23_275 ();
 FILLCELL_X8 FILLER_23_290 ();
 FILLCELL_X2 FILLER_23_298 ();
 FILLCELL_X16 FILLER_23_305 ();
 FILLCELL_X2 FILLER_23_321 ();
 FILLCELL_X4 FILLER_23_332 ();
 FILLCELL_X2 FILLER_23_359 ();
 FILLCELL_X1 FILLER_23_368 ();
 FILLCELL_X1 FILLER_23_371 ();
 FILLCELL_X1 FILLER_23_381 ();
 FILLCELL_X8 FILLER_23_416 ();
 FILLCELL_X1 FILLER_23_424 ();
 FILLCELL_X4 FILLER_23_442 ();
 FILLCELL_X2 FILLER_23_446 ();
 FILLCELL_X4 FILLER_23_471 ();
 FILLCELL_X1 FILLER_23_475 ();
 FILLCELL_X2 FILLER_23_485 ();
 FILLCELL_X1 FILLER_23_487 ();
 FILLCELL_X32 FILLER_23_494 ();
 FILLCELL_X16 FILLER_23_526 ();
 FILLCELL_X2 FILLER_23_542 ();
 FILLCELL_X4 FILLER_23_556 ();
 FILLCELL_X1 FILLER_23_560 ();
 FILLCELL_X4 FILLER_23_571 ();
 FILLCELL_X2 FILLER_23_604 ();
 FILLCELL_X1 FILLER_23_606 ();
 FILLCELL_X1 FILLER_23_616 ();
 FILLCELL_X4 FILLER_23_627 ();
 FILLCELL_X2 FILLER_23_631 ();
 FILLCELL_X1 FILLER_23_633 ();
 FILLCELL_X32 FILLER_23_644 ();
 FILLCELL_X1 FILLER_23_676 ();
 FILLCELL_X4 FILLER_23_686 ();
 FILLCELL_X2 FILLER_23_690 ();
 FILLCELL_X1 FILLER_23_692 ();
 FILLCELL_X8 FILLER_23_698 ();
 FILLCELL_X1 FILLER_23_720 ();
 FILLCELL_X8 FILLER_23_724 ();
 FILLCELL_X2 FILLER_23_732 ();
 FILLCELL_X16 FILLER_23_741 ();
 FILLCELL_X2 FILLER_23_757 ();
 FILLCELL_X1 FILLER_23_772 ();
 FILLCELL_X2 FILLER_23_782 ();
 FILLCELL_X2 FILLER_23_822 ();
 FILLCELL_X32 FILLER_23_834 ();
 FILLCELL_X32 FILLER_23_866 ();
 FILLCELL_X32 FILLER_23_898 ();
 FILLCELL_X32 FILLER_23_930 ();
 FILLCELL_X16 FILLER_23_962 ();
 FILLCELL_X4 FILLER_23_978 ();
 FILLCELL_X16 FILLER_24_1 ();
 FILLCELL_X4 FILLER_24_17 ();
 FILLCELL_X1 FILLER_24_21 ();
 FILLCELL_X32 FILLER_24_43 ();
 FILLCELL_X8 FILLER_24_75 ();
 FILLCELL_X2 FILLER_24_83 ();
 FILLCELL_X16 FILLER_24_92 ();
 FILLCELL_X8 FILLER_24_108 ();
 FILLCELL_X4 FILLER_24_116 ();
 FILLCELL_X2 FILLER_24_120 ();
 FILLCELL_X1 FILLER_24_122 ();
 FILLCELL_X8 FILLER_24_130 ();
 FILLCELL_X2 FILLER_24_138 ();
 FILLCELL_X1 FILLER_24_140 ();
 FILLCELL_X2 FILLER_24_162 ();
 FILLCELL_X1 FILLER_24_170 ();
 FILLCELL_X32 FILLER_24_174 ();
 FILLCELL_X4 FILLER_24_206 ();
 FILLCELL_X1 FILLER_24_210 ();
 FILLCELL_X16 FILLER_24_220 ();
 FILLCELL_X8 FILLER_24_236 ();
 FILLCELL_X2 FILLER_24_244 ();
 FILLCELL_X1 FILLER_24_246 ();
 FILLCELL_X1 FILLER_24_254 ();
 FILLCELL_X1 FILLER_24_260 ();
 FILLCELL_X8 FILLER_24_268 ();
 FILLCELL_X4 FILLER_24_276 ();
 FILLCELL_X1 FILLER_24_280 ();
 FILLCELL_X8 FILLER_24_286 ();
 FILLCELL_X4 FILLER_24_294 ();
 FILLCELL_X1 FILLER_24_298 ();
 FILLCELL_X8 FILLER_24_308 ();
 FILLCELL_X1 FILLER_24_316 ();
 FILLCELL_X2 FILLER_24_364 ();
 FILLCELL_X4 FILLER_24_378 ();
 FILLCELL_X8 FILLER_24_386 ();
 FILLCELL_X2 FILLER_24_394 ();
 FILLCELL_X1 FILLER_24_396 ();
 FILLCELL_X4 FILLER_24_434 ();
 FILLCELL_X8 FILLER_24_442 ();
 FILLCELL_X4 FILLER_24_450 ();
 FILLCELL_X1 FILLER_24_454 ();
 FILLCELL_X4 FILLER_24_459 ();
 FILLCELL_X2 FILLER_24_463 ();
 FILLCELL_X1 FILLER_24_465 ();
 FILLCELL_X8 FILLER_24_471 ();
 FILLCELL_X32 FILLER_24_508 ();
 FILLCELL_X16 FILLER_24_540 ();
 FILLCELL_X4 FILLER_24_556 ();
 FILLCELL_X2 FILLER_24_560 ();
 FILLCELL_X8 FILLER_24_569 ();
 FILLCELL_X1 FILLER_24_577 ();
 FILLCELL_X8 FILLER_24_587 ();
 FILLCELL_X2 FILLER_24_595 ();
 FILLCELL_X1 FILLER_24_602 ();
 FILLCELL_X8 FILLER_24_607 ();
 FILLCELL_X4 FILLER_24_615 ();
 FILLCELL_X2 FILLER_24_619 ();
 FILLCELL_X1 FILLER_24_621 ();
 FILLCELL_X4 FILLER_24_627 ();
 FILLCELL_X16 FILLER_24_652 ();
 FILLCELL_X4 FILLER_24_668 ();
 FILLCELL_X1 FILLER_24_672 ();
 FILLCELL_X16 FILLER_24_675 ();
 FILLCELL_X8 FILLER_24_691 ();
 FILLCELL_X1 FILLER_24_699 ();
 FILLCELL_X1 FILLER_24_702 ();
 FILLCELL_X8 FILLER_24_727 ();
 FILLCELL_X1 FILLER_24_735 ();
 FILLCELL_X16 FILLER_24_747 ();
 FILLCELL_X2 FILLER_24_763 ();
 FILLCELL_X1 FILLER_24_765 ();
 FILLCELL_X4 FILLER_24_782 ();
 FILLCELL_X2 FILLER_24_786 ();
 FILLCELL_X4 FILLER_24_792 ();
 FILLCELL_X2 FILLER_24_796 ();
 FILLCELL_X2 FILLER_24_816 ();
 FILLCELL_X1 FILLER_24_818 ();
 FILLCELL_X32 FILLER_24_832 ();
 FILLCELL_X32 FILLER_24_864 ();
 FILLCELL_X32 FILLER_24_896 ();
 FILLCELL_X32 FILLER_24_928 ();
 FILLCELL_X16 FILLER_24_960 ();
 FILLCELL_X4 FILLER_24_976 ();
 FILLCELL_X2 FILLER_24_980 ();
 FILLCELL_X8 FILLER_25_1 ();
 FILLCELL_X4 FILLER_25_9 ();
 FILLCELL_X2 FILLER_25_13 ();
 FILLCELL_X2 FILLER_25_25 ();
 FILLCELL_X1 FILLER_25_29 ();
 FILLCELL_X1 FILLER_25_39 ();
 FILLCELL_X16 FILLER_25_53 ();
 FILLCELL_X2 FILLER_25_69 ();
 FILLCELL_X32 FILLER_25_85 ();
 FILLCELL_X32 FILLER_25_117 ();
 FILLCELL_X2 FILLER_25_149 ();
 FILLCELL_X1 FILLER_25_151 ();
 FILLCELL_X1 FILLER_25_164 ();
 FILLCELL_X16 FILLER_25_172 ();
 FILLCELL_X8 FILLER_25_188 ();
 FILLCELL_X2 FILLER_25_196 ();
 FILLCELL_X1 FILLER_25_198 ();
 FILLCELL_X2 FILLER_25_212 ();
 FILLCELL_X1 FILLER_25_214 ();
 FILLCELL_X4 FILLER_25_220 ();
 FILLCELL_X2 FILLER_25_224 ();
 FILLCELL_X1 FILLER_25_226 ();
 FILLCELL_X2 FILLER_25_255 ();
 FILLCELL_X1 FILLER_25_257 ();
 FILLCELL_X2 FILLER_25_271 ();
 FILLCELL_X1 FILLER_25_277 ();
 FILLCELL_X2 FILLER_25_290 ();
 FILLCELL_X1 FILLER_25_306 ();
 FILLCELL_X2 FILLER_25_317 ();
 FILLCELL_X1 FILLER_25_324 ();
 FILLCELL_X4 FILLER_25_330 ();
 FILLCELL_X2 FILLER_25_334 ();
 FILLCELL_X1 FILLER_25_343 ();
 FILLCELL_X8 FILLER_25_355 ();
 FILLCELL_X4 FILLER_25_363 ();
 FILLCELL_X2 FILLER_25_367 ();
 FILLCELL_X1 FILLER_25_369 ();
 FILLCELL_X16 FILLER_25_388 ();
 FILLCELL_X2 FILLER_25_404 ();
 FILLCELL_X4 FILLER_25_409 ();
 FILLCELL_X2 FILLER_25_413 ();
 FILLCELL_X1 FILLER_25_415 ();
 FILLCELL_X2 FILLER_25_427 ();
 FILLCELL_X4 FILLER_25_444 ();
 FILLCELL_X1 FILLER_25_452 ();
 FILLCELL_X2 FILLER_25_457 ();
 FILLCELL_X1 FILLER_25_459 ();
 FILLCELL_X2 FILLER_25_465 ();
 FILLCELL_X4 FILLER_25_474 ();
 FILLCELL_X2 FILLER_25_478 ();
 FILLCELL_X1 FILLER_25_480 ();
 FILLCELL_X4 FILLER_25_497 ();
 FILLCELL_X32 FILLER_25_507 ();
 FILLCELL_X8 FILLER_25_539 ();
 FILLCELL_X32 FILLER_25_559 ();
 FILLCELL_X32 FILLER_25_591 ();
 FILLCELL_X4 FILLER_25_623 ();
 FILLCELL_X2 FILLER_25_627 ();
 FILLCELL_X8 FILLER_25_633 ();
 FILLCELL_X4 FILLER_25_641 ();
 FILLCELL_X1 FILLER_25_645 ();
 FILLCELL_X2 FILLER_25_657 ();
 FILLCELL_X1 FILLER_25_659 ();
 FILLCELL_X2 FILLER_25_676 ();
 FILLCELL_X1 FILLER_25_678 ();
 FILLCELL_X1 FILLER_25_699 ();
 FILLCELL_X1 FILLER_25_722 ();
 FILLCELL_X2 FILLER_25_727 ();
 FILLCELL_X4 FILLER_25_755 ();
 FILLCELL_X1 FILLER_25_759 ();
 FILLCELL_X16 FILLER_25_785 ();
 FILLCELL_X4 FILLER_25_801 ();
 FILLCELL_X2 FILLER_25_805 ();
 FILLCELL_X1 FILLER_25_807 ();
 FILLCELL_X2 FILLER_25_822 ();
 FILLCELL_X1 FILLER_25_824 ();
 FILLCELL_X32 FILLER_25_832 ();
 FILLCELL_X32 FILLER_25_864 ();
 FILLCELL_X32 FILLER_25_896 ();
 FILLCELL_X32 FILLER_25_928 ();
 FILLCELL_X16 FILLER_25_960 ();
 FILLCELL_X4 FILLER_25_976 ();
 FILLCELL_X2 FILLER_25_980 ();
 FILLCELL_X1 FILLER_26_1 ();
 FILLCELL_X4 FILLER_26_25 ();
 FILLCELL_X2 FILLER_26_36 ();
 FILLCELL_X1 FILLER_26_40 ();
 FILLCELL_X1 FILLER_26_60 ();
 FILLCELL_X4 FILLER_26_64 ();
 FILLCELL_X2 FILLER_26_68 ();
 FILLCELL_X1 FILLER_26_103 ();
 FILLCELL_X1 FILLER_26_106 ();
 FILLCELL_X1 FILLER_26_121 ();
 FILLCELL_X8 FILLER_26_132 ();
 FILLCELL_X2 FILLER_26_140 ();
 FILLCELL_X1 FILLER_26_142 ();
 FILLCELL_X4 FILLER_26_159 ();
 FILLCELL_X1 FILLER_26_163 ();
 FILLCELL_X4 FILLER_26_174 ();
 FILLCELL_X2 FILLER_26_178 ();
 FILLCELL_X1 FILLER_26_180 ();
 FILLCELL_X4 FILLER_26_196 ();
 FILLCELL_X1 FILLER_26_225 ();
 FILLCELL_X8 FILLER_26_233 ();
 FILLCELL_X4 FILLER_26_241 ();
 FILLCELL_X4 FILLER_26_248 ();
 FILLCELL_X2 FILLER_26_252 ();
 FILLCELL_X1 FILLER_26_254 ();
 FILLCELL_X4 FILLER_26_262 ();
 FILLCELL_X2 FILLER_26_266 ();
 FILLCELL_X1 FILLER_26_268 ();
 FILLCELL_X4 FILLER_26_278 ();
 FILLCELL_X1 FILLER_26_282 ();
 FILLCELL_X16 FILLER_26_308 ();
 FILLCELL_X32 FILLER_26_338 ();
 FILLCELL_X8 FILLER_26_370 ();
 FILLCELL_X4 FILLER_26_378 ();
 FILLCELL_X4 FILLER_26_398 ();
 FILLCELL_X1 FILLER_26_402 ();
 FILLCELL_X2 FILLER_26_421 ();
 FILLCELL_X1 FILLER_26_479 ();
 FILLCELL_X32 FILLER_26_500 ();
 FILLCELL_X4 FILLER_26_532 ();
 FILLCELL_X32 FILLER_26_564 ();
 FILLCELL_X32 FILLER_26_596 ();
 FILLCELL_X2 FILLER_26_628 ();
 FILLCELL_X1 FILLER_26_630 ();
 FILLCELL_X16 FILLER_26_632 ();
 FILLCELL_X8 FILLER_26_648 ();
 FILLCELL_X4 FILLER_26_656 ();
 FILLCELL_X16 FILLER_26_675 ();
 FILLCELL_X8 FILLER_26_691 ();
 FILLCELL_X2 FILLER_26_699 ();
 FILLCELL_X1 FILLER_26_701 ();
 FILLCELL_X2 FILLER_26_709 ();
 FILLCELL_X8 FILLER_26_721 ();
 FILLCELL_X2 FILLER_26_729 ();
 FILLCELL_X1 FILLER_26_731 ();
 FILLCELL_X2 FILLER_26_741 ();
 FILLCELL_X4 FILLER_26_789 ();
 FILLCELL_X2 FILLER_26_793 ();
 FILLCELL_X1 FILLER_26_795 ();
 FILLCELL_X32 FILLER_26_833 ();
 FILLCELL_X32 FILLER_26_865 ();
 FILLCELL_X32 FILLER_26_897 ();
 FILLCELL_X32 FILLER_26_929 ();
 FILLCELL_X16 FILLER_26_961 ();
 FILLCELL_X4 FILLER_26_977 ();
 FILLCELL_X1 FILLER_26_981 ();
 FILLCELL_X8 FILLER_27_1 ();
 FILLCELL_X4 FILLER_27_9 ();
 FILLCELL_X2 FILLER_27_13 ();
 FILLCELL_X1 FILLER_27_15 ();
 FILLCELL_X2 FILLER_27_48 ();
 FILLCELL_X1 FILLER_27_57 ();
 FILLCELL_X1 FILLER_27_61 ();
 FILLCELL_X4 FILLER_27_66 ();
 FILLCELL_X1 FILLER_27_70 ();
 FILLCELL_X4 FILLER_27_81 ();
 FILLCELL_X2 FILLER_27_85 ();
 FILLCELL_X1 FILLER_27_104 ();
 FILLCELL_X1 FILLER_27_109 ();
 FILLCELL_X1 FILLER_27_112 ();
 FILLCELL_X1 FILLER_27_119 ();
 FILLCELL_X2 FILLER_27_127 ();
 FILLCELL_X8 FILLER_27_135 ();
 FILLCELL_X4 FILLER_27_143 ();
 FILLCELL_X1 FILLER_27_157 ();
 FILLCELL_X1 FILLER_27_163 ();
 FILLCELL_X1 FILLER_27_171 ();
 FILLCELL_X2 FILLER_27_178 ();
 FILLCELL_X8 FILLER_27_188 ();
 FILLCELL_X2 FILLER_27_196 ();
 FILLCELL_X1 FILLER_27_198 ();
 FILLCELL_X2 FILLER_27_202 ();
 FILLCELL_X1 FILLER_27_204 ();
 FILLCELL_X4 FILLER_27_215 ();
 FILLCELL_X2 FILLER_27_228 ();
 FILLCELL_X32 FILLER_27_234 ();
 FILLCELL_X32 FILLER_27_266 ();
 FILLCELL_X32 FILLER_27_298 ();
 FILLCELL_X16 FILLER_27_330 ();
 FILLCELL_X4 FILLER_27_346 ();
 FILLCELL_X2 FILLER_27_350 ();
 FILLCELL_X32 FILLER_27_361 ();
 FILLCELL_X8 FILLER_27_393 ();
 FILLCELL_X2 FILLER_27_401 ();
 FILLCELL_X1 FILLER_27_403 ();
 FILLCELL_X2 FILLER_27_411 ();
 FILLCELL_X2 FILLER_27_416 ();
 FILLCELL_X2 FILLER_27_424 ();
 FILLCELL_X1 FILLER_27_434 ();
 FILLCELL_X8 FILLER_27_442 ();
 FILLCELL_X4 FILLER_27_450 ();
 FILLCELL_X1 FILLER_27_454 ();
 FILLCELL_X1 FILLER_27_468 ();
 FILLCELL_X16 FILLER_27_475 ();
 FILLCELL_X8 FILLER_27_491 ();
 FILLCELL_X8 FILLER_27_527 ();
 FILLCELL_X2 FILLER_27_535 ();
 FILLCELL_X1 FILLER_27_568 ();
 FILLCELL_X8 FILLER_27_592 ();
 FILLCELL_X4 FILLER_27_622 ();
 FILLCELL_X2 FILLER_27_626 ();
 FILLCELL_X1 FILLER_27_628 ();
 FILLCELL_X32 FILLER_27_646 ();
 FILLCELL_X8 FILLER_27_691 ();
 FILLCELL_X4 FILLER_27_699 ();
 FILLCELL_X2 FILLER_27_703 ();
 FILLCELL_X1 FILLER_27_705 ();
 FILLCELL_X8 FILLER_27_727 ();
 FILLCELL_X4 FILLER_27_735 ();
 FILLCELL_X2 FILLER_27_739 ();
 FILLCELL_X1 FILLER_27_741 ();
 FILLCELL_X2 FILLER_27_758 ();
 FILLCELL_X2 FILLER_27_764 ();
 FILLCELL_X4 FILLER_27_787 ();
 FILLCELL_X2 FILLER_27_791 ();
 FILLCELL_X1 FILLER_27_821 ();
 FILLCELL_X32 FILLER_27_829 ();
 FILLCELL_X32 FILLER_27_861 ();
 FILLCELL_X32 FILLER_27_893 ();
 FILLCELL_X32 FILLER_27_925 ();
 FILLCELL_X16 FILLER_27_957 ();
 FILLCELL_X8 FILLER_27_973 ();
 FILLCELL_X1 FILLER_27_981 ();
 FILLCELL_X4 FILLER_28_1 ();
 FILLCELL_X1 FILLER_28_5 ();
 FILLCELL_X16 FILLER_28_27 ();
 FILLCELL_X4 FILLER_28_43 ();
 FILLCELL_X2 FILLER_28_47 ();
 FILLCELL_X16 FILLER_28_66 ();
 FILLCELL_X2 FILLER_28_123 ();
 FILLCELL_X8 FILLER_28_132 ();
 FILLCELL_X4 FILLER_28_140 ();
 FILLCELL_X1 FILLER_28_144 ();
 FILLCELL_X1 FILLER_28_162 ();
 FILLCELL_X16 FILLER_28_167 ();
 FILLCELL_X8 FILLER_28_183 ();
 FILLCELL_X4 FILLER_28_191 ();
 FILLCELL_X2 FILLER_28_195 ();
 FILLCELL_X2 FILLER_28_210 ();
 FILLCELL_X1 FILLER_28_212 ();
 FILLCELL_X32 FILLER_28_235 ();
 FILLCELL_X8 FILLER_28_267 ();
 FILLCELL_X4 FILLER_28_275 ();
 FILLCELL_X1 FILLER_28_279 ();
 FILLCELL_X2 FILLER_28_282 ();
 FILLCELL_X32 FILLER_28_286 ();
 FILLCELL_X2 FILLER_28_318 ();
 FILLCELL_X8 FILLER_28_332 ();
 FILLCELL_X1 FILLER_28_340 ();
 FILLCELL_X4 FILLER_28_351 ();
 FILLCELL_X16 FILLER_28_368 ();
 FILLCELL_X8 FILLER_28_384 ();
 FILLCELL_X4 FILLER_28_392 ();
 FILLCELL_X1 FILLER_28_396 ();
 FILLCELL_X8 FILLER_28_407 ();
 FILLCELL_X4 FILLER_28_415 ();
 FILLCELL_X1 FILLER_28_419 ();
 FILLCELL_X32 FILLER_28_445 ();
 FILLCELL_X16 FILLER_28_477 ();
 FILLCELL_X8 FILLER_28_493 ();
 FILLCELL_X2 FILLER_28_501 ();
 FILLCELL_X16 FILLER_28_528 ();
 FILLCELL_X1 FILLER_28_549 ();
 FILLCELL_X1 FILLER_28_556 ();
 FILLCELL_X8 FILLER_28_564 ();
 FILLCELL_X2 FILLER_28_572 ();
 FILLCELL_X1 FILLER_28_574 ();
 FILLCELL_X8 FILLER_28_585 ();
 FILLCELL_X4 FILLER_28_593 ();
 FILLCELL_X2 FILLER_28_597 ();
 FILLCELL_X4 FILLER_28_606 ();
 FILLCELL_X1 FILLER_28_610 ();
 FILLCELL_X4 FILLER_28_623 ();
 FILLCELL_X2 FILLER_28_629 ();
 FILLCELL_X4 FILLER_28_632 ();
 FILLCELL_X1 FILLER_28_636 ();
 FILLCELL_X1 FILLER_28_639 ();
 FILLCELL_X1 FILLER_28_653 ();
 FILLCELL_X16 FILLER_28_661 ();
 FILLCELL_X1 FILLER_28_687 ();
 FILLCELL_X2 FILLER_28_703 ();
 FILLCELL_X1 FILLER_28_718 ();
 FILLCELL_X2 FILLER_28_725 ();
 FILLCELL_X1 FILLER_28_727 ();
 FILLCELL_X2 FILLER_28_740 ();
 FILLCELL_X1 FILLER_28_742 ();
 FILLCELL_X4 FILLER_28_785 ();
 FILLCELL_X2 FILLER_28_789 ();
 FILLCELL_X1 FILLER_28_791 ();
 FILLCELL_X4 FILLER_28_796 ();
 FILLCELL_X2 FILLER_28_800 ();
 FILLCELL_X1 FILLER_28_802 ();
 FILLCELL_X2 FILLER_28_824 ();
 FILLCELL_X32 FILLER_28_830 ();
 FILLCELL_X32 FILLER_28_862 ();
 FILLCELL_X32 FILLER_28_894 ();
 FILLCELL_X32 FILLER_28_926 ();
 FILLCELL_X16 FILLER_28_958 ();
 FILLCELL_X8 FILLER_28_974 ();
 FILLCELL_X8 FILLER_29_1 ();
 FILLCELL_X2 FILLER_29_9 ();
 FILLCELL_X8 FILLER_29_15 ();
 FILLCELL_X4 FILLER_29_37 ();
 FILLCELL_X1 FILLER_29_41 ();
 FILLCELL_X4 FILLER_29_61 ();
 FILLCELL_X2 FILLER_29_65 ();
 FILLCELL_X16 FILLER_29_72 ();
 FILLCELL_X16 FILLER_29_99 ();
 FILLCELL_X8 FILLER_29_115 ();
 FILLCELL_X4 FILLER_29_123 ();
 FILLCELL_X2 FILLER_29_127 ();
 FILLCELL_X1 FILLER_29_129 ();
 FILLCELL_X8 FILLER_29_143 ();
 FILLCELL_X1 FILLER_29_151 ();
 FILLCELL_X4 FILLER_29_172 ();
 FILLCELL_X2 FILLER_29_176 ();
 FILLCELL_X1 FILLER_29_178 ();
 FILLCELL_X16 FILLER_29_182 ();
 FILLCELL_X1 FILLER_29_198 ();
 FILLCELL_X4 FILLER_29_206 ();
 FILLCELL_X1 FILLER_29_210 ();
 FILLCELL_X8 FILLER_29_223 ();
 FILLCELL_X4 FILLER_29_231 ();
 FILLCELL_X16 FILLER_29_247 ();
 FILLCELL_X8 FILLER_29_263 ();
 FILLCELL_X2 FILLER_29_271 ();
 FILLCELL_X1 FILLER_29_273 ();
 FILLCELL_X1 FILLER_29_280 ();
 FILLCELL_X1 FILLER_29_285 ();
 FILLCELL_X1 FILLER_29_290 ();
 FILLCELL_X2 FILLER_29_296 ();
 FILLCELL_X8 FILLER_29_308 ();
 FILLCELL_X2 FILLER_29_316 ();
 FILLCELL_X1 FILLER_29_318 ();
 FILLCELL_X8 FILLER_29_336 ();
 FILLCELL_X2 FILLER_29_344 ();
 FILLCELL_X1 FILLER_29_346 ();
 FILLCELL_X16 FILLER_29_371 ();
 FILLCELL_X32 FILLER_29_409 ();
 FILLCELL_X16 FILLER_29_441 ();
 FILLCELL_X8 FILLER_29_457 ();
 FILLCELL_X2 FILLER_29_465 ();
 FILLCELL_X1 FILLER_29_467 ();
 FILLCELL_X16 FILLER_29_480 ();
 FILLCELL_X8 FILLER_29_496 ();
 FILLCELL_X2 FILLER_29_504 ();
 FILLCELL_X1 FILLER_29_506 ();
 FILLCELL_X4 FILLER_29_510 ();
 FILLCELL_X1 FILLER_29_514 ();
 FILLCELL_X4 FILLER_29_535 ();
 FILLCELL_X1 FILLER_29_539 ();
 FILLCELL_X2 FILLER_29_550 ();
 FILLCELL_X2 FILLER_29_556 ();
 FILLCELL_X1 FILLER_29_558 ();
 FILLCELL_X8 FILLER_29_566 ();
 FILLCELL_X2 FILLER_29_578 ();
 FILLCELL_X1 FILLER_29_587 ();
 FILLCELL_X8 FILLER_29_594 ();
 FILLCELL_X1 FILLER_29_602 ();
 FILLCELL_X1 FILLER_29_637 ();
 FILLCELL_X4 FILLER_29_654 ();
 FILLCELL_X16 FILLER_29_664 ();
 FILLCELL_X2 FILLER_29_686 ();
 FILLCELL_X1 FILLER_29_688 ();
 FILLCELL_X4 FILLER_29_707 ();
 FILLCELL_X2 FILLER_29_711 ();
 FILLCELL_X2 FILLER_29_730 ();
 FILLCELL_X4 FILLER_29_736 ();
 FILLCELL_X2 FILLER_29_747 ();
 FILLCELL_X4 FILLER_29_756 ();
 FILLCELL_X4 FILLER_29_765 ();
 FILLCELL_X1 FILLER_29_769 ();
 FILLCELL_X2 FILLER_29_790 ();
 FILLCELL_X2 FILLER_29_799 ();
 FILLCELL_X1 FILLER_29_801 ();
 FILLCELL_X8 FILLER_29_809 ();
 FILLCELL_X1 FILLER_29_817 ();
 FILLCELL_X32 FILLER_29_828 ();
 FILLCELL_X32 FILLER_29_860 ();
 FILLCELL_X32 FILLER_29_892 ();
 FILLCELL_X32 FILLER_29_924 ();
 FILLCELL_X16 FILLER_29_956 ();
 FILLCELL_X8 FILLER_29_972 ();
 FILLCELL_X2 FILLER_29_980 ();
 FILLCELL_X4 FILLER_30_1 ();
 FILLCELL_X1 FILLER_30_12 ();
 FILLCELL_X1 FILLER_30_26 ();
 FILLCELL_X8 FILLER_30_30 ();
 FILLCELL_X4 FILLER_30_59 ();
 FILLCELL_X2 FILLER_30_63 ();
 FILLCELL_X1 FILLER_30_65 ();
 FILLCELL_X2 FILLER_30_72 ();
 FILLCELL_X32 FILLER_30_80 ();
 FILLCELL_X8 FILLER_30_112 ();
 FILLCELL_X1 FILLER_30_120 ();
 FILLCELL_X1 FILLER_30_139 ();
 FILLCELL_X8 FILLER_30_150 ();
 FILLCELL_X8 FILLER_30_161 ();
 FILLCELL_X1 FILLER_30_169 ();
 FILLCELL_X4 FILLER_30_183 ();
 FILLCELL_X8 FILLER_30_191 ();
 FILLCELL_X4 FILLER_30_199 ();
 FILLCELL_X1 FILLER_30_211 ();
 FILLCELL_X2 FILLER_30_221 ();
 FILLCELL_X1 FILLER_30_223 ();
 FILLCELL_X4 FILLER_30_234 ();
 FILLCELL_X8 FILLER_30_253 ();
 FILLCELL_X2 FILLER_30_261 ();
 FILLCELL_X1 FILLER_30_263 ();
 FILLCELL_X1 FILLER_30_284 ();
 FILLCELL_X16 FILLER_30_296 ();
 FILLCELL_X4 FILLER_30_312 ();
 FILLCELL_X1 FILLER_30_316 ();
 FILLCELL_X4 FILLER_30_323 ();
 FILLCELL_X4 FILLER_30_346 ();
 FILLCELL_X1 FILLER_30_359 ();
 FILLCELL_X8 FILLER_30_372 ();
 FILLCELL_X4 FILLER_30_380 ();
 FILLCELL_X2 FILLER_30_384 ();
 FILLCELL_X1 FILLER_30_398 ();
 FILLCELL_X16 FILLER_30_421 ();
 FILLCELL_X8 FILLER_30_437 ();
 FILLCELL_X2 FILLER_30_445 ();
 FILLCELL_X16 FILLER_30_487 ();
 FILLCELL_X4 FILLER_30_503 ();
 FILLCELL_X1 FILLER_30_507 ();
 FILLCELL_X4 FILLER_30_512 ();
 FILLCELL_X8 FILLER_30_534 ();
 FILLCELL_X2 FILLER_30_542 ();
 FILLCELL_X16 FILLER_30_559 ();
 FILLCELL_X1 FILLER_30_577 ();
 FILLCELL_X1 FILLER_30_601 ();
 FILLCELL_X8 FILLER_30_609 ();
 FILLCELL_X1 FILLER_30_617 ();
 FILLCELL_X1 FILLER_30_635 ();
 FILLCELL_X32 FILLER_30_650 ();
 FILLCELL_X2 FILLER_30_682 ();
 FILLCELL_X1 FILLER_30_684 ();
 FILLCELL_X1 FILLER_30_688 ();
 FILLCELL_X4 FILLER_30_702 ();
 FILLCELL_X2 FILLER_30_706 ();
 FILLCELL_X4 FILLER_30_724 ();
 FILLCELL_X8 FILLER_30_735 ();
 FILLCELL_X1 FILLER_30_743 ();
 FILLCELL_X8 FILLER_30_765 ();
 FILLCELL_X4 FILLER_30_773 ();
 FILLCELL_X1 FILLER_30_781 ();
 FILLCELL_X1 FILLER_30_795 ();
 FILLCELL_X1 FILLER_30_801 ();
 FILLCELL_X32 FILLER_30_828 ();
 FILLCELL_X32 FILLER_30_860 ();
 FILLCELL_X32 FILLER_30_892 ();
 FILLCELL_X32 FILLER_30_924 ();
 FILLCELL_X16 FILLER_30_956 ();
 FILLCELL_X8 FILLER_30_972 ();
 FILLCELL_X2 FILLER_30_980 ();
 FILLCELL_X4 FILLER_31_1 ();
 FILLCELL_X1 FILLER_31_5 ();
 FILLCELL_X8 FILLER_31_33 ();
 FILLCELL_X4 FILLER_31_41 ();
 FILLCELL_X2 FILLER_31_45 ();
 FILLCELL_X8 FILLER_31_53 ();
 FILLCELL_X2 FILLER_31_61 ();
 FILLCELL_X1 FILLER_31_63 ();
 FILLCELL_X8 FILLER_31_82 ();
 FILLCELL_X16 FILLER_31_94 ();
 FILLCELL_X8 FILLER_31_110 ();
 FILLCELL_X2 FILLER_31_118 ();
 FILLCELL_X1 FILLER_31_120 ();
 FILLCELL_X1 FILLER_31_138 ();
 FILLCELL_X4 FILLER_31_152 ();
 FILLCELL_X2 FILLER_31_156 ();
 FILLCELL_X1 FILLER_31_158 ();
 FILLCELL_X1 FILLER_31_171 ();
 FILLCELL_X1 FILLER_31_177 ();
 FILLCELL_X4 FILLER_31_183 ();
 FILLCELL_X2 FILLER_31_187 ();
 FILLCELL_X1 FILLER_31_189 ();
 FILLCELL_X16 FILLER_31_192 ();
 FILLCELL_X1 FILLER_31_214 ();
 FILLCELL_X1 FILLER_31_222 ();
 FILLCELL_X2 FILLER_31_245 ();
 FILLCELL_X1 FILLER_31_247 ();
 FILLCELL_X8 FILLER_31_252 ();
 FILLCELL_X2 FILLER_31_260 ();
 FILLCELL_X1 FILLER_31_262 ();
 FILLCELL_X1 FILLER_31_286 ();
 FILLCELL_X4 FILLER_31_305 ();
 FILLCELL_X2 FILLER_31_309 ();
 FILLCELL_X1 FILLER_31_311 ();
 FILLCELL_X8 FILLER_31_338 ();
 FILLCELL_X4 FILLER_31_346 ();
 FILLCELL_X2 FILLER_31_350 ();
 FILLCELL_X16 FILLER_31_368 ();
 FILLCELL_X8 FILLER_31_384 ();
 FILLCELL_X4 FILLER_31_392 ();
 FILLCELL_X2 FILLER_31_396 ();
 FILLCELL_X4 FILLER_31_417 ();
 FILLCELL_X1 FILLER_31_421 ();
 FILLCELL_X4 FILLER_31_429 ();
 FILLCELL_X1 FILLER_31_433 ();
 FILLCELL_X2 FILLER_31_463 ();
 FILLCELL_X1 FILLER_31_473 ();
 FILLCELL_X1 FILLER_31_483 ();
 FILLCELL_X16 FILLER_31_488 ();
 FILLCELL_X4 FILLER_31_504 ();
 FILLCELL_X2 FILLER_31_508 ();
 FILLCELL_X16 FILLER_31_524 ();
 FILLCELL_X8 FILLER_31_540 ();
 FILLCELL_X2 FILLER_31_558 ();
 FILLCELL_X1 FILLER_31_590 ();
 FILLCELL_X32 FILLER_31_598 ();
 FILLCELL_X8 FILLER_31_630 ();
 FILLCELL_X1 FILLER_31_638 ();
 FILLCELL_X16 FILLER_31_660 ();
 FILLCELL_X4 FILLER_31_676 ();
 FILLCELL_X1 FILLER_31_680 ();
 FILLCELL_X16 FILLER_31_683 ();
 FILLCELL_X8 FILLER_31_699 ();
 FILLCELL_X4 FILLER_31_724 ();
 FILLCELL_X2 FILLER_31_728 ();
 FILLCELL_X1 FILLER_31_730 ();
 FILLCELL_X4 FILLER_31_738 ();
 FILLCELL_X2 FILLER_31_742 ();
 FILLCELL_X4 FILLER_31_749 ();
 FILLCELL_X2 FILLER_31_753 ();
 FILLCELL_X1 FILLER_31_777 ();
 FILLCELL_X2 FILLER_31_780 ();
 FILLCELL_X4 FILLER_31_813 ();
 FILLCELL_X1 FILLER_31_817 ();
 FILLCELL_X32 FILLER_31_832 ();
 FILLCELL_X32 FILLER_31_864 ();
 FILLCELL_X32 FILLER_31_896 ();
 FILLCELL_X32 FILLER_31_928 ();
 FILLCELL_X16 FILLER_31_960 ();
 FILLCELL_X4 FILLER_31_976 ();
 FILLCELL_X2 FILLER_31_980 ();
 FILLCELL_X4 FILLER_32_1 ();
 FILLCELL_X8 FILLER_32_35 ();
 FILLCELL_X4 FILLER_32_43 ();
 FILLCELL_X2 FILLER_32_56 ();
 FILLCELL_X16 FILLER_32_69 ();
 FILLCELL_X8 FILLER_32_85 ();
 FILLCELL_X2 FILLER_32_93 ();
 FILLCELL_X1 FILLER_32_122 ();
 FILLCELL_X1 FILLER_32_134 ();
 FILLCELL_X16 FILLER_32_141 ();
 FILLCELL_X1 FILLER_32_157 ();
 FILLCELL_X16 FILLER_32_181 ();
 FILLCELL_X2 FILLER_32_207 ();
 FILLCELL_X2 FILLER_32_216 ();
 FILLCELL_X4 FILLER_32_231 ();
 FILLCELL_X2 FILLER_32_235 ();
 FILLCELL_X1 FILLER_32_242 ();
 FILLCELL_X8 FILLER_32_250 ();
 FILLCELL_X4 FILLER_32_258 ();
 FILLCELL_X16 FILLER_32_281 ();
 FILLCELL_X8 FILLER_32_297 ();
 FILLCELL_X4 FILLER_32_305 ();
 FILLCELL_X2 FILLER_32_309 ();
 FILLCELL_X1 FILLER_32_311 ();
 FILLCELL_X2 FILLER_32_317 ();
 FILLCELL_X1 FILLER_32_319 ();
 FILLCELL_X16 FILLER_32_327 ();
 FILLCELL_X8 FILLER_32_343 ();
 FILLCELL_X32 FILLER_32_371 ();
 FILLCELL_X1 FILLER_32_403 ();
 FILLCELL_X16 FILLER_32_413 ();
 FILLCELL_X4 FILLER_32_429 ();
 FILLCELL_X1 FILLER_32_433 ();
 FILLCELL_X2 FILLER_32_441 ();
 FILLCELL_X1 FILLER_32_443 ();
 FILLCELL_X8 FILLER_32_497 ();
 FILLCELL_X2 FILLER_32_505 ();
 FILLCELL_X16 FILLER_32_537 ();
 FILLCELL_X4 FILLER_32_553 ();
 FILLCELL_X1 FILLER_32_588 ();
 FILLCELL_X4 FILLER_32_595 ();
 FILLCELL_X2 FILLER_32_599 ();
 FILLCELL_X1 FILLER_32_601 ();
 FILLCELL_X4 FILLER_32_612 ();
 FILLCELL_X2 FILLER_32_616 ();
 FILLCELL_X2 FILLER_32_621 ();
 FILLCELL_X4 FILLER_32_626 ();
 FILLCELL_X1 FILLER_32_630 ();
 FILLCELL_X2 FILLER_32_632 ();
 FILLCELL_X4 FILLER_32_666 ();
 FILLCELL_X2 FILLER_32_670 ();
 FILLCELL_X8 FILLER_32_684 ();
 FILLCELL_X4 FILLER_32_692 ();
 FILLCELL_X1 FILLER_32_696 ();
 FILLCELL_X2 FILLER_32_707 ();
 FILLCELL_X8 FILLER_32_732 ();
 FILLCELL_X1 FILLER_32_740 ();
 FILLCELL_X4 FILLER_32_748 ();
 FILLCELL_X4 FILLER_32_759 ();
 FILLCELL_X8 FILLER_32_784 ();
 FILLCELL_X8 FILLER_32_799 ();
 FILLCELL_X4 FILLER_32_807 ();
 FILLCELL_X1 FILLER_32_811 ();
 FILLCELL_X32 FILLER_32_828 ();
 FILLCELL_X32 FILLER_32_860 ();
 FILLCELL_X32 FILLER_32_892 ();
 FILLCELL_X32 FILLER_32_924 ();
 FILLCELL_X16 FILLER_32_956 ();
 FILLCELL_X8 FILLER_32_972 ();
 FILLCELL_X2 FILLER_32_980 ();
 FILLCELL_X4 FILLER_33_1 ();
 FILLCELL_X1 FILLER_33_19 ();
 FILLCELL_X1 FILLER_33_31 ();
 FILLCELL_X2 FILLER_33_36 ();
 FILLCELL_X1 FILLER_33_45 ();
 FILLCELL_X16 FILLER_33_75 ();
 FILLCELL_X2 FILLER_33_91 ();
 FILLCELL_X32 FILLER_33_113 ();
 FILLCELL_X16 FILLER_33_145 ();
 FILLCELL_X1 FILLER_33_161 ();
 FILLCELL_X8 FILLER_33_172 ();
 FILLCELL_X4 FILLER_33_180 ();
 FILLCELL_X32 FILLER_33_201 ();
 FILLCELL_X1 FILLER_33_233 ();
 FILLCELL_X16 FILLER_33_240 ();
 FILLCELL_X2 FILLER_33_256 ();
 FILLCELL_X2 FILLER_33_268 ();
 FILLCELL_X16 FILLER_33_280 ();
 FILLCELL_X8 FILLER_33_296 ();
 FILLCELL_X2 FILLER_33_304 ();
 FILLCELL_X1 FILLER_33_316 ();
 FILLCELL_X4 FILLER_33_334 ();
 FILLCELL_X2 FILLER_33_338 ();
 FILLCELL_X1 FILLER_33_340 ();
 FILLCELL_X8 FILLER_33_368 ();
 FILLCELL_X4 FILLER_33_376 ();
 FILLCELL_X2 FILLER_33_380 ();
 FILLCELL_X1 FILLER_33_382 ();
 FILLCELL_X16 FILLER_33_419 ();
 FILLCELL_X8 FILLER_33_435 ();
 FILLCELL_X4 FILLER_33_454 ();
 FILLCELL_X1 FILLER_33_458 ();
 FILLCELL_X16 FILLER_33_461 ();
 FILLCELL_X8 FILLER_33_477 ();
 FILLCELL_X4 FILLER_33_485 ();
 FILLCELL_X1 FILLER_33_489 ();
 FILLCELL_X8 FILLER_33_497 ();
 FILLCELL_X4 FILLER_33_505 ();
 FILLCELL_X2 FILLER_33_509 ();
 FILLCELL_X16 FILLER_33_536 ();
 FILLCELL_X4 FILLER_33_552 ();
 FILLCELL_X2 FILLER_33_556 ();
 FILLCELL_X8 FILLER_33_560 ();
 FILLCELL_X4 FILLER_33_568 ();
 FILLCELL_X2 FILLER_33_572 ();
 FILLCELL_X2 FILLER_33_580 ();
 FILLCELL_X2 FILLER_33_584 ();
 FILLCELL_X1 FILLER_33_586 ();
 FILLCELL_X8 FILLER_33_592 ();
 FILLCELL_X2 FILLER_33_600 ();
 FILLCELL_X8 FILLER_33_632 ();
 FILLCELL_X2 FILLER_33_640 ();
 FILLCELL_X1 FILLER_33_642 ();
 FILLCELL_X4 FILLER_33_671 ();
 FILLCELL_X1 FILLER_33_675 ();
 FILLCELL_X8 FILLER_33_687 ();
 FILLCELL_X4 FILLER_33_695 ();
 FILLCELL_X1 FILLER_33_699 ();
 FILLCELL_X4 FILLER_33_735 ();
 FILLCELL_X1 FILLER_33_739 ();
 FILLCELL_X1 FILLER_33_766 ();
 FILLCELL_X32 FILLER_33_813 ();
 FILLCELL_X32 FILLER_33_845 ();
 FILLCELL_X32 FILLER_33_877 ();
 FILLCELL_X32 FILLER_33_909 ();
 FILLCELL_X32 FILLER_33_941 ();
 FILLCELL_X8 FILLER_33_973 ();
 FILLCELL_X1 FILLER_33_981 ();
 FILLCELL_X2 FILLER_34_1 ();
 FILLCELL_X1 FILLER_34_45 ();
 FILLCELL_X1 FILLER_34_64 ();
 FILLCELL_X4 FILLER_34_74 ();
 FILLCELL_X1 FILLER_34_78 ();
 FILLCELL_X4 FILLER_34_89 ();
 FILLCELL_X2 FILLER_34_93 ();
 FILLCELL_X2 FILLER_34_97 ();
 FILLCELL_X1 FILLER_34_99 ();
 FILLCELL_X8 FILLER_34_121 ();
 FILLCELL_X16 FILLER_34_167 ();
 FILLCELL_X1 FILLER_34_183 ();
 FILLCELL_X2 FILLER_34_194 ();
 FILLCELL_X1 FILLER_34_196 ();
 FILLCELL_X8 FILLER_34_208 ();
 FILLCELL_X2 FILLER_34_216 ();
 FILLCELL_X1 FILLER_34_218 ();
 FILLCELL_X4 FILLER_34_229 ();
 FILLCELL_X8 FILLER_34_249 ();
 FILLCELL_X2 FILLER_34_257 ();
 FILLCELL_X4 FILLER_34_262 ();
 FILLCELL_X1 FILLER_34_266 ();
 FILLCELL_X16 FILLER_34_291 ();
 FILLCELL_X4 FILLER_34_307 ();
 FILLCELL_X1 FILLER_34_311 ();
 FILLCELL_X8 FILLER_34_333 ();
 FILLCELL_X4 FILLER_34_341 ();
 FILLCELL_X16 FILLER_34_364 ();
 FILLCELL_X8 FILLER_34_380 ();
 FILLCELL_X4 FILLER_34_388 ();
 FILLCELL_X2 FILLER_34_392 ();
 FILLCELL_X1 FILLER_34_394 ();
 FILLCELL_X16 FILLER_34_425 ();
 FILLCELL_X8 FILLER_34_441 ();
 FILLCELL_X4 FILLER_34_449 ();
 FILLCELL_X16 FILLER_34_455 ();
 FILLCELL_X2 FILLER_34_471 ();
 FILLCELL_X8 FILLER_34_483 ();
 FILLCELL_X1 FILLER_34_491 ();
 FILLCELL_X4 FILLER_34_506 ();
 FILLCELL_X4 FILLER_34_513 ();
 FILLCELL_X2 FILLER_34_517 ();
 FILLCELL_X1 FILLER_34_519 ();
 FILLCELL_X32 FILLER_34_542 ();
 FILLCELL_X4 FILLER_34_574 ();
 FILLCELL_X1 FILLER_34_578 ();
 FILLCELL_X2 FILLER_34_586 ();
 FILLCELL_X4 FILLER_34_598 ();
 FILLCELL_X1 FILLER_34_602 ();
 FILLCELL_X1 FILLER_34_616 ();
 FILLCELL_X1 FILLER_34_626 ();
 FILLCELL_X4 FILLER_34_639 ();
 FILLCELL_X2 FILLER_34_643 ();
 FILLCELL_X1 FILLER_34_654 ();
 FILLCELL_X4 FILLER_34_666 ();
 FILLCELL_X2 FILLER_34_670 ();
 FILLCELL_X2 FILLER_34_704 ();
 FILLCELL_X4 FILLER_34_733 ();
 FILLCELL_X2 FILLER_34_737 ();
 FILLCELL_X1 FILLER_34_739 ();
 FILLCELL_X8 FILLER_34_758 ();
 FILLCELL_X1 FILLER_34_766 ();
 FILLCELL_X4 FILLER_34_772 ();
 FILLCELL_X2 FILLER_34_776 ();
 FILLCELL_X4 FILLER_34_782 ();
 FILLCELL_X32 FILLER_34_826 ();
 FILLCELL_X32 FILLER_34_858 ();
 FILLCELL_X32 FILLER_34_890 ();
 FILLCELL_X32 FILLER_34_922 ();
 FILLCELL_X16 FILLER_34_954 ();
 FILLCELL_X8 FILLER_34_970 ();
 FILLCELL_X4 FILLER_34_978 ();
 FILLCELL_X16 FILLER_35_1 ();
 FILLCELL_X2 FILLER_35_17 ();
 FILLCELL_X16 FILLER_35_24 ();
 FILLCELL_X1 FILLER_35_40 ();
 FILLCELL_X1 FILLER_35_59 ();
 FILLCELL_X16 FILLER_35_112 ();
 FILLCELL_X4 FILLER_35_128 ();
 FILLCELL_X1 FILLER_35_132 ();
 FILLCELL_X2 FILLER_35_136 ();
 FILLCELL_X1 FILLER_35_138 ();
 FILLCELL_X32 FILLER_35_150 ();
 FILLCELL_X2 FILLER_35_182 ();
 FILLCELL_X1 FILLER_35_184 ();
 FILLCELL_X8 FILLER_35_200 ();
 FILLCELL_X4 FILLER_35_208 ();
 FILLCELL_X2 FILLER_35_212 ();
 FILLCELL_X1 FILLER_35_214 ();
 FILLCELL_X2 FILLER_35_222 ();
 FILLCELL_X1 FILLER_35_224 ();
 FILLCELL_X8 FILLER_35_243 ();
 FILLCELL_X2 FILLER_35_251 ();
 FILLCELL_X1 FILLER_35_253 ();
 FILLCELL_X1 FILLER_35_271 ();
 FILLCELL_X16 FILLER_35_278 ();
 FILLCELL_X4 FILLER_35_294 ();
 FILLCELL_X2 FILLER_35_298 ();
 FILLCELL_X1 FILLER_35_300 ();
 FILLCELL_X8 FILLER_35_311 ();
 FILLCELL_X16 FILLER_35_325 ();
 FILLCELL_X4 FILLER_35_341 ();
 FILLCELL_X2 FILLER_35_345 ();
 FILLCELL_X1 FILLER_35_347 ();
 FILLCELL_X16 FILLER_35_370 ();
 FILLCELL_X8 FILLER_35_386 ();
 FILLCELL_X4 FILLER_35_394 ();
 FILLCELL_X2 FILLER_35_403 ();
 FILLCELL_X1 FILLER_35_405 ();
 FILLCELL_X16 FILLER_35_415 ();
 FILLCELL_X8 FILLER_35_431 ();
 FILLCELL_X2 FILLER_35_439 ();
 FILLCELL_X1 FILLER_35_441 ();
 FILLCELL_X1 FILLER_35_456 ();
 FILLCELL_X1 FILLER_35_460 ();
 FILLCELL_X1 FILLER_35_465 ();
 FILLCELL_X8 FILLER_35_470 ();
 FILLCELL_X4 FILLER_35_478 ();
 FILLCELL_X2 FILLER_35_482 ();
 FILLCELL_X2 FILLER_35_496 ();
 FILLCELL_X2 FILLER_35_501 ();
 FILLCELL_X16 FILLER_35_515 ();
 FILLCELL_X8 FILLER_35_531 ();
 FILLCELL_X2 FILLER_35_539 ();
 FILLCELL_X1 FILLER_35_541 ();
 FILLCELL_X8 FILLER_35_564 ();
 FILLCELL_X2 FILLER_35_572 ();
 FILLCELL_X1 FILLER_35_574 ();
 FILLCELL_X4 FILLER_35_585 ();
 FILLCELL_X1 FILLER_35_589 ();
 FILLCELL_X1 FILLER_35_604 ();
 FILLCELL_X1 FILLER_35_609 ();
 FILLCELL_X1 FILLER_35_615 ();
 FILLCELL_X16 FILLER_35_623 ();
 FILLCELL_X8 FILLER_35_639 ();
 FILLCELL_X4 FILLER_35_647 ();
 FILLCELL_X1 FILLER_35_651 ();
 FILLCELL_X4 FILLER_35_659 ();
 FILLCELL_X2 FILLER_35_663 ();
 FILLCELL_X1 FILLER_35_668 ();
 FILLCELL_X8 FILLER_35_683 ();
 FILLCELL_X4 FILLER_35_691 ();
 FILLCELL_X2 FILLER_35_695 ();
 FILLCELL_X8 FILLER_35_729 ();
 FILLCELL_X2 FILLER_35_737 ();
 FILLCELL_X1 FILLER_35_739 ();
 FILLCELL_X1 FILLER_35_749 ();
 FILLCELL_X1 FILLER_35_757 ();
 FILLCELL_X1 FILLER_35_764 ();
 FILLCELL_X1 FILLER_35_774 ();
 FILLCELL_X1 FILLER_35_788 ();
 FILLCELL_X2 FILLER_35_812 ();
 FILLCELL_X1 FILLER_35_814 ();
 FILLCELL_X32 FILLER_35_832 ();
 FILLCELL_X32 FILLER_35_864 ();
 FILLCELL_X32 FILLER_35_896 ();
 FILLCELL_X32 FILLER_35_928 ();
 FILLCELL_X16 FILLER_35_960 ();
 FILLCELL_X4 FILLER_35_976 ();
 FILLCELL_X2 FILLER_35_980 ();
 FILLCELL_X1 FILLER_36_1 ();
 FILLCELL_X16 FILLER_36_12 ();
 FILLCELL_X8 FILLER_36_28 ();
 FILLCELL_X4 FILLER_36_36 ();
 FILLCELL_X1 FILLER_36_40 ();
 FILLCELL_X8 FILLER_36_45 ();
 FILLCELL_X4 FILLER_36_53 ();
 FILLCELL_X2 FILLER_36_57 ();
 FILLCELL_X32 FILLER_36_62 ();
 FILLCELL_X1 FILLER_36_94 ();
 FILLCELL_X16 FILLER_36_104 ();
 FILLCELL_X2 FILLER_36_120 ();
 FILLCELL_X1 FILLER_36_122 ();
 FILLCELL_X2 FILLER_36_136 ();
 FILLCELL_X1 FILLER_36_138 ();
 FILLCELL_X2 FILLER_36_146 ();
 FILLCELL_X16 FILLER_36_155 ();
 FILLCELL_X2 FILLER_36_171 ();
 FILLCELL_X1 FILLER_36_173 ();
 FILLCELL_X2 FILLER_36_184 ();
 FILLCELL_X1 FILLER_36_186 ();
 FILLCELL_X4 FILLER_36_191 ();
 FILLCELL_X2 FILLER_36_195 ();
 FILLCELL_X16 FILLER_36_204 ();
 FILLCELL_X2 FILLER_36_232 ();
 FILLCELL_X1 FILLER_36_234 ();
 FILLCELL_X8 FILLER_36_246 ();
 FILLCELL_X2 FILLER_36_254 ();
 FILLCELL_X8 FILLER_36_303 ();
 FILLCELL_X1 FILLER_36_324 ();
 FILLCELL_X8 FILLER_36_332 ();
 FILLCELL_X2 FILLER_36_340 ();
 FILLCELL_X2 FILLER_36_359 ();
 FILLCELL_X1 FILLER_36_361 ();
 FILLCELL_X8 FILLER_36_387 ();
 FILLCELL_X2 FILLER_36_395 ();
 FILLCELL_X1 FILLER_36_397 ();
 FILLCELL_X8 FILLER_36_409 ();
 FILLCELL_X4 FILLER_36_417 ();
 FILLCELL_X2 FILLER_36_421 ();
 FILLCELL_X8 FILLER_36_435 ();
 FILLCELL_X2 FILLER_36_443 ();
 FILLCELL_X2 FILLER_36_452 ();
 FILLCELL_X4 FILLER_36_456 ();
 FILLCELL_X2 FILLER_36_460 ();
 FILLCELL_X2 FILLER_36_466 ();
 FILLCELL_X1 FILLER_36_468 ();
 FILLCELL_X2 FILLER_36_471 ();
 FILLCELL_X8 FILLER_36_479 ();
 FILLCELL_X4 FILLER_36_487 ();
 FILLCELL_X32 FILLER_36_495 ();
 FILLCELL_X4 FILLER_36_527 ();
 FILLCELL_X1 FILLER_36_531 ();
 FILLCELL_X2 FILLER_36_541 ();
 FILLCELL_X1 FILLER_36_543 ();
 FILLCELL_X16 FILLER_36_562 ();
 FILLCELL_X8 FILLER_36_578 ();
 FILLCELL_X2 FILLER_36_586 ();
 FILLCELL_X1 FILLER_36_588 ();
 FILLCELL_X8 FILLER_36_618 ();
 FILLCELL_X4 FILLER_36_626 ();
 FILLCELL_X1 FILLER_36_630 ();
 FILLCELL_X16 FILLER_36_632 ();
 FILLCELL_X8 FILLER_36_648 ();
 FILLCELL_X2 FILLER_36_656 ();
 FILLCELL_X8 FILLER_36_682 ();
 FILLCELL_X4 FILLER_36_690 ();
 FILLCELL_X1 FILLER_36_694 ();
 FILLCELL_X2 FILLER_36_718 ();
 FILLCELL_X1 FILLER_36_720 ();
 FILLCELL_X4 FILLER_36_725 ();
 FILLCELL_X1 FILLER_36_729 ();
 FILLCELL_X2 FILLER_36_743 ();
 FILLCELL_X1 FILLER_36_758 ();
 FILLCELL_X1 FILLER_36_766 ();
 FILLCELL_X1 FILLER_36_785 ();
 FILLCELL_X2 FILLER_36_803 ();
 FILLCELL_X1 FILLER_36_808 ();
 FILLCELL_X2 FILLER_36_814 ();
 FILLCELL_X4 FILLER_36_829 ();
 FILLCELL_X32 FILLER_36_838 ();
 FILLCELL_X32 FILLER_36_870 ();
 FILLCELL_X32 FILLER_36_902 ();
 FILLCELL_X32 FILLER_36_934 ();
 FILLCELL_X16 FILLER_36_966 ();
 FILLCELL_X4 FILLER_37_1 ();
 FILLCELL_X2 FILLER_37_5 ();
 FILLCELL_X1 FILLER_37_7 ();
 FILLCELL_X4 FILLER_37_21 ();
 FILLCELL_X2 FILLER_37_25 ();
 FILLCELL_X1 FILLER_37_27 ();
 FILLCELL_X4 FILLER_37_53 ();
 FILLCELL_X2 FILLER_37_57 ();
 FILLCELL_X32 FILLER_37_73 ();
 FILLCELL_X2 FILLER_37_105 ();
 FILLCELL_X8 FILLER_37_114 ();
 FILLCELL_X1 FILLER_37_122 ();
 FILLCELL_X1 FILLER_37_126 ();
 FILLCELL_X8 FILLER_37_132 ();
 FILLCELL_X8 FILLER_37_168 ();
 FILLCELL_X1 FILLER_37_176 ();
 FILLCELL_X1 FILLER_37_185 ();
 FILLCELL_X16 FILLER_37_189 ();
 FILLCELL_X8 FILLER_37_205 ();
 FILLCELL_X4 FILLER_37_213 ();
 FILLCELL_X2 FILLER_37_217 ();
 FILLCELL_X1 FILLER_37_219 ();
 FILLCELL_X16 FILLER_37_236 ();
 FILLCELL_X4 FILLER_37_252 ();
 FILLCELL_X2 FILLER_37_256 ();
 FILLCELL_X16 FILLER_37_264 ();
 FILLCELL_X2 FILLER_37_280 ();
 FILLCELL_X1 FILLER_37_282 ();
 FILLCELL_X8 FILLER_37_290 ();
 FILLCELL_X16 FILLER_37_307 ();
 FILLCELL_X4 FILLER_37_323 ();
 FILLCELL_X16 FILLER_37_331 ();
 FILLCELL_X1 FILLER_37_351 ();
 FILLCELL_X16 FILLER_37_374 ();
 FILLCELL_X1 FILLER_37_390 ();
 FILLCELL_X1 FILLER_37_412 ();
 FILLCELL_X16 FILLER_37_420 ();
 FILLCELL_X8 FILLER_37_436 ();
 FILLCELL_X1 FILLER_37_444 ();
 FILLCELL_X4 FILLER_37_447 ();
 FILLCELL_X1 FILLER_37_451 ();
 FILLCELL_X4 FILLER_37_458 ();
 FILLCELL_X1 FILLER_37_462 ();
 FILLCELL_X2 FILLER_37_480 ();
 FILLCELL_X4 FILLER_37_484 ();
 FILLCELL_X1 FILLER_37_501 ();
 FILLCELL_X2 FILLER_37_505 ();
 FILLCELL_X1 FILLER_37_507 ();
 FILLCELL_X8 FILLER_37_512 ();
 FILLCELL_X8 FILLER_37_534 ();
 FILLCELL_X4 FILLER_37_542 ();
 FILLCELL_X2 FILLER_37_546 ();
 FILLCELL_X16 FILLER_37_571 ();
 FILLCELL_X4 FILLER_37_587 ();
 FILLCELL_X2 FILLER_37_607 ();
 FILLCELL_X1 FILLER_37_609 ();
 FILLCELL_X4 FILLER_37_623 ();
 FILLCELL_X2 FILLER_37_627 ();
 FILLCELL_X8 FILLER_37_633 ();
 FILLCELL_X16 FILLER_37_647 ();
 FILLCELL_X4 FILLER_37_663 ();
 FILLCELL_X2 FILLER_37_667 ();
 FILLCELL_X2 FILLER_37_679 ();
 FILLCELL_X8 FILLER_37_691 ();
 FILLCELL_X4 FILLER_37_699 ();
 FILLCELL_X1 FILLER_37_703 ();
 FILLCELL_X1 FILLER_37_708 ();
 FILLCELL_X4 FILLER_37_721 ();
 FILLCELL_X2 FILLER_37_725 ();
 FILLCELL_X4 FILLER_37_734 ();
 FILLCELL_X1 FILLER_37_774 ();
 FILLCELL_X4 FILLER_37_793 ();
 FILLCELL_X2 FILLER_37_797 ();
 FILLCELL_X2 FILLER_37_819 ();
 FILLCELL_X1 FILLER_37_821 ();
 FILLCELL_X32 FILLER_37_832 ();
 FILLCELL_X32 FILLER_37_864 ();
 FILLCELL_X32 FILLER_37_896 ();
 FILLCELL_X32 FILLER_37_928 ();
 FILLCELL_X16 FILLER_37_960 ();
 FILLCELL_X4 FILLER_37_976 ();
 FILLCELL_X2 FILLER_37_980 ();
 FILLCELL_X8 FILLER_38_1 ();
 FILLCELL_X4 FILLER_38_9 ();
 FILLCELL_X1 FILLER_38_13 ();
 FILLCELL_X2 FILLER_38_20 ();
 FILLCELL_X1 FILLER_38_22 ();
 FILLCELL_X1 FILLER_38_50 ();
 FILLCELL_X8 FILLER_38_65 ();
 FILLCELL_X1 FILLER_38_73 ();
 FILLCELL_X16 FILLER_38_80 ();
 FILLCELL_X4 FILLER_38_96 ();
 FILLCELL_X2 FILLER_38_100 ();
 FILLCELL_X1 FILLER_38_102 ();
 FILLCELL_X4 FILLER_38_106 ();
 FILLCELL_X1 FILLER_38_126 ();
 FILLCELL_X1 FILLER_38_131 ();
 FILLCELL_X2 FILLER_38_137 ();
 FILLCELL_X1 FILLER_38_139 ();
 FILLCELL_X2 FILLER_38_167 ();
 FILLCELL_X1 FILLER_38_169 ();
 FILLCELL_X2 FILLER_38_186 ();
 FILLCELL_X8 FILLER_38_201 ();
 FILLCELL_X2 FILLER_38_242 ();
 FILLCELL_X1 FILLER_38_244 ();
 FILLCELL_X8 FILLER_38_247 ();
 FILLCELL_X1 FILLER_38_260 ();
 FILLCELL_X8 FILLER_38_272 ();
 FILLCELL_X4 FILLER_38_286 ();
 FILLCELL_X1 FILLER_38_290 ();
 FILLCELL_X2 FILLER_38_317 ();
 FILLCELL_X1 FILLER_38_319 ();
 FILLCELL_X16 FILLER_38_332 ();
 FILLCELL_X2 FILLER_38_352 ();
 FILLCELL_X1 FILLER_38_354 ();
 FILLCELL_X8 FILLER_38_368 ();
 FILLCELL_X2 FILLER_38_376 ();
 FILLCELL_X8 FILLER_38_381 ();
 FILLCELL_X2 FILLER_38_389 ();
 FILLCELL_X1 FILLER_38_391 ();
 FILLCELL_X4 FILLER_38_412 ();
 FILLCELL_X2 FILLER_38_416 ();
 FILLCELL_X1 FILLER_38_418 ();
 FILLCELL_X1 FILLER_38_421 ();
 FILLCELL_X4 FILLER_38_437 ();
 FILLCELL_X2 FILLER_38_441 ();
 FILLCELL_X1 FILLER_38_443 ();
 FILLCELL_X1 FILLER_38_457 ();
 FILLCELL_X1 FILLER_38_477 ();
 FILLCELL_X1 FILLER_38_491 ();
 FILLCELL_X4 FILLER_38_495 ();
 FILLCELL_X1 FILLER_38_499 ();
 FILLCELL_X4 FILLER_38_513 ();
 FILLCELL_X2 FILLER_38_517 ();
 FILLCELL_X1 FILLER_38_519 ();
 FILLCELL_X4 FILLER_38_550 ();
 FILLCELL_X2 FILLER_38_554 ();
 FILLCELL_X16 FILLER_38_569 ();
 FILLCELL_X4 FILLER_38_585 ();
 FILLCELL_X1 FILLER_38_589 ();
 FILLCELL_X16 FILLER_38_608 ();
 FILLCELL_X4 FILLER_38_624 ();
 FILLCELL_X2 FILLER_38_628 ();
 FILLCELL_X1 FILLER_38_630 ();
 FILLCELL_X8 FILLER_38_632 ();
 FILLCELL_X4 FILLER_38_640 ();
 FILLCELL_X1 FILLER_38_644 ();
 FILLCELL_X2 FILLER_38_649 ();
 FILLCELL_X1 FILLER_38_651 ();
 FILLCELL_X1 FILLER_38_656 ();
 FILLCELL_X8 FILLER_38_661 ();
 FILLCELL_X1 FILLER_38_669 ();
 FILLCELL_X2 FILLER_38_673 ();
 FILLCELL_X2 FILLER_38_680 ();
 FILLCELL_X1 FILLER_38_682 ();
 FILLCELL_X1 FILLER_38_693 ();
 FILLCELL_X4 FILLER_38_732 ();
 FILLCELL_X2 FILLER_38_736 ();
 FILLCELL_X1 FILLER_38_738 ();
 FILLCELL_X1 FILLER_38_757 ();
 FILLCELL_X8 FILLER_38_765 ();
 FILLCELL_X2 FILLER_38_773 ();
 FILLCELL_X1 FILLER_38_775 ();
 FILLCELL_X1 FILLER_38_781 ();
 FILLCELL_X2 FILLER_38_799 ();
 FILLCELL_X1 FILLER_38_801 ();
 FILLCELL_X32 FILLER_38_828 ();
 FILLCELL_X32 FILLER_38_860 ();
 FILLCELL_X32 FILLER_38_892 ();
 FILLCELL_X32 FILLER_38_924 ();
 FILLCELL_X16 FILLER_38_956 ();
 FILLCELL_X8 FILLER_38_972 ();
 FILLCELL_X2 FILLER_38_980 ();
 FILLCELL_X1 FILLER_39_18 ();
 FILLCELL_X8 FILLER_39_29 ();
 FILLCELL_X4 FILLER_39_69 ();
 FILLCELL_X2 FILLER_39_76 ();
 FILLCELL_X8 FILLER_39_87 ();
 FILLCELL_X1 FILLER_39_95 ();
 FILLCELL_X32 FILLER_39_101 ();
 FILLCELL_X8 FILLER_39_133 ();
 FILLCELL_X4 FILLER_39_141 ();
 FILLCELL_X2 FILLER_39_145 ();
 FILLCELL_X1 FILLER_39_147 ();
 FILLCELL_X8 FILLER_39_162 ();
 FILLCELL_X4 FILLER_39_170 ();
 FILLCELL_X2 FILLER_39_174 ();
 FILLCELL_X1 FILLER_39_176 ();
 FILLCELL_X16 FILLER_39_185 ();
 FILLCELL_X4 FILLER_39_201 ();
 FILLCELL_X1 FILLER_39_205 ();
 FILLCELL_X4 FILLER_39_210 ();
 FILLCELL_X2 FILLER_39_214 ();
 FILLCELL_X2 FILLER_39_242 ();
 FILLCELL_X1 FILLER_39_244 ();
 FILLCELL_X2 FILLER_39_252 ();
 FILLCELL_X4 FILLER_39_267 ();
 FILLCELL_X1 FILLER_39_271 ();
 FILLCELL_X2 FILLER_39_288 ();
 FILLCELL_X4 FILLER_39_307 ();
 FILLCELL_X4 FILLER_39_324 ();
 FILLCELL_X8 FILLER_39_335 ();
 FILLCELL_X4 FILLER_39_355 ();
 FILLCELL_X1 FILLER_39_359 ();
 FILLCELL_X16 FILLER_39_369 ();
 FILLCELL_X8 FILLER_39_385 ();
 FILLCELL_X4 FILLER_39_393 ();
 FILLCELL_X1 FILLER_39_397 ();
 FILLCELL_X2 FILLER_39_402 ();
 FILLCELL_X1 FILLER_39_404 ();
 FILLCELL_X1 FILLER_39_436 ();
 FILLCELL_X1 FILLER_39_444 ();
 FILLCELL_X2 FILLER_39_457 ();
 FILLCELL_X1 FILLER_39_459 ();
 FILLCELL_X2 FILLER_39_467 ();
 FILLCELL_X1 FILLER_39_478 ();
 FILLCELL_X1 FILLER_39_483 ();
 FILLCELL_X4 FILLER_39_492 ();
 FILLCELL_X2 FILLER_39_496 ();
 FILLCELL_X1 FILLER_39_498 ();
 FILLCELL_X2 FILLER_39_530 ();
 FILLCELL_X16 FILLER_39_536 ();
 FILLCELL_X4 FILLER_39_552 ();
 FILLCELL_X1 FILLER_39_556 ();
 FILLCELL_X2 FILLER_39_571 ();
 FILLCELL_X8 FILLER_39_577 ();
 FILLCELL_X1 FILLER_39_585 ();
 FILLCELL_X4 FILLER_39_588 ();
 FILLCELL_X2 FILLER_39_609 ();
 FILLCELL_X1 FILLER_39_611 ();
 FILLCELL_X16 FILLER_39_621 ();
 FILLCELL_X2 FILLER_39_637 ();
 FILLCELL_X1 FILLER_39_639 ();
 FILLCELL_X32 FILLER_39_653 ();
 FILLCELL_X2 FILLER_39_685 ();
 FILLCELL_X8 FILLER_39_690 ();
 FILLCELL_X1 FILLER_39_698 ();
 FILLCELL_X4 FILLER_39_706 ();
 FILLCELL_X1 FILLER_39_714 ();
 FILLCELL_X8 FILLER_39_722 ();
 FILLCELL_X1 FILLER_39_739 ();
 FILLCELL_X2 FILLER_39_753 ();
 FILLCELL_X2 FILLER_39_760 ();
 FILLCELL_X16 FILLER_39_776 ();
 FILLCELL_X4 FILLER_39_792 ();
 FILLCELL_X2 FILLER_39_796 ();
 FILLCELL_X1 FILLER_39_801 ();
 FILLCELL_X2 FILLER_39_823 ();
 FILLCELL_X32 FILLER_39_832 ();
 FILLCELL_X32 FILLER_39_864 ();
 FILLCELL_X32 FILLER_39_896 ();
 FILLCELL_X32 FILLER_39_928 ();
 FILLCELL_X16 FILLER_39_960 ();
 FILLCELL_X4 FILLER_39_976 ();
 FILLCELL_X2 FILLER_39_980 ();
 FILLCELL_X4 FILLER_40_1 ();
 FILLCELL_X2 FILLER_40_5 ();
 FILLCELL_X1 FILLER_40_7 ();
 FILLCELL_X1 FILLER_40_11 ();
 FILLCELL_X2 FILLER_40_15 ();
 FILLCELL_X1 FILLER_40_17 ();
 FILLCELL_X1 FILLER_40_23 ();
 FILLCELL_X4 FILLER_40_31 ();
 FILLCELL_X2 FILLER_40_35 ();
 FILLCELL_X1 FILLER_40_71 ();
 FILLCELL_X16 FILLER_40_94 ();
 FILLCELL_X16 FILLER_40_133 ();
 FILLCELL_X2 FILLER_40_149 ();
 FILLCELL_X4 FILLER_40_169 ();
 FILLCELL_X1 FILLER_40_173 ();
 FILLCELL_X4 FILLER_40_182 ();
 FILLCELL_X2 FILLER_40_186 ();
 FILLCELL_X1 FILLER_40_208 ();
 FILLCELL_X2 FILLER_40_239 ();
 FILLCELL_X1 FILLER_40_241 ();
 FILLCELL_X1 FILLER_40_252 ();
 FILLCELL_X1 FILLER_40_257 ();
 FILLCELL_X1 FILLER_40_279 ();
 FILLCELL_X1 FILLER_40_329 ();
 FILLCELL_X2 FILLER_40_333 ();
 FILLCELL_X1 FILLER_40_335 ();
 FILLCELL_X32 FILLER_40_343 ();
 FILLCELL_X1 FILLER_40_375 ();
 FILLCELL_X1 FILLER_40_380 ();
 FILLCELL_X1 FILLER_40_391 ();
 FILLCELL_X1 FILLER_40_396 ();
 FILLCELL_X1 FILLER_40_403 ();
 FILLCELL_X8 FILLER_40_411 ();
 FILLCELL_X4 FILLER_40_419 ();
 FILLCELL_X1 FILLER_40_423 ();
 FILLCELL_X16 FILLER_40_428 ();
 FILLCELL_X4 FILLER_40_444 ();
 FILLCELL_X2 FILLER_40_448 ();
 FILLCELL_X16 FILLER_40_455 ();
 FILLCELL_X1 FILLER_40_471 ();
 FILLCELL_X2 FILLER_40_476 ();
 FILLCELL_X8 FILLER_40_497 ();
 FILLCELL_X2 FILLER_40_505 ();
 FILLCELL_X1 FILLER_40_507 ();
 FILLCELL_X4 FILLER_40_526 ();
 FILLCELL_X8 FILLER_40_542 ();
 FILLCELL_X2 FILLER_40_550 ();
 FILLCELL_X8 FILLER_40_579 ();
 FILLCELL_X16 FILLER_40_610 ();
 FILLCELL_X2 FILLER_40_626 ();
 FILLCELL_X1 FILLER_40_630 ();
 FILLCELL_X1 FILLER_40_632 ();
 FILLCELL_X16 FILLER_40_642 ();
 FILLCELL_X4 FILLER_40_658 ();
 FILLCELL_X2 FILLER_40_662 ();
 FILLCELL_X4 FILLER_40_674 ();
 FILLCELL_X2 FILLER_40_678 ();
 FILLCELL_X4 FILLER_40_723 ();
 FILLCELL_X1 FILLER_40_727 ();
 FILLCELL_X1 FILLER_40_786 ();
 FILLCELL_X4 FILLER_40_800 ();
 FILLCELL_X32 FILLER_40_822 ();
 FILLCELL_X32 FILLER_40_854 ();
 FILLCELL_X32 FILLER_40_886 ();
 FILLCELL_X32 FILLER_40_918 ();
 FILLCELL_X32 FILLER_40_950 ();
 FILLCELL_X8 FILLER_41_1 ();
 FILLCELL_X8 FILLER_41_16 ();
 FILLCELL_X4 FILLER_41_24 ();
 FILLCELL_X1 FILLER_41_41 ();
 FILLCELL_X1 FILLER_41_63 ();
 FILLCELL_X1 FILLER_41_73 ();
 FILLCELL_X1 FILLER_41_83 ();
 FILLCELL_X8 FILLER_41_102 ();
 FILLCELL_X2 FILLER_41_110 ();
 FILLCELL_X8 FILLER_41_155 ();
 FILLCELL_X4 FILLER_41_163 ();
 FILLCELL_X2 FILLER_41_167 ();
 FILLCELL_X32 FILLER_41_194 ();
 FILLCELL_X32 FILLER_41_226 ();
 FILLCELL_X8 FILLER_41_258 ();
 FILLCELL_X1 FILLER_41_266 ();
 FILLCELL_X4 FILLER_41_276 ();
 FILLCELL_X8 FILLER_41_312 ();
 FILLCELL_X4 FILLER_41_320 ();
 FILLCELL_X2 FILLER_41_324 ();
 FILLCELL_X8 FILLER_41_340 ();
 FILLCELL_X2 FILLER_41_348 ();
 FILLCELL_X1 FILLER_41_350 ();
 FILLCELL_X4 FILLER_41_360 ();
 FILLCELL_X1 FILLER_41_373 ();
 FILLCELL_X1 FILLER_41_388 ();
 FILLCELL_X1 FILLER_41_392 ();
 FILLCELL_X2 FILLER_41_423 ();
 FILLCELL_X16 FILLER_41_430 ();
 FILLCELL_X2 FILLER_41_446 ();
 FILLCELL_X8 FILLER_41_457 ();
 FILLCELL_X1 FILLER_41_465 ();
 FILLCELL_X1 FILLER_41_485 ();
 FILLCELL_X8 FILLER_41_491 ();
 FILLCELL_X1 FILLER_41_499 ();
 FILLCELL_X8 FILLER_41_516 ();
 FILLCELL_X1 FILLER_41_542 ();
 FILLCELL_X32 FILLER_41_553 ();
 FILLCELL_X16 FILLER_41_585 ();
 FILLCELL_X8 FILLER_41_601 ();
 FILLCELL_X2 FILLER_41_609 ();
 FILLCELL_X1 FILLER_41_611 ();
 FILLCELL_X1 FILLER_41_615 ();
 FILLCELL_X1 FILLER_41_620 ();
 FILLCELL_X2 FILLER_41_624 ();
 FILLCELL_X4 FILLER_41_640 ();
 FILLCELL_X2 FILLER_41_644 ();
 FILLCELL_X1 FILLER_41_662 ();
 FILLCELL_X2 FILLER_41_674 ();
 FILLCELL_X1 FILLER_41_686 ();
 FILLCELL_X1 FILLER_41_700 ();
 FILLCELL_X1 FILLER_41_705 ();
 FILLCELL_X16 FILLER_41_710 ();
 FILLCELL_X4 FILLER_41_726 ();
 FILLCELL_X2 FILLER_41_730 ();
 FILLCELL_X1 FILLER_41_732 ();
 FILLCELL_X1 FILLER_41_740 ();
 FILLCELL_X1 FILLER_41_748 ();
 FILLCELL_X1 FILLER_41_753 ();
 FILLCELL_X2 FILLER_41_758 ();
 FILLCELL_X1 FILLER_41_760 ();
 FILLCELL_X1 FILLER_41_790 ();
 FILLCELL_X8 FILLER_41_803 ();
 FILLCELL_X4 FILLER_41_811 ();
 FILLCELL_X1 FILLER_41_815 ();
 FILLCELL_X32 FILLER_41_826 ();
 FILLCELL_X32 FILLER_41_858 ();
 FILLCELL_X32 FILLER_41_890 ();
 FILLCELL_X32 FILLER_41_922 ();
 FILLCELL_X16 FILLER_41_954 ();
 FILLCELL_X8 FILLER_41_970 ();
 FILLCELL_X4 FILLER_41_978 ();
 FILLCELL_X8 FILLER_42_1 ();
 FILLCELL_X1 FILLER_42_9 ();
 FILLCELL_X4 FILLER_42_25 ();
 FILLCELL_X8 FILLER_42_58 ();
 FILLCELL_X4 FILLER_42_66 ();
 FILLCELL_X4 FILLER_42_75 ();
 FILLCELL_X2 FILLER_42_79 ();
 FILLCELL_X8 FILLER_42_101 ();
 FILLCELL_X2 FILLER_42_109 ();
 FILLCELL_X1 FILLER_42_111 ();
 FILLCELL_X4 FILLER_42_115 ();
 FILLCELL_X2 FILLER_42_119 ();
 FILLCELL_X16 FILLER_42_123 ();
 FILLCELL_X4 FILLER_42_139 ();
 FILLCELL_X2 FILLER_42_143 ();
 FILLCELL_X1 FILLER_42_145 ();
 FILLCELL_X8 FILLER_42_153 ();
 FILLCELL_X4 FILLER_42_161 ();
 FILLCELL_X2 FILLER_42_165 ();
 FILLCELL_X1 FILLER_42_167 ();
 FILLCELL_X4 FILLER_42_181 ();
 FILLCELL_X2 FILLER_42_208 ();
 FILLCELL_X16 FILLER_42_218 ();
 FILLCELL_X2 FILLER_42_234 ();
 FILLCELL_X1 FILLER_42_236 ();
 FILLCELL_X2 FILLER_42_242 ();
 FILLCELL_X4 FILLER_42_247 ();
 FILLCELL_X32 FILLER_42_263 ();
 FILLCELL_X8 FILLER_42_295 ();
 FILLCELL_X4 FILLER_42_303 ();
 FILLCELL_X1 FILLER_42_307 ();
 FILLCELL_X1 FILLER_42_317 ();
 FILLCELL_X16 FILLER_42_323 ();
 FILLCELL_X4 FILLER_42_339 ();
 FILLCELL_X2 FILLER_42_343 ();
 FILLCELL_X1 FILLER_42_345 ();
 FILLCELL_X8 FILLER_42_369 ();
 FILLCELL_X4 FILLER_42_377 ();
 FILLCELL_X2 FILLER_42_381 ();
 FILLCELL_X1 FILLER_42_383 ();
 FILLCELL_X1 FILLER_42_393 ();
 FILLCELL_X1 FILLER_42_402 ();
 FILLCELL_X4 FILLER_42_436 ();
 FILLCELL_X2 FILLER_42_440 ();
 FILLCELL_X1 FILLER_42_446 ();
 FILLCELL_X8 FILLER_42_458 ();
 FILLCELL_X4 FILLER_42_466 ();
 FILLCELL_X2 FILLER_42_470 ();
 FILLCELL_X1 FILLER_42_472 ();
 FILLCELL_X2 FILLER_42_488 ();
 FILLCELL_X1 FILLER_42_490 ();
 FILLCELL_X16 FILLER_42_493 ();
 FILLCELL_X1 FILLER_42_509 ();
 FILLCELL_X2 FILLER_42_516 ();
 FILLCELL_X1 FILLER_42_518 ();
 FILLCELL_X2 FILLER_42_533 ();
 FILLCELL_X16 FILLER_42_538 ();
 FILLCELL_X8 FILLER_42_554 ();
 FILLCELL_X2 FILLER_42_562 ();
 FILLCELL_X1 FILLER_42_564 ();
 FILLCELL_X8 FILLER_42_593 ();
 FILLCELL_X4 FILLER_42_601 ();
 FILLCELL_X2 FILLER_42_643 ();
 FILLCELL_X1 FILLER_42_648 ();
 FILLCELL_X1 FILLER_42_651 ();
 FILLCELL_X2 FILLER_42_661 ();
 FILLCELL_X2 FILLER_42_666 ();
 FILLCELL_X2 FILLER_42_675 ();
 FILLCELL_X8 FILLER_42_690 ();
 FILLCELL_X2 FILLER_42_698 ();
 FILLCELL_X1 FILLER_42_700 ();
 FILLCELL_X2 FILLER_42_705 ();
 FILLCELL_X1 FILLER_42_707 ();
 FILLCELL_X2 FILLER_42_719 ();
 FILLCELL_X1 FILLER_42_731 ();
 FILLCELL_X1 FILLER_42_741 ();
 FILLCELL_X2 FILLER_42_774 ();
 FILLCELL_X32 FILLER_42_806 ();
 FILLCELL_X32 FILLER_42_838 ();
 FILLCELL_X32 FILLER_42_870 ();
 FILLCELL_X32 FILLER_42_902 ();
 FILLCELL_X32 FILLER_42_934 ();
 FILLCELL_X16 FILLER_42_966 ();
 FILLCELL_X8 FILLER_43_1 ();
 FILLCELL_X2 FILLER_43_9 ();
 FILLCELL_X2 FILLER_43_30 ();
 FILLCELL_X4 FILLER_43_38 ();
 FILLCELL_X1 FILLER_43_42 ();
 FILLCELL_X2 FILLER_43_52 ();
 FILLCELL_X1 FILLER_43_54 ();
 FILLCELL_X16 FILLER_43_74 ();
 FILLCELL_X4 FILLER_43_90 ();
 FILLCELL_X2 FILLER_43_94 ();
 FILLCELL_X1 FILLER_43_96 ();
 FILLCELL_X8 FILLER_43_100 ();
 FILLCELL_X4 FILLER_43_122 ();
 FILLCELL_X2 FILLER_43_126 ();
 FILLCELL_X1 FILLER_43_128 ();
 FILLCELL_X8 FILLER_43_138 ();
 FILLCELL_X1 FILLER_43_146 ();
 FILLCELL_X4 FILLER_43_162 ();
 FILLCELL_X1 FILLER_43_166 ();
 FILLCELL_X4 FILLER_43_174 ();
 FILLCELL_X2 FILLER_43_178 ();
 FILLCELL_X4 FILLER_43_203 ();
 FILLCELL_X1 FILLER_43_207 ();
 FILLCELL_X1 FILLER_43_210 ();
 FILLCELL_X4 FILLER_43_234 ();
 FILLCELL_X2 FILLER_43_262 ();
 FILLCELL_X4 FILLER_43_268 ();
 FILLCELL_X1 FILLER_43_275 ();
 FILLCELL_X16 FILLER_43_281 ();
 FILLCELL_X4 FILLER_43_297 ();
 FILLCELL_X2 FILLER_43_320 ();
 FILLCELL_X1 FILLER_43_322 ();
 FILLCELL_X1 FILLER_43_339 ();
 FILLCELL_X2 FILLER_43_343 ();
 FILLCELL_X1 FILLER_43_345 ();
 FILLCELL_X16 FILLER_43_365 ();
 FILLCELL_X8 FILLER_43_381 ();
 FILLCELL_X4 FILLER_43_389 ();
 FILLCELL_X2 FILLER_43_393 ();
 FILLCELL_X1 FILLER_43_409 ();
 FILLCELL_X2 FILLER_43_429 ();
 FILLCELL_X1 FILLER_43_431 ();
 FILLCELL_X1 FILLER_43_449 ();
 FILLCELL_X16 FILLER_43_463 ();
 FILLCELL_X8 FILLER_43_479 ();
 FILLCELL_X4 FILLER_43_487 ();
 FILLCELL_X2 FILLER_43_491 ();
 FILLCELL_X2 FILLER_43_501 ();
 FILLCELL_X2 FILLER_43_506 ();
 FILLCELL_X1 FILLER_43_524 ();
 FILLCELL_X2 FILLER_43_547 ();
 FILLCELL_X16 FILLER_43_554 ();
 FILLCELL_X8 FILLER_43_570 ();
 FILLCELL_X1 FILLER_43_578 ();
 FILLCELL_X16 FILLER_43_591 ();
 FILLCELL_X8 FILLER_43_607 ();
 FILLCELL_X2 FILLER_43_629 ();
 FILLCELL_X1 FILLER_43_631 ();
 FILLCELL_X4 FILLER_43_643 ();
 FILLCELL_X1 FILLER_43_647 ();
 FILLCELL_X2 FILLER_43_651 ();
 FILLCELL_X4 FILLER_43_659 ();
 FILLCELL_X16 FILLER_43_667 ();
 FILLCELL_X2 FILLER_43_683 ();
 FILLCELL_X1 FILLER_43_685 ();
 FILLCELL_X2 FILLER_43_702 ();
 FILLCELL_X8 FILLER_43_713 ();
 FILLCELL_X1 FILLER_43_732 ();
 FILLCELL_X4 FILLER_43_745 ();
 FILLCELL_X2 FILLER_43_749 ();
 FILLCELL_X1 FILLER_43_751 ();
 FILLCELL_X32 FILLER_43_798 ();
 FILLCELL_X32 FILLER_43_830 ();
 FILLCELL_X32 FILLER_43_862 ();
 FILLCELL_X32 FILLER_43_894 ();
 FILLCELL_X32 FILLER_43_926 ();
 FILLCELL_X16 FILLER_43_958 ();
 FILLCELL_X8 FILLER_43_974 ();
 FILLCELL_X1 FILLER_44_43 ();
 FILLCELL_X1 FILLER_44_53 ();
 FILLCELL_X1 FILLER_44_59 ();
 FILLCELL_X1 FILLER_44_63 ();
 FILLCELL_X1 FILLER_44_75 ();
 FILLCELL_X1 FILLER_44_79 ();
 FILLCELL_X1 FILLER_44_107 ();
 FILLCELL_X8 FILLER_44_134 ();
 FILLCELL_X4 FILLER_44_142 ();
 FILLCELL_X1 FILLER_44_146 ();
 FILLCELL_X32 FILLER_44_177 ();
 FILLCELL_X16 FILLER_44_209 ();
 FILLCELL_X16 FILLER_44_238 ();
 FILLCELL_X8 FILLER_44_254 ();
 FILLCELL_X8 FILLER_44_283 ();
 FILLCELL_X2 FILLER_44_291 ();
 FILLCELL_X1 FILLER_44_293 ();
 FILLCELL_X8 FILLER_44_312 ();
 FILLCELL_X2 FILLER_44_320 ();
 FILLCELL_X2 FILLER_44_335 ();
 FILLCELL_X1 FILLER_44_341 ();
 FILLCELL_X2 FILLER_44_349 ();
 FILLCELL_X1 FILLER_44_351 ();
 FILLCELL_X8 FILLER_44_362 ();
 FILLCELL_X1 FILLER_44_370 ();
 FILLCELL_X16 FILLER_44_395 ();
 FILLCELL_X8 FILLER_44_411 ();
 FILLCELL_X4 FILLER_44_419 ();
 FILLCELL_X8 FILLER_44_436 ();
 FILLCELL_X8 FILLER_44_462 ();
 FILLCELL_X4 FILLER_44_470 ();
 FILLCELL_X2 FILLER_44_474 ();
 FILLCELL_X2 FILLER_44_482 ();
 FILLCELL_X4 FILLER_44_495 ();
 FILLCELL_X1 FILLER_44_509 ();
 FILLCELL_X2 FILLER_44_521 ();
 FILLCELL_X2 FILLER_44_532 ();
 FILLCELL_X1 FILLER_44_534 ();
 FILLCELL_X1 FILLER_44_543 ();
 FILLCELL_X32 FILLER_44_563 ();
 FILLCELL_X8 FILLER_44_595 ();
 FILLCELL_X4 FILLER_44_603 ();
 FILLCELL_X4 FILLER_44_614 ();
 FILLCELL_X8 FILLER_44_622 ();
 FILLCELL_X1 FILLER_44_630 ();
 FILLCELL_X4 FILLER_44_632 ();
 FILLCELL_X2 FILLER_44_636 ();
 FILLCELL_X2 FILLER_44_644 ();
 FILLCELL_X1 FILLER_44_653 ();
 FILLCELL_X16 FILLER_44_665 ();
 FILLCELL_X2 FILLER_44_681 ();
 FILLCELL_X1 FILLER_44_683 ();
 FILLCELL_X2 FILLER_44_687 ();
 FILLCELL_X1 FILLER_44_689 ();
 FILLCELL_X1 FILLER_44_703 ();
 FILLCELL_X16 FILLER_44_709 ();
 FILLCELL_X8 FILLER_44_742 ();
 FILLCELL_X1 FILLER_44_750 ();
 FILLCELL_X1 FILLER_44_780 ();
 FILLCELL_X32 FILLER_44_806 ();
 FILLCELL_X32 FILLER_44_838 ();
 FILLCELL_X32 FILLER_44_870 ();
 FILLCELL_X32 FILLER_44_902 ();
 FILLCELL_X32 FILLER_44_934 ();
 FILLCELL_X16 FILLER_44_966 ();
 FILLCELL_X4 FILLER_45_1 ();
 FILLCELL_X2 FILLER_45_5 ();
 FILLCELL_X8 FILLER_45_43 ();
 FILLCELL_X4 FILLER_45_93 ();
 FILLCELL_X16 FILLER_45_111 ();
 FILLCELL_X8 FILLER_45_127 ();
 FILLCELL_X1 FILLER_45_135 ();
 FILLCELL_X4 FILLER_45_146 ();
 FILLCELL_X1 FILLER_45_150 ();
 FILLCELL_X4 FILLER_45_160 ();
 FILLCELL_X2 FILLER_45_164 ();
 FILLCELL_X1 FILLER_45_166 ();
 FILLCELL_X8 FILLER_45_172 ();
 FILLCELL_X1 FILLER_45_180 ();
 FILLCELL_X8 FILLER_45_200 ();
 FILLCELL_X4 FILLER_45_208 ();
 FILLCELL_X2 FILLER_45_221 ();
 FILLCELL_X1 FILLER_45_223 ();
 FILLCELL_X8 FILLER_45_246 ();
 FILLCELL_X2 FILLER_45_254 ();
 FILLCELL_X8 FILLER_45_263 ();
 FILLCELL_X2 FILLER_45_279 ();
 FILLCELL_X8 FILLER_45_290 ();
 FILLCELL_X4 FILLER_45_298 ();
 FILLCELL_X2 FILLER_45_302 ();
 FILLCELL_X1 FILLER_45_304 ();
 FILLCELL_X1 FILLER_45_312 ();
 FILLCELL_X1 FILLER_45_330 ();
 FILLCELL_X4 FILLER_45_353 ();
 FILLCELL_X2 FILLER_45_357 ();
 FILLCELL_X8 FILLER_45_362 ();
 FILLCELL_X4 FILLER_45_370 ();
 FILLCELL_X1 FILLER_45_401 ();
 FILLCELL_X1 FILLER_45_409 ();
 FILLCELL_X1 FILLER_45_424 ();
 FILLCELL_X8 FILLER_45_431 ();
 FILLCELL_X4 FILLER_45_439 ();
 FILLCELL_X2 FILLER_45_443 ();
 FILLCELL_X8 FILLER_45_467 ();
 FILLCELL_X1 FILLER_45_475 ();
 FILLCELL_X1 FILLER_45_499 ();
 FILLCELL_X1 FILLER_45_545 ();
 FILLCELL_X4 FILLER_45_554 ();
 FILLCELL_X2 FILLER_45_558 ();
 FILLCELL_X1 FILLER_45_560 ();
 FILLCELL_X1 FILLER_45_579 ();
 FILLCELL_X8 FILLER_45_583 ();
 FILLCELL_X1 FILLER_45_598 ();
 FILLCELL_X16 FILLER_45_605 ();
 FILLCELL_X8 FILLER_45_621 ();
 FILLCELL_X2 FILLER_45_629 ();
 FILLCELL_X1 FILLER_45_651 ();
 FILLCELL_X2 FILLER_45_668 ();
 FILLCELL_X1 FILLER_45_674 ();
 FILLCELL_X1 FILLER_45_678 ();
 FILLCELL_X4 FILLER_45_695 ();
 FILLCELL_X1 FILLER_45_699 ();
 FILLCELL_X1 FILLER_45_707 ();
 FILLCELL_X1 FILLER_45_717 ();
 FILLCELL_X4 FILLER_45_733 ();
 FILLCELL_X2 FILLER_45_737 ();
 FILLCELL_X1 FILLER_45_739 ();
 FILLCELL_X1 FILLER_45_760 ();
 FILLCELL_X1 FILLER_45_779 ();
 FILLCELL_X1 FILLER_45_794 ();
 FILLCELL_X1 FILLER_45_798 ();
 FILLCELL_X32 FILLER_45_808 ();
 FILLCELL_X32 FILLER_45_840 ();
 FILLCELL_X32 FILLER_45_872 ();
 FILLCELL_X32 FILLER_45_904 ();
 FILLCELL_X32 FILLER_45_936 ();
 FILLCELL_X8 FILLER_45_968 ();
 FILLCELL_X4 FILLER_45_976 ();
 FILLCELL_X2 FILLER_45_980 ();
 FILLCELL_X16 FILLER_46_1 ();
 FILLCELL_X2 FILLER_46_31 ();
 FILLCELL_X1 FILLER_46_33 ();
 FILLCELL_X2 FILLER_46_36 ();
 FILLCELL_X1 FILLER_46_38 ();
 FILLCELL_X1 FILLER_46_56 ();
 FILLCELL_X1 FILLER_46_60 ();
 FILLCELL_X16 FILLER_46_73 ();
 FILLCELL_X8 FILLER_46_89 ();
 FILLCELL_X1 FILLER_46_97 ();
 FILLCELL_X8 FILLER_46_123 ();
 FILLCELL_X4 FILLER_46_131 ();
 FILLCELL_X4 FILLER_46_146 ();
 FILLCELL_X2 FILLER_46_150 ();
 FILLCELL_X8 FILLER_46_159 ();
 FILLCELL_X4 FILLER_46_167 ();
 FILLCELL_X2 FILLER_46_171 ();
 FILLCELL_X4 FILLER_46_202 ();
 FILLCELL_X1 FILLER_46_206 ();
 FILLCELL_X1 FILLER_46_231 ();
 FILLCELL_X4 FILLER_46_249 ();
 FILLCELL_X1 FILLER_46_253 ();
 FILLCELL_X8 FILLER_46_256 ();
 FILLCELL_X2 FILLER_46_264 ();
 FILLCELL_X1 FILLER_46_266 ();
 FILLCELL_X2 FILLER_46_279 ();
 FILLCELL_X1 FILLER_46_281 ();
 FILLCELL_X2 FILLER_46_286 ();
 FILLCELL_X8 FILLER_46_291 ();
 FILLCELL_X4 FILLER_46_299 ();
 FILLCELL_X1 FILLER_46_303 ();
 FILLCELL_X4 FILLER_46_310 ();
 FILLCELL_X2 FILLER_46_314 ();
 FILLCELL_X1 FILLER_46_316 ();
 FILLCELL_X2 FILLER_46_326 ();
 FILLCELL_X2 FILLER_46_335 ();
 FILLCELL_X8 FILLER_46_346 ();
 FILLCELL_X2 FILLER_46_354 ();
 FILLCELL_X1 FILLER_46_356 ();
 FILLCELL_X1 FILLER_46_364 ();
 FILLCELL_X4 FILLER_46_369 ();
 FILLCELL_X2 FILLER_46_384 ();
 FILLCELL_X32 FILLER_46_395 ();
 FILLCELL_X8 FILLER_46_427 ();
 FILLCELL_X4 FILLER_46_435 ();
 FILLCELL_X1 FILLER_46_439 ();
 FILLCELL_X1 FILLER_46_449 ();
 FILLCELL_X4 FILLER_46_469 ();
 FILLCELL_X1 FILLER_46_473 ();
 FILLCELL_X2 FILLER_46_483 ();
 FILLCELL_X2 FILLER_46_492 ();
 FILLCELL_X8 FILLER_46_505 ();
 FILLCELL_X4 FILLER_46_513 ();
 FILLCELL_X2 FILLER_46_517 ();
 FILLCELL_X1 FILLER_46_519 ();
 FILLCELL_X16 FILLER_46_536 ();
 FILLCELL_X8 FILLER_46_552 ();
 FILLCELL_X4 FILLER_46_560 ();
 FILLCELL_X2 FILLER_46_564 ();
 FILLCELL_X1 FILLER_46_566 ();
 FILLCELL_X2 FILLER_46_577 ();
 FILLCELL_X4 FILLER_46_596 ();
 FILLCELL_X2 FILLER_46_610 ();
 FILLCELL_X1 FILLER_46_612 ();
 FILLCELL_X1 FILLER_46_630 ();
 FILLCELL_X8 FILLER_46_654 ();
 FILLCELL_X2 FILLER_46_662 ();
 FILLCELL_X2 FILLER_46_670 ();
 FILLCELL_X4 FILLER_46_694 ();
 FILLCELL_X2 FILLER_46_698 ();
 FILLCELL_X1 FILLER_46_700 ();
 FILLCELL_X4 FILLER_46_710 ();
 FILLCELL_X2 FILLER_46_714 ();
 FILLCELL_X1 FILLER_46_716 ();
 FILLCELL_X8 FILLER_46_736 ();
 FILLCELL_X1 FILLER_46_744 ();
 FILLCELL_X4 FILLER_46_750 ();
 FILLCELL_X1 FILLER_46_754 ();
 FILLCELL_X1 FILLER_46_759 ();
 FILLCELL_X4 FILLER_46_767 ();
 FILLCELL_X2 FILLER_46_771 ();
 FILLCELL_X1 FILLER_46_773 ();
 FILLCELL_X32 FILLER_46_803 ();
 FILLCELL_X32 FILLER_46_835 ();
 FILLCELL_X32 FILLER_46_867 ();
 FILLCELL_X32 FILLER_46_899 ();
 FILLCELL_X32 FILLER_46_931 ();
 FILLCELL_X16 FILLER_46_963 ();
 FILLCELL_X2 FILLER_46_979 ();
 FILLCELL_X1 FILLER_46_981 ();
 FILLCELL_X16 FILLER_47_1 ();
 FILLCELL_X4 FILLER_47_17 ();
 FILLCELL_X4 FILLER_47_23 ();
 FILLCELL_X16 FILLER_47_31 ();
 FILLCELL_X2 FILLER_47_47 ();
 FILLCELL_X1 FILLER_47_49 ();
 FILLCELL_X4 FILLER_47_81 ();
 FILLCELL_X1 FILLER_47_96 ();
 FILLCELL_X8 FILLER_47_101 ();
 FILLCELL_X4 FILLER_47_109 ();
 FILLCELL_X2 FILLER_47_113 ();
 FILLCELL_X1 FILLER_47_115 ();
 FILLCELL_X32 FILLER_47_131 ();
 FILLCELL_X16 FILLER_47_163 ();
 FILLCELL_X4 FILLER_47_179 ();
 FILLCELL_X2 FILLER_47_183 ();
 FILLCELL_X1 FILLER_47_185 ();
 FILLCELL_X1 FILLER_47_201 ();
 FILLCELL_X16 FILLER_47_225 ();
 FILLCELL_X1 FILLER_47_241 ();
 FILLCELL_X16 FILLER_47_246 ();
 FILLCELL_X4 FILLER_47_262 ();
 FILLCELL_X1 FILLER_47_278 ();
 FILLCELL_X2 FILLER_47_296 ();
 FILLCELL_X2 FILLER_47_302 ();
 FILLCELL_X2 FILLER_47_314 ();
 FILLCELL_X1 FILLER_47_316 ();
 FILLCELL_X2 FILLER_47_324 ();
 FILLCELL_X1 FILLER_47_326 ();
 FILLCELL_X8 FILLER_47_358 ();
 FILLCELL_X1 FILLER_47_366 ();
 FILLCELL_X2 FILLER_47_374 ();
 FILLCELL_X16 FILLER_47_389 ();
 FILLCELL_X1 FILLER_47_405 ();
 FILLCELL_X8 FILLER_47_412 ();
 FILLCELL_X4 FILLER_47_420 ();
 FILLCELL_X1 FILLER_47_424 ();
 FILLCELL_X4 FILLER_47_434 ();
 FILLCELL_X2 FILLER_47_485 ();
 FILLCELL_X8 FILLER_47_497 ();
 FILLCELL_X4 FILLER_47_505 ();
 FILLCELL_X2 FILLER_47_509 ();
 FILLCELL_X2 FILLER_47_518 ();
 FILLCELL_X8 FILLER_47_529 ();
 FILLCELL_X4 FILLER_47_537 ();
 FILLCELL_X1 FILLER_47_562 ();
 FILLCELL_X2 FILLER_47_570 ();
 FILLCELL_X1 FILLER_47_572 ();
 FILLCELL_X2 FILLER_47_583 ();
 FILLCELL_X4 FILLER_47_607 ();
 FILLCELL_X1 FILLER_47_624 ();
 FILLCELL_X1 FILLER_47_629 ();
 FILLCELL_X1 FILLER_47_650 ();
 FILLCELL_X8 FILLER_47_669 ();
 FILLCELL_X4 FILLER_47_677 ();
 FILLCELL_X4 FILLER_47_690 ();
 FILLCELL_X1 FILLER_47_694 ();
 FILLCELL_X4 FILLER_47_714 ();
 FILLCELL_X1 FILLER_47_725 ();
 FILLCELL_X2 FILLER_47_737 ();
 FILLCELL_X8 FILLER_47_761 ();
 FILLCELL_X2 FILLER_47_769 ();
 FILLCELL_X2 FILLER_47_778 ();
 FILLCELL_X1 FILLER_47_780 ();
 FILLCELL_X2 FILLER_47_798 ();
 FILLCELL_X1 FILLER_47_800 ();
 FILLCELL_X32 FILLER_47_805 ();
 FILLCELL_X32 FILLER_47_837 ();
 FILLCELL_X32 FILLER_47_869 ();
 FILLCELL_X32 FILLER_47_901 ();
 FILLCELL_X32 FILLER_47_933 ();
 FILLCELL_X16 FILLER_47_965 ();
 FILLCELL_X1 FILLER_47_981 ();
 FILLCELL_X16 FILLER_48_1 ();
 FILLCELL_X1 FILLER_48_17 ();
 FILLCELL_X2 FILLER_48_26 ();
 FILLCELL_X1 FILLER_48_28 ();
 FILLCELL_X8 FILLER_48_43 ();
 FILLCELL_X4 FILLER_48_51 ();
 FILLCELL_X2 FILLER_48_55 ();
 FILLCELL_X16 FILLER_48_129 ();
 FILLCELL_X8 FILLER_48_145 ();
 FILLCELL_X2 FILLER_48_153 ();
 FILLCELL_X1 FILLER_48_155 ();
 FILLCELL_X32 FILLER_48_158 ();
 FILLCELL_X16 FILLER_48_190 ();
 FILLCELL_X2 FILLER_48_206 ();
 FILLCELL_X1 FILLER_48_208 ();
 FILLCELL_X1 FILLER_48_226 ();
 FILLCELL_X1 FILLER_48_234 ();
 FILLCELL_X8 FILLER_48_247 ();
 FILLCELL_X2 FILLER_48_255 ();
 FILLCELL_X4 FILLER_48_264 ();
 FILLCELL_X1 FILLER_48_299 ();
 FILLCELL_X1 FILLER_48_335 ();
 FILLCELL_X4 FILLER_48_355 ();
 FILLCELL_X1 FILLER_48_359 ();
 FILLCELL_X2 FILLER_48_371 ();
 FILLCELL_X1 FILLER_48_373 ();
 FILLCELL_X2 FILLER_48_386 ();
 FILLCELL_X2 FILLER_48_391 ();
 FILLCELL_X1 FILLER_48_414 ();
 FILLCELL_X1 FILLER_48_419 ();
 FILLCELL_X16 FILLER_48_427 ();
 FILLCELL_X8 FILLER_48_443 ();
 FILLCELL_X4 FILLER_48_451 ();
 FILLCELL_X2 FILLER_48_455 ();
 FILLCELL_X16 FILLER_48_464 ();
 FILLCELL_X1 FILLER_48_480 ();
 FILLCELL_X4 FILLER_48_484 ();
 FILLCELL_X16 FILLER_48_493 ();
 FILLCELL_X2 FILLER_48_509 ();
 FILLCELL_X16 FILLER_48_530 ();
 FILLCELL_X4 FILLER_48_546 ();
 FILLCELL_X2 FILLER_48_550 ();
 FILLCELL_X1 FILLER_48_552 ();
 FILLCELL_X2 FILLER_48_582 ();
 FILLCELL_X1 FILLER_48_584 ();
 FILLCELL_X1 FILLER_48_599 ();
 FILLCELL_X4 FILLER_48_607 ();
 FILLCELL_X2 FILLER_48_628 ();
 FILLCELL_X1 FILLER_48_630 ();
 FILLCELL_X16 FILLER_48_632 ();
 FILLCELL_X1 FILLER_48_648 ();
 FILLCELL_X2 FILLER_48_675 ();
 FILLCELL_X1 FILLER_48_677 ();
 FILLCELL_X2 FILLER_48_683 ();
 FILLCELL_X16 FILLER_48_695 ();
 FILLCELL_X8 FILLER_48_711 ();
 FILLCELL_X2 FILLER_48_719 ();
 FILLCELL_X8 FILLER_48_725 ();
 FILLCELL_X2 FILLER_48_733 ();
 FILLCELL_X1 FILLER_48_760 ();
 FILLCELL_X4 FILLER_48_774 ();
 FILLCELL_X32 FILLER_48_796 ();
 FILLCELL_X32 FILLER_48_828 ();
 FILLCELL_X32 FILLER_48_860 ();
 FILLCELL_X32 FILLER_48_892 ();
 FILLCELL_X32 FILLER_48_924 ();
 FILLCELL_X16 FILLER_48_956 ();
 FILLCELL_X8 FILLER_48_972 ();
 FILLCELL_X2 FILLER_48_980 ();
 FILLCELL_X16 FILLER_49_1 ();
 FILLCELL_X1 FILLER_49_17 ();
 FILLCELL_X8 FILLER_49_39 ();
 FILLCELL_X1 FILLER_49_47 ();
 FILLCELL_X2 FILLER_49_61 ();
 FILLCELL_X1 FILLER_49_63 ();
 FILLCELL_X2 FILLER_49_84 ();
 FILLCELL_X2 FILLER_49_92 ();
 FILLCELL_X1 FILLER_49_94 ();
 FILLCELL_X1 FILLER_49_108 ();
 FILLCELL_X1 FILLER_49_116 ();
 FILLCELL_X1 FILLER_49_121 ();
 FILLCELL_X4 FILLER_49_129 ();
 FILLCELL_X1 FILLER_49_136 ();
 FILLCELL_X2 FILLER_49_179 ();
 FILLCELL_X1 FILLER_49_181 ();
 FILLCELL_X8 FILLER_49_185 ();
 FILLCELL_X2 FILLER_49_199 ();
 FILLCELL_X1 FILLER_49_201 ();
 FILLCELL_X4 FILLER_49_208 ();
 FILLCELL_X8 FILLER_49_224 ();
 FILLCELL_X4 FILLER_49_232 ();
 FILLCELL_X2 FILLER_49_236 ();
 FILLCELL_X1 FILLER_49_238 ();
 FILLCELL_X8 FILLER_49_242 ();
 FILLCELL_X4 FILLER_49_303 ();
 FILLCELL_X2 FILLER_49_307 ();
 FILLCELL_X2 FILLER_49_319 ();
 FILLCELL_X8 FILLER_49_353 ();
 FILLCELL_X2 FILLER_49_361 ();
 FILLCELL_X1 FILLER_49_363 ();
 FILLCELL_X1 FILLER_49_387 ();
 FILLCELL_X8 FILLER_49_397 ();
 FILLCELL_X1 FILLER_49_415 ();
 FILLCELL_X1 FILLER_49_433 ();
 FILLCELL_X8 FILLER_49_465 ();
 FILLCELL_X4 FILLER_49_473 ();
 FILLCELL_X4 FILLER_49_486 ();
 FILLCELL_X1 FILLER_49_490 ();
 FILLCELL_X4 FILLER_49_504 ();
 FILLCELL_X1 FILLER_49_508 ();
 FILLCELL_X4 FILLER_49_534 ();
 FILLCELL_X2 FILLER_49_538 ();
 FILLCELL_X8 FILLER_49_546 ();
 FILLCELL_X2 FILLER_49_554 ();
 FILLCELL_X16 FILLER_49_588 ();
 FILLCELL_X8 FILLER_49_604 ();
 FILLCELL_X4 FILLER_49_612 ();
 FILLCELL_X2 FILLER_49_616 ();
 FILLCELL_X16 FILLER_49_635 ();
 FILLCELL_X8 FILLER_49_651 ();
 FILLCELL_X4 FILLER_49_659 ();
 FILLCELL_X1 FILLER_49_676 ();
 FILLCELL_X1 FILLER_49_724 ();
 FILLCELL_X8 FILLER_49_733 ();
 FILLCELL_X8 FILLER_49_746 ();
 FILLCELL_X1 FILLER_49_778 ();
 FILLCELL_X1 FILLER_49_784 ();
 FILLCELL_X2 FILLER_49_792 ();
 FILLCELL_X32 FILLER_49_799 ();
 FILLCELL_X32 FILLER_49_831 ();
 FILLCELL_X8 FILLER_49_863 ();
 FILLCELL_X1 FILLER_49_871 ();
 FILLCELL_X32 FILLER_49_886 ();
 FILLCELL_X32 FILLER_49_918 ();
 FILLCELL_X32 FILLER_49_950 ();
 FILLCELL_X16 FILLER_50_1 ();
 FILLCELL_X2 FILLER_50_17 ();
 FILLCELL_X8 FILLER_50_52 ();
 FILLCELL_X4 FILLER_50_60 ();
 FILLCELL_X2 FILLER_50_64 ();
 FILLCELL_X16 FILLER_50_77 ();
 FILLCELL_X2 FILLER_50_102 ();
 FILLCELL_X4 FILLER_50_115 ();
 FILLCELL_X2 FILLER_50_119 ();
 FILLCELL_X1 FILLER_50_121 ();
 FILLCELL_X1 FILLER_50_153 ();
 FILLCELL_X4 FILLER_50_193 ();
 FILLCELL_X1 FILLER_50_197 ();
 FILLCELL_X2 FILLER_50_207 ();
 FILLCELL_X1 FILLER_50_209 ();
 FILLCELL_X8 FILLER_50_218 ();
 FILLCELL_X4 FILLER_50_226 ();
 FILLCELL_X2 FILLER_50_230 ();
 FILLCELL_X2 FILLER_50_234 ();
 FILLCELL_X8 FILLER_50_246 ();
 FILLCELL_X8 FILLER_50_275 ();
 FILLCELL_X1 FILLER_50_283 ();
 FILLCELL_X4 FILLER_50_295 ();
 FILLCELL_X1 FILLER_50_299 ();
 FILLCELL_X4 FILLER_50_309 ();
 FILLCELL_X1 FILLER_50_313 ();
 FILLCELL_X4 FILLER_50_319 ();
 FILLCELL_X2 FILLER_50_327 ();
 FILLCELL_X1 FILLER_50_329 ();
 FILLCELL_X4 FILLER_50_347 ();
 FILLCELL_X1 FILLER_50_351 ();
 FILLCELL_X2 FILLER_50_358 ();
 FILLCELL_X1 FILLER_50_369 ();
 FILLCELL_X1 FILLER_50_383 ();
 FILLCELL_X1 FILLER_50_393 ();
 FILLCELL_X1 FILLER_50_412 ();
 FILLCELL_X1 FILLER_50_417 ();
 FILLCELL_X4 FILLER_50_425 ();
 FILLCELL_X16 FILLER_50_436 ();
 FILLCELL_X4 FILLER_50_452 ();
 FILLCELL_X2 FILLER_50_456 ();
 FILLCELL_X1 FILLER_50_467 ();
 FILLCELL_X1 FILLER_50_487 ();
 FILLCELL_X8 FILLER_50_552 ();
 FILLCELL_X2 FILLER_50_560 ();
 FILLCELL_X4 FILLER_50_566 ();
 FILLCELL_X2 FILLER_50_570 ();
 FILLCELL_X1 FILLER_50_572 ();
 FILLCELL_X1 FILLER_50_591 ();
 FILLCELL_X4 FILLER_50_604 ();
 FILLCELL_X2 FILLER_50_608 ();
 FILLCELL_X1 FILLER_50_610 ();
 FILLCELL_X8 FILLER_50_620 ();
 FILLCELL_X2 FILLER_50_628 ();
 FILLCELL_X1 FILLER_50_630 ();
 FILLCELL_X4 FILLER_50_632 ();
 FILLCELL_X2 FILLER_50_654 ();
 FILLCELL_X1 FILLER_50_656 ();
 FILLCELL_X8 FILLER_50_661 ();
 FILLCELL_X4 FILLER_50_676 ();
 FILLCELL_X1 FILLER_50_691 ();
 FILLCELL_X2 FILLER_50_712 ();
 FILLCELL_X1 FILLER_50_730 ();
 FILLCELL_X8 FILLER_50_738 ();
 FILLCELL_X1 FILLER_50_746 ();
 FILLCELL_X1 FILLER_50_754 ();
 FILLCELL_X8 FILLER_50_761 ();
 FILLCELL_X4 FILLER_50_769 ();
 FILLCELL_X32 FILLER_50_795 ();
 FILLCELL_X16 FILLER_50_827 ();
 FILLCELL_X2 FILLER_50_843 ();
 FILLCELL_X1 FILLER_50_845 ();
 FILLCELL_X8 FILLER_50_856 ();
 FILLCELL_X4 FILLER_50_866 ();
 FILLCELL_X2 FILLER_50_870 ();
 FILLCELL_X2 FILLER_50_894 ();
 FILLCELL_X32 FILLER_50_914 ();
 FILLCELL_X32 FILLER_50_946 ();
 FILLCELL_X4 FILLER_50_978 ();
 FILLCELL_X8 FILLER_51_1 ();
 FILLCELL_X1 FILLER_51_9 ();
 FILLCELL_X2 FILLER_51_16 ();
 FILLCELL_X4 FILLER_51_60 ();
 FILLCELL_X2 FILLER_51_64 ();
 FILLCELL_X8 FILLER_51_82 ();
 FILLCELL_X4 FILLER_51_90 ();
 FILLCELL_X1 FILLER_51_94 ();
 FILLCELL_X8 FILLER_51_102 ();
 FILLCELL_X16 FILLER_51_123 ();
 FILLCELL_X4 FILLER_51_139 ();
 FILLCELL_X1 FILLER_51_152 ();
 FILLCELL_X2 FILLER_51_156 ();
 FILLCELL_X2 FILLER_51_171 ();
 FILLCELL_X1 FILLER_51_173 ();
 FILLCELL_X2 FILLER_51_181 ();
 FILLCELL_X4 FILLER_51_194 ();
 FILLCELL_X2 FILLER_51_198 ();
 FILLCELL_X2 FILLER_51_210 ();
 FILLCELL_X2 FILLER_51_217 ();
 FILLCELL_X1 FILLER_51_222 ();
 FILLCELL_X8 FILLER_51_227 ();
 FILLCELL_X1 FILLER_51_235 ();
 FILLCELL_X8 FILLER_51_252 ();
 FILLCELL_X4 FILLER_51_264 ();
 FILLCELL_X2 FILLER_51_286 ();
 FILLCELL_X2 FILLER_51_295 ();
 FILLCELL_X2 FILLER_51_302 ();
 FILLCELL_X8 FILLER_51_307 ();
 FILLCELL_X2 FILLER_51_315 ();
 FILLCELL_X1 FILLER_51_327 ();
 FILLCELL_X4 FILLER_51_335 ();
 FILLCELL_X2 FILLER_51_343 ();
 FILLCELL_X1 FILLER_51_345 ();
 FILLCELL_X1 FILLER_51_380 ();
 FILLCELL_X2 FILLER_51_409 ();
 FILLCELL_X2 FILLER_51_418 ();
 FILLCELL_X1 FILLER_51_420 ();
 FILLCELL_X8 FILLER_51_444 ();
 FILLCELL_X1 FILLER_51_492 ();
 FILLCELL_X8 FILLER_51_503 ();
 FILLCELL_X4 FILLER_51_517 ();
 FILLCELL_X1 FILLER_51_521 ();
 FILLCELL_X32 FILLER_51_525 ();
 FILLCELL_X2 FILLER_51_564 ();
 FILLCELL_X2 FILLER_51_570 ();
 FILLCELL_X1 FILLER_51_572 ();
 FILLCELL_X2 FILLER_51_580 ();
 FILLCELL_X1 FILLER_51_582 ();
 FILLCELL_X4 FILLER_51_587 ();
 FILLCELL_X8 FILLER_51_598 ();
 FILLCELL_X2 FILLER_51_611 ();
 FILLCELL_X8 FILLER_51_624 ();
 FILLCELL_X4 FILLER_51_632 ();
 FILLCELL_X2 FILLER_51_636 ();
 FILLCELL_X4 FILLER_51_649 ();
 FILLCELL_X8 FILLER_51_670 ();
 FILLCELL_X2 FILLER_51_678 ();
 FILLCELL_X4 FILLER_51_698 ();
 FILLCELL_X1 FILLER_51_718 ();
 FILLCELL_X8 FILLER_51_732 ();
 FILLCELL_X4 FILLER_51_740 ();
 FILLCELL_X1 FILLER_51_744 ();
 FILLCELL_X1 FILLER_51_775 ();
 FILLCELL_X4 FILLER_51_781 ();
 FILLCELL_X1 FILLER_51_785 ();
 FILLCELL_X8 FILLER_51_796 ();
 FILLCELL_X1 FILLER_51_804 ();
 FILLCELL_X8 FILLER_51_831 ();
 FILLCELL_X2 FILLER_51_839 ();
 FILLCELL_X1 FILLER_51_841 ();
 FILLCELL_X2 FILLER_51_879 ();
 FILLCELL_X1 FILLER_51_881 ();
 FILLCELL_X4 FILLER_51_890 ();
 FILLCELL_X2 FILLER_51_894 ();
 FILLCELL_X1 FILLER_51_896 ();
 FILLCELL_X16 FILLER_51_902 ();
 FILLCELL_X8 FILLER_51_918 ();
 FILLCELL_X8 FILLER_51_942 ();
 FILLCELL_X2 FILLER_51_956 ();
 FILLCELL_X1 FILLER_51_958 ();
 FILLCELL_X16 FILLER_51_961 ();
 FILLCELL_X4 FILLER_51_977 ();
 FILLCELL_X1 FILLER_51_981 ();
 FILLCELL_X8 FILLER_52_4 ();
 FILLCELL_X4 FILLER_52_12 ();
 FILLCELL_X1 FILLER_52_16 ();
 FILLCELL_X1 FILLER_52_20 ();
 FILLCELL_X1 FILLER_52_41 ();
 FILLCELL_X4 FILLER_52_47 ();
 FILLCELL_X1 FILLER_52_51 ();
 FILLCELL_X8 FILLER_52_63 ();
 FILLCELL_X2 FILLER_52_71 ();
 FILLCELL_X4 FILLER_52_102 ();
 FILLCELL_X1 FILLER_52_106 ();
 FILLCELL_X4 FILLER_52_145 ();
 FILLCELL_X1 FILLER_52_149 ();
 FILLCELL_X4 FILLER_52_153 ();
 FILLCELL_X2 FILLER_52_157 ();
 FILLCELL_X1 FILLER_52_159 ();
 FILLCELL_X2 FILLER_52_169 ();
 FILLCELL_X16 FILLER_52_185 ();
 FILLCELL_X1 FILLER_52_245 ();
 FILLCELL_X4 FILLER_52_253 ();
 FILLCELL_X1 FILLER_52_257 ();
 FILLCELL_X1 FILLER_52_267 ();
 FILLCELL_X16 FILLER_52_277 ();
 FILLCELL_X2 FILLER_52_293 ();
 FILLCELL_X2 FILLER_52_304 ();
 FILLCELL_X4 FILLER_52_315 ();
 FILLCELL_X1 FILLER_52_319 ();
 FILLCELL_X2 FILLER_52_356 ();
 FILLCELL_X1 FILLER_52_358 ();
 FILLCELL_X2 FILLER_52_381 ();
 FILLCELL_X1 FILLER_52_400 ();
 FILLCELL_X4 FILLER_52_443 ();
 FILLCELL_X2 FILLER_52_447 ();
 FILLCELL_X2 FILLER_52_460 ();
 FILLCELL_X2 FILLER_52_491 ();
 FILLCELL_X4 FILLER_52_506 ();
 FILLCELL_X8 FILLER_52_515 ();
 FILLCELL_X4 FILLER_52_523 ();
 FILLCELL_X1 FILLER_52_527 ();
 FILLCELL_X16 FILLER_52_532 ();
 FILLCELL_X2 FILLER_52_548 ();
 FILLCELL_X1 FILLER_52_550 ();
 FILLCELL_X16 FILLER_52_562 ();
 FILLCELL_X4 FILLER_52_578 ();
 FILLCELL_X2 FILLER_52_582 ();
 FILLCELL_X16 FILLER_52_591 ();
 FILLCELL_X2 FILLER_52_607 ();
 FILLCELL_X1 FILLER_52_609 ();
 FILLCELL_X4 FILLER_52_626 ();
 FILLCELL_X1 FILLER_52_630 ();
 FILLCELL_X1 FILLER_52_663 ();
 FILLCELL_X4 FILLER_52_687 ();
 FILLCELL_X2 FILLER_52_691 ();
 FILLCELL_X4 FILLER_52_698 ();
 FILLCELL_X1 FILLER_52_722 ();
 FILLCELL_X2 FILLER_52_734 ();
 FILLCELL_X4 FILLER_52_750 ();
 FILLCELL_X1 FILLER_52_754 ();
 FILLCELL_X4 FILLER_52_770 ();
 FILLCELL_X16 FILLER_52_781 ();
 FILLCELL_X2 FILLER_52_797 ();
 FILLCELL_X1 FILLER_52_799 ();
 FILLCELL_X4 FILLER_52_810 ();
 FILLCELL_X2 FILLER_52_814 ();
 FILLCELL_X2 FILLER_52_832 ();
 FILLCELL_X8 FILLER_52_836 ();
 FILLCELL_X4 FILLER_52_844 ();
 FILLCELL_X1 FILLER_52_848 ();
 FILLCELL_X2 FILLER_52_865 ();
 FILLCELL_X16 FILLER_52_869 ();
 FILLCELL_X2 FILLER_52_885 ();
 FILLCELL_X1 FILLER_52_887 ();
 FILLCELL_X16 FILLER_52_962 ();
 FILLCELL_X4 FILLER_52_978 ();
 FILLCELL_X2 FILLER_53_1 ();
 FILLCELL_X1 FILLER_53_3 ();
 FILLCELL_X1 FILLER_53_7 ();
 FILLCELL_X8 FILLER_53_11 ();
 FILLCELL_X2 FILLER_53_19 ();
 FILLCELL_X4 FILLER_53_27 ();
 FILLCELL_X2 FILLER_53_31 ();
 FILLCELL_X2 FILLER_53_63 ();
 FILLCELL_X2 FILLER_53_85 ();
 FILLCELL_X2 FILLER_53_97 ();
 FILLCELL_X2 FILLER_53_105 ();
 FILLCELL_X1 FILLER_53_107 ();
 FILLCELL_X1 FILLER_53_118 ();
 FILLCELL_X4 FILLER_53_132 ();
 FILLCELL_X1 FILLER_53_136 ();
 FILLCELL_X2 FILLER_53_150 ();
 FILLCELL_X4 FILLER_53_165 ();
 FILLCELL_X1 FILLER_53_169 ();
 FILLCELL_X4 FILLER_53_177 ();
 FILLCELL_X4 FILLER_53_217 ();
 FILLCELL_X16 FILLER_53_226 ();
 FILLCELL_X2 FILLER_53_242 ();
 FILLCELL_X8 FILLER_53_250 ();
 FILLCELL_X2 FILLER_53_258 ();
 FILLCELL_X1 FILLER_53_260 ();
 FILLCELL_X1 FILLER_53_286 ();
 FILLCELL_X4 FILLER_53_292 ();
 FILLCELL_X2 FILLER_53_296 ();
 FILLCELL_X4 FILLER_53_316 ();
 FILLCELL_X2 FILLER_53_320 ();
 FILLCELL_X1 FILLER_53_322 ();
 FILLCELL_X16 FILLER_53_349 ();
 FILLCELL_X8 FILLER_53_372 ();
 FILLCELL_X1 FILLER_53_380 ();
 FILLCELL_X4 FILLER_53_394 ();
 FILLCELL_X1 FILLER_53_398 ();
 FILLCELL_X8 FILLER_53_420 ();
 FILLCELL_X4 FILLER_53_428 ();
 FILLCELL_X2 FILLER_53_439 ();
 FILLCELL_X4 FILLER_53_464 ();
 FILLCELL_X1 FILLER_53_484 ();
 FILLCELL_X1 FILLER_53_501 ();
 FILLCELL_X2 FILLER_53_519 ();
 FILLCELL_X1 FILLER_53_532 ();
 FILLCELL_X1 FILLER_53_537 ();
 FILLCELL_X2 FILLER_53_555 ();
 FILLCELL_X8 FILLER_53_564 ();
 FILLCELL_X4 FILLER_53_572 ();
 FILLCELL_X1 FILLER_53_576 ();
 FILLCELL_X1 FILLER_53_580 ();
 FILLCELL_X8 FILLER_53_592 ();
 FILLCELL_X1 FILLER_53_600 ();
 FILLCELL_X2 FILLER_53_606 ();
 FILLCELL_X8 FILLER_53_622 ();
 FILLCELL_X4 FILLER_53_630 ();
 FILLCELL_X1 FILLER_53_634 ();
 FILLCELL_X1 FILLER_53_640 ();
 FILLCELL_X2 FILLER_53_669 ();
 FILLCELL_X8 FILLER_53_689 ();
 FILLCELL_X1 FILLER_53_697 ();
 FILLCELL_X2 FILLER_53_720 ();
 FILLCELL_X4 FILLER_53_729 ();
 FILLCELL_X32 FILLER_53_762 ();
 FILLCELL_X8 FILLER_53_794 ();
 FILLCELL_X1 FILLER_53_802 ();
 FILLCELL_X2 FILLER_53_805 ();
 FILLCELL_X8 FILLER_53_823 ();
 FILLCELL_X4 FILLER_53_831 ();
 FILLCELL_X1 FILLER_53_835 ();
 FILLCELL_X2 FILLER_53_846 ();
 FILLCELL_X8 FILLER_53_858 ();
 FILLCELL_X4 FILLER_53_866 ();
 FILLCELL_X1 FILLER_53_870 ();
 FILLCELL_X4 FILLER_53_873 ();
 FILLCELL_X1 FILLER_53_887 ();
 FILLCELL_X16 FILLER_53_890 ();
 FILLCELL_X4 FILLER_53_906 ();
 FILLCELL_X4 FILLER_53_920 ();
 FILLCELL_X1 FILLER_53_924 ();
 FILLCELL_X8 FILLER_53_927 ();
 FILLCELL_X2 FILLER_53_935 ();
 FILLCELL_X4 FILLER_53_939 ();
 FILLCELL_X1 FILLER_53_943 ();
 FILLCELL_X1 FILLER_53_960 ();
 FILLCELL_X4 FILLER_53_975 ();
 FILLCELL_X2 FILLER_53_979 ();
 FILLCELL_X1 FILLER_53_981 ();
 FILLCELL_X32 FILLER_54_1 ();
 FILLCELL_X4 FILLER_54_33 ();
 FILLCELL_X2 FILLER_54_45 ();
 FILLCELL_X2 FILLER_54_73 ();
 FILLCELL_X2 FILLER_54_85 ();
 FILLCELL_X1 FILLER_54_87 ();
 FILLCELL_X1 FILLER_54_101 ();
 FILLCELL_X8 FILLER_54_127 ();
 FILLCELL_X4 FILLER_54_135 ();
 FILLCELL_X4 FILLER_54_161 ();
 FILLCELL_X2 FILLER_54_208 ();
 FILLCELL_X2 FILLER_54_232 ();
 FILLCELL_X2 FILLER_54_238 ();
 FILLCELL_X1 FILLER_54_249 ();
 FILLCELL_X4 FILLER_54_274 ();
 FILLCELL_X1 FILLER_54_285 ();
 FILLCELL_X2 FILLER_54_295 ();
 FILLCELL_X4 FILLER_54_311 ();
 FILLCELL_X1 FILLER_54_333 ();
 FILLCELL_X1 FILLER_54_339 ();
 FILLCELL_X1 FILLER_54_351 ();
 FILLCELL_X4 FILLER_54_360 ();
 FILLCELL_X2 FILLER_54_367 ();
 FILLCELL_X1 FILLER_54_373 ();
 FILLCELL_X2 FILLER_54_383 ();
 FILLCELL_X2 FILLER_54_397 ();
 FILLCELL_X2 FILLER_54_421 ();
 FILLCELL_X1 FILLER_54_423 ();
 FILLCELL_X16 FILLER_54_436 ();
 FILLCELL_X4 FILLER_54_452 ();
 FILLCELL_X2 FILLER_54_456 ();
 FILLCELL_X8 FILLER_54_472 ();
 FILLCELL_X2 FILLER_54_480 ();
 FILLCELL_X1 FILLER_54_489 ();
 FILLCELL_X8 FILLER_54_494 ();
 FILLCELL_X1 FILLER_54_508 ();
 FILLCELL_X1 FILLER_54_514 ();
 FILLCELL_X1 FILLER_54_528 ();
 FILLCELL_X2 FILLER_54_546 ();
 FILLCELL_X1 FILLER_54_551 ();
 FILLCELL_X2 FILLER_54_595 ();
 FILLCELL_X1 FILLER_54_597 ();
 FILLCELL_X4 FILLER_54_604 ();
 FILLCELL_X2 FILLER_54_608 ();
 FILLCELL_X2 FILLER_54_614 ();
 FILLCELL_X8 FILLER_54_619 ();
 FILLCELL_X4 FILLER_54_627 ();
 FILLCELL_X2 FILLER_54_632 ();
 FILLCELL_X1 FILLER_54_643 ();
 FILLCELL_X2 FILLER_54_648 ();
 FILLCELL_X2 FILLER_54_654 ();
 FILLCELL_X4 FILLER_54_669 ();
 FILLCELL_X2 FILLER_54_673 ();
 FILLCELL_X2 FILLER_54_684 ();
 FILLCELL_X1 FILLER_54_686 ();
 FILLCELL_X1 FILLER_54_704 ();
 FILLCELL_X2 FILLER_54_723 ();
 FILLCELL_X2 FILLER_54_731 ();
 FILLCELL_X1 FILLER_54_746 ();
 FILLCELL_X32 FILLER_54_762 ();
 FILLCELL_X8 FILLER_54_794 ();
 FILLCELL_X8 FILLER_54_818 ();
 FILLCELL_X2 FILLER_54_826 ();
 FILLCELL_X2 FILLER_54_844 ();
 FILLCELL_X4 FILLER_54_862 ();
 FILLCELL_X2 FILLER_54_866 ();
 FILLCELL_X16 FILLER_54_878 ();
 FILLCELL_X8 FILLER_54_894 ();
 FILLCELL_X2 FILLER_54_920 ();
 FILLCELL_X16 FILLER_54_938 ();
 FILLCELL_X4 FILLER_54_954 ();
 FILLCELL_X1 FILLER_54_958 ();
 FILLCELL_X4 FILLER_54_975 ();
 FILLCELL_X2 FILLER_54_979 ();
 FILLCELL_X1 FILLER_54_981 ();
 FILLCELL_X32 FILLER_55_1 ();
 FILLCELL_X16 FILLER_55_33 ();
 FILLCELL_X1 FILLER_55_59 ();
 FILLCELL_X1 FILLER_55_69 ();
 FILLCELL_X1 FILLER_55_81 ();
 FILLCELL_X2 FILLER_55_121 ();
 FILLCELL_X4 FILLER_55_136 ();
 FILLCELL_X1 FILLER_55_144 ();
 FILLCELL_X1 FILLER_55_239 ();
 FILLCELL_X16 FILLER_55_262 ();
 FILLCELL_X4 FILLER_55_278 ();
 FILLCELL_X2 FILLER_55_282 ();
 FILLCELL_X1 FILLER_55_284 ();
 FILLCELL_X4 FILLER_55_295 ();
 FILLCELL_X1 FILLER_55_325 ();
 FILLCELL_X4 FILLER_55_331 ();
 FILLCELL_X2 FILLER_55_335 ();
 FILLCELL_X4 FILLER_55_342 ();
 FILLCELL_X2 FILLER_55_346 ();
 FILLCELL_X8 FILLER_55_364 ();
 FILLCELL_X1 FILLER_55_372 ();
 FILLCELL_X4 FILLER_55_383 ();
 FILLCELL_X1 FILLER_55_387 ();
 FILLCELL_X1 FILLER_55_398 ();
 FILLCELL_X1 FILLER_55_403 ();
 FILLCELL_X4 FILLER_55_408 ();
 FILLCELL_X1 FILLER_55_412 ();
 FILLCELL_X4 FILLER_55_420 ();
 FILLCELL_X1 FILLER_55_437 ();
 FILLCELL_X4 FILLER_55_448 ();
 FILLCELL_X2 FILLER_55_452 ();
 FILLCELL_X4 FILLER_55_481 ();
 FILLCELL_X16 FILLER_55_500 ();
 FILLCELL_X4 FILLER_55_516 ();
 FILLCELL_X2 FILLER_55_540 ();
 FILLCELL_X1 FILLER_55_542 ();
 FILLCELL_X4 FILLER_55_566 ();
 FILLCELL_X4 FILLER_55_575 ();
 FILLCELL_X2 FILLER_55_579 ();
 FILLCELL_X1 FILLER_55_581 ();
 FILLCELL_X1 FILLER_55_589 ();
 FILLCELL_X1 FILLER_55_595 ();
 FILLCELL_X8 FILLER_55_606 ();
 FILLCELL_X1 FILLER_55_618 ();
 FILLCELL_X4 FILLER_55_645 ();
 FILLCELL_X2 FILLER_55_649 ();
 FILLCELL_X1 FILLER_55_664 ();
 FILLCELL_X1 FILLER_55_668 ();
 FILLCELL_X2 FILLER_55_697 ();
 FILLCELL_X1 FILLER_55_699 ();
 FILLCELL_X1 FILLER_55_712 ();
 FILLCELL_X1 FILLER_55_722 ();
 FILLCELL_X4 FILLER_55_750 ();
 FILLCELL_X8 FILLER_55_772 ();
 FILLCELL_X2 FILLER_55_780 ();
 FILLCELL_X8 FILLER_55_798 ();
 FILLCELL_X4 FILLER_55_806 ();
 FILLCELL_X1 FILLER_55_810 ();
 FILLCELL_X16 FILLER_55_813 ();
 FILLCELL_X2 FILLER_55_849 ();
 FILLCELL_X8 FILLER_55_877 ();
 FILLCELL_X2 FILLER_55_885 ();
 FILLCELL_X1 FILLER_55_887 ();
 FILLCELL_X2 FILLER_55_904 ();
 FILLCELL_X16 FILLER_55_908 ();
 FILLCELL_X4 FILLER_55_924 ();
 FILLCELL_X1 FILLER_55_928 ();
 FILLCELL_X4 FILLER_55_931 ();
 FILLCELL_X2 FILLER_55_935 ();
 FILLCELL_X1 FILLER_55_937 ();
 FILLCELL_X16 FILLER_55_948 ();
 FILLCELL_X1 FILLER_55_964 ();
 FILLCELL_X4 FILLER_55_975 ();
 FILLCELL_X2 FILLER_55_979 ();
 FILLCELL_X1 FILLER_55_981 ();
 FILLCELL_X32 FILLER_56_1 ();
 FILLCELL_X32 FILLER_56_33 ();
 FILLCELL_X2 FILLER_56_65 ();
 FILLCELL_X1 FILLER_56_67 ();
 FILLCELL_X8 FILLER_56_78 ();
 FILLCELL_X1 FILLER_56_86 ();
 FILLCELL_X2 FILLER_56_94 ();
 FILLCELL_X1 FILLER_56_106 ();
 FILLCELL_X2 FILLER_56_136 ();
 FILLCELL_X1 FILLER_56_151 ();
 FILLCELL_X1 FILLER_56_181 ();
 FILLCELL_X2 FILLER_56_202 ();
 FILLCELL_X1 FILLER_56_204 ();
 FILLCELL_X4 FILLER_56_262 ();
 FILLCELL_X2 FILLER_56_266 ();
 FILLCELL_X2 FILLER_56_288 ();
 FILLCELL_X1 FILLER_56_290 ();
 FILLCELL_X16 FILLER_56_296 ();
 FILLCELL_X4 FILLER_56_312 ();
 FILLCELL_X2 FILLER_56_316 ();
 FILLCELL_X1 FILLER_56_318 ();
 FILLCELL_X4 FILLER_56_332 ();
 FILLCELL_X2 FILLER_56_353 ();
 FILLCELL_X1 FILLER_56_362 ();
 FILLCELL_X2 FILLER_56_367 ();
 FILLCELL_X2 FILLER_56_388 ();
 FILLCELL_X8 FILLER_56_404 ();
 FILLCELL_X1 FILLER_56_412 ();
 FILLCELL_X2 FILLER_56_418 ();
 FILLCELL_X4 FILLER_56_424 ();
 FILLCELL_X4 FILLER_56_435 ();
 FILLCELL_X2 FILLER_56_439 ();
 FILLCELL_X8 FILLER_56_447 ();
 FILLCELL_X4 FILLER_56_455 ();
 FILLCELL_X2 FILLER_56_459 ();
 FILLCELL_X1 FILLER_56_461 ();
 FILLCELL_X2 FILLER_56_508 ();
 FILLCELL_X1 FILLER_56_510 ();
 FILLCELL_X4 FILLER_56_524 ();
 FILLCELL_X1 FILLER_56_535 ();
 FILLCELL_X4 FILLER_56_540 ();
 FILLCELL_X2 FILLER_56_544 ();
 FILLCELL_X1 FILLER_56_559 ();
 FILLCELL_X4 FILLER_56_585 ();
 FILLCELL_X1 FILLER_56_589 ();
 FILLCELL_X1 FILLER_56_614 ();
 FILLCELL_X4 FILLER_56_620 ();
 FILLCELL_X2 FILLER_56_624 ();
 FILLCELL_X2 FILLER_56_645 ();
 FILLCELL_X2 FILLER_56_660 ();
 FILLCELL_X4 FILLER_56_667 ();
 FILLCELL_X2 FILLER_56_671 ();
 FILLCELL_X1 FILLER_56_673 ();
 FILLCELL_X2 FILLER_56_704 ();
 FILLCELL_X1 FILLER_56_706 ();
 FILLCELL_X4 FILLER_56_714 ();
 FILLCELL_X4 FILLER_56_725 ();
 FILLCELL_X1 FILLER_56_729 ();
 FILLCELL_X1 FILLER_56_734 ();
 FILLCELL_X8 FILLER_56_750 ();
 FILLCELL_X4 FILLER_56_778 ();
 FILLCELL_X1 FILLER_56_782 ();
 FILLCELL_X2 FILLER_56_785 ();
 FILLCELL_X2 FILLER_56_825 ();
 FILLCELL_X1 FILLER_56_843 ();
 FILLCELL_X2 FILLER_56_872 ();
 FILLCELL_X1 FILLER_56_874 ();
 FILLCELL_X4 FILLER_56_891 ();
 FILLCELL_X2 FILLER_56_895 ();
 FILLCELL_X2 FILLER_56_907 ();
 FILLCELL_X1 FILLER_56_909 ();
 FILLCELL_X2 FILLER_56_926 ();
 FILLCELL_X1 FILLER_56_928 ();
 FILLCELL_X2 FILLER_56_939 ();
 FILLCELL_X2 FILLER_56_943 ();
 FILLCELL_X1 FILLER_56_945 ();
 FILLCELL_X8 FILLER_56_948 ();
 FILLCELL_X4 FILLER_56_956 ();
 FILLCELL_X2 FILLER_56_960 ();
 FILLCELL_X4 FILLER_56_978 ();
 FILLCELL_X32 FILLER_57_1 ();
 FILLCELL_X32 FILLER_57_33 ();
 FILLCELL_X4 FILLER_57_65 ();
 FILLCELL_X1 FILLER_57_138 ();
 FILLCELL_X1 FILLER_57_150 ();
 FILLCELL_X1 FILLER_57_156 ();
 FILLCELL_X1 FILLER_57_170 ();
 FILLCELL_X1 FILLER_57_173 ();
 FILLCELL_X1 FILLER_57_177 ();
 FILLCELL_X1 FILLER_57_191 ();
 FILLCELL_X1 FILLER_57_197 ();
 FILLCELL_X2 FILLER_57_205 ();
 FILLCELL_X1 FILLER_57_211 ();
 FILLCELL_X1 FILLER_57_224 ();
 FILLCELL_X1 FILLER_57_231 ();
 FILLCELL_X1 FILLER_57_239 ();
 FILLCELL_X1 FILLER_57_251 ();
 FILLCELL_X1 FILLER_57_256 ();
 FILLCELL_X16 FILLER_57_264 ();
 FILLCELL_X4 FILLER_57_280 ();
 FILLCELL_X8 FILLER_57_290 ();
 FILLCELL_X4 FILLER_57_298 ();
 FILLCELL_X2 FILLER_57_302 ();
 FILLCELL_X4 FILLER_57_347 ();
 FILLCELL_X2 FILLER_57_351 ();
 FILLCELL_X2 FILLER_57_359 ();
 FILLCELL_X1 FILLER_57_361 ();
 FILLCELL_X2 FILLER_57_376 ();
 FILLCELL_X1 FILLER_57_378 ();
 FILLCELL_X4 FILLER_57_384 ();
 FILLCELL_X1 FILLER_57_394 ();
 FILLCELL_X1 FILLER_57_400 ();
 FILLCELL_X2 FILLER_57_406 ();
 FILLCELL_X1 FILLER_57_421 ();
 FILLCELL_X1 FILLER_57_431 ();
 FILLCELL_X1 FILLER_57_434 ();
 FILLCELL_X2 FILLER_57_438 ();
 FILLCELL_X16 FILLER_57_444 ();
 FILLCELL_X2 FILLER_57_460 ();
 FILLCELL_X1 FILLER_57_462 ();
 FILLCELL_X1 FILLER_57_485 ();
 FILLCELL_X2 FILLER_57_489 ();
 FILLCELL_X8 FILLER_57_494 ();
 FILLCELL_X8 FILLER_57_519 ();
 FILLCELL_X2 FILLER_57_527 ();
 FILLCELL_X1 FILLER_57_529 ();
 FILLCELL_X2 FILLER_57_534 ();
 FILLCELL_X16 FILLER_57_560 ();
 FILLCELL_X8 FILLER_57_576 ();
 FILLCELL_X2 FILLER_57_584 ();
 FILLCELL_X16 FILLER_57_606 ();
 FILLCELL_X1 FILLER_57_622 ();
 FILLCELL_X1 FILLER_57_661 ();
 FILLCELL_X2 FILLER_57_665 ();
 FILLCELL_X1 FILLER_57_686 ();
 FILLCELL_X1 FILLER_57_691 ();
 FILLCELL_X1 FILLER_57_699 ();
 FILLCELL_X1 FILLER_57_704 ();
 FILLCELL_X16 FILLER_57_717 ();
 FILLCELL_X2 FILLER_57_733 ();
 FILLCELL_X1 FILLER_57_735 ();
 FILLCELL_X16 FILLER_57_745 ();
 FILLCELL_X2 FILLER_57_761 ();
 FILLCELL_X32 FILLER_57_783 ();
 FILLCELL_X4 FILLER_57_815 ();
 FILLCELL_X2 FILLER_57_819 ();
 FILLCELL_X1 FILLER_57_821 ();
 FILLCELL_X16 FILLER_57_824 ();
 FILLCELL_X2 FILLER_57_840 ();
 FILLCELL_X16 FILLER_57_844 ();
 FILLCELL_X8 FILLER_57_860 ();
 FILLCELL_X4 FILLER_57_868 ();
 FILLCELL_X4 FILLER_57_874 ();
 FILLCELL_X2 FILLER_57_878 ();
 FILLCELL_X1 FILLER_57_880 ();
 FILLCELL_X4 FILLER_57_909 ();
 FILLCELL_X2 FILLER_57_939 ();
 FILLCELL_X1 FILLER_57_941 ();
 FILLCELL_X4 FILLER_57_962 ();
 FILLCELL_X32 FILLER_58_1 ();
 FILLCELL_X32 FILLER_58_33 ();
 FILLCELL_X16 FILLER_58_65 ();
 FILLCELL_X4 FILLER_58_81 ();
 FILLCELL_X4 FILLER_58_117 ();
 FILLCELL_X1 FILLER_58_121 ();
 FILLCELL_X4 FILLER_58_135 ();
 FILLCELL_X2 FILLER_58_148 ();
 FILLCELL_X1 FILLER_58_150 ();
 FILLCELL_X2 FILLER_58_158 ();
 FILLCELL_X1 FILLER_58_160 ();
 FILLCELL_X2 FILLER_58_209 ();
 FILLCELL_X1 FILLER_58_211 ();
 FILLCELL_X2 FILLER_58_226 ();
 FILLCELL_X1 FILLER_58_228 ();
 FILLCELL_X8 FILLER_58_243 ();
 FILLCELL_X2 FILLER_58_251 ();
 FILLCELL_X2 FILLER_58_258 ();
 FILLCELL_X1 FILLER_58_260 ();
 FILLCELL_X2 FILLER_58_270 ();
 FILLCELL_X4 FILLER_58_275 ();
 FILLCELL_X1 FILLER_58_279 ();
 FILLCELL_X2 FILLER_58_289 ();
 FILLCELL_X2 FILLER_58_301 ();
 FILLCELL_X8 FILLER_58_321 ();
 FILLCELL_X4 FILLER_58_329 ();
 FILLCELL_X2 FILLER_58_337 ();
 FILLCELL_X1 FILLER_58_339 ();
 FILLCELL_X4 FILLER_58_344 ();
 FILLCELL_X4 FILLER_58_366 ();
 FILLCELL_X1 FILLER_58_370 ();
 FILLCELL_X1 FILLER_58_380 ();
 FILLCELL_X1 FILLER_58_388 ();
 FILLCELL_X1 FILLER_58_398 ();
 FILLCELL_X1 FILLER_58_406 ();
 FILLCELL_X2 FILLER_58_435 ();
 FILLCELL_X1 FILLER_58_437 ();
 FILLCELL_X2 FILLER_58_443 ();
 FILLCELL_X1 FILLER_58_470 ();
 FILLCELL_X2 FILLER_58_475 ();
 FILLCELL_X4 FILLER_58_480 ();
 FILLCELL_X2 FILLER_58_484 ();
 FILLCELL_X8 FILLER_58_493 ();
 FILLCELL_X1 FILLER_58_501 ();
 FILLCELL_X4 FILLER_58_510 ();
 FILLCELL_X8 FILLER_58_517 ();
 FILLCELL_X4 FILLER_58_534 ();
 FILLCELL_X2 FILLER_58_538 ();
 FILLCELL_X4 FILLER_58_547 ();
 FILLCELL_X2 FILLER_58_551 ();
 FILLCELL_X8 FILLER_58_567 ();
 FILLCELL_X16 FILLER_58_589 ();
 FILLCELL_X8 FILLER_58_605 ();
 FILLCELL_X4 FILLER_58_613 ();
 FILLCELL_X4 FILLER_58_632 ();
 FILLCELL_X2 FILLER_58_659 ();
 FILLCELL_X8 FILLER_58_666 ();
 FILLCELL_X2 FILLER_58_674 ();
 FILLCELL_X2 FILLER_58_687 ();
 FILLCELL_X4 FILLER_58_702 ();
 FILLCELL_X2 FILLER_58_706 ();
 FILLCELL_X1 FILLER_58_708 ();
 FILLCELL_X4 FILLER_58_722 ();
 FILLCELL_X1 FILLER_58_726 ();
 FILLCELL_X4 FILLER_58_742 ();
 FILLCELL_X4 FILLER_58_749 ();
 FILLCELL_X1 FILLER_58_753 ();
 FILLCELL_X4 FILLER_58_764 ();
 FILLCELL_X1 FILLER_58_768 ();
 FILLCELL_X16 FILLER_58_783 ();
 FILLCELL_X2 FILLER_58_799 ();
 FILLCELL_X1 FILLER_58_801 ();
 FILLCELL_X32 FILLER_58_804 ();
 FILLCELL_X2 FILLER_58_836 ();
 FILLCELL_X8 FILLER_58_854 ();
 FILLCELL_X2 FILLER_58_862 ();
 FILLCELL_X1 FILLER_58_864 ();
 FILLCELL_X4 FILLER_58_867 ();
 FILLCELL_X32 FILLER_58_889 ();
 FILLCELL_X2 FILLER_58_921 ();
 FILLCELL_X1 FILLER_58_923 ();
 FILLCELL_X16 FILLER_58_940 ();
 FILLCELL_X8 FILLER_58_972 ();
 FILLCELL_X2 FILLER_58_980 ();
 FILLCELL_X32 FILLER_59_1 ();
 FILLCELL_X32 FILLER_59_33 ();
 FILLCELL_X16 FILLER_59_65 ();
 FILLCELL_X8 FILLER_59_81 ();
 FILLCELL_X4 FILLER_59_89 ();
 FILLCELL_X4 FILLER_59_97 ();
 FILLCELL_X2 FILLER_59_101 ();
 FILLCELL_X1 FILLER_59_103 ();
 FILLCELL_X4 FILLER_59_113 ();
 FILLCELL_X2 FILLER_59_117 ();
 FILLCELL_X1 FILLER_59_128 ();
 FILLCELL_X8 FILLER_59_140 ();
 FILLCELL_X1 FILLER_59_161 ();
 FILLCELL_X2 FILLER_59_182 ();
 FILLCELL_X2 FILLER_59_216 ();
 FILLCELL_X1 FILLER_59_218 ();
 FILLCELL_X2 FILLER_59_224 ();
 FILLCELL_X4 FILLER_59_255 ();
 FILLCELL_X1 FILLER_59_259 ();
 FILLCELL_X4 FILLER_59_276 ();
 FILLCELL_X2 FILLER_59_280 ();
 FILLCELL_X1 FILLER_59_282 ();
 FILLCELL_X2 FILLER_59_290 ();
 FILLCELL_X2 FILLER_59_301 ();
 FILLCELL_X1 FILLER_59_303 ();
 FILLCELL_X2 FILLER_59_307 ();
 FILLCELL_X2 FILLER_59_320 ();
 FILLCELL_X1 FILLER_59_322 ();
 FILLCELL_X1 FILLER_59_336 ();
 FILLCELL_X1 FILLER_59_341 ();
 FILLCELL_X4 FILLER_59_346 ();
 FILLCELL_X1 FILLER_59_350 ();
 FILLCELL_X1 FILLER_59_385 ();
 FILLCELL_X8 FILLER_59_395 ();
 FILLCELL_X2 FILLER_59_403 ();
 FILLCELL_X1 FILLER_59_405 ();
 FILLCELL_X4 FILLER_59_411 ();
 FILLCELL_X2 FILLER_59_425 ();
 FILLCELL_X1 FILLER_59_427 ();
 FILLCELL_X8 FILLER_59_441 ();
 FILLCELL_X4 FILLER_59_449 ();
 FILLCELL_X1 FILLER_59_453 ();
 FILLCELL_X1 FILLER_59_458 ();
 FILLCELL_X2 FILLER_59_466 ();
 FILLCELL_X1 FILLER_59_468 ();
 FILLCELL_X8 FILLER_59_474 ();
 FILLCELL_X2 FILLER_59_482 ();
 FILLCELL_X2 FILLER_59_496 ();
 FILLCELL_X2 FILLER_59_501 ();
 FILLCELL_X1 FILLER_59_503 ();
 FILLCELL_X2 FILLER_59_508 ();
 FILLCELL_X1 FILLER_59_510 ();
 FILLCELL_X8 FILLER_59_526 ();
 FILLCELL_X2 FILLER_59_534 ();
 FILLCELL_X1 FILLER_59_536 ();
 FILLCELL_X4 FILLER_59_550 ();
 FILLCELL_X2 FILLER_59_569 ();
 FILLCELL_X1 FILLER_59_571 ();
 FILLCELL_X8 FILLER_59_595 ();
 FILLCELL_X4 FILLER_59_603 ();
 FILLCELL_X2 FILLER_59_607 ();
 FILLCELL_X1 FILLER_59_609 ();
 FILLCELL_X4 FILLER_59_639 ();
 FILLCELL_X2 FILLER_59_643 ();
 FILLCELL_X1 FILLER_59_645 ();
 FILLCELL_X1 FILLER_59_653 ();
 FILLCELL_X4 FILLER_59_723 ();
 FILLCELL_X1 FILLER_59_738 ();
 FILLCELL_X8 FILLER_59_744 ();
 FILLCELL_X2 FILLER_59_752 ();
 FILLCELL_X2 FILLER_59_764 ();
 FILLCELL_X1 FILLER_59_766 ();
 FILLCELL_X1 FILLER_59_769 ();
 FILLCELL_X1 FILLER_59_786 ();
 FILLCELL_X1 FILLER_59_789 ();
 FILLCELL_X1 FILLER_59_822 ();
 FILLCELL_X32 FILLER_59_839 ();
 FILLCELL_X32 FILLER_59_871 ();
 FILLCELL_X16 FILLER_59_903 ();
 FILLCELL_X8 FILLER_59_919 ();
 FILLCELL_X4 FILLER_59_927 ();
 FILLCELL_X8 FILLER_59_970 ();
 FILLCELL_X4 FILLER_59_978 ();
 FILLCELL_X16 FILLER_60_1 ();
 FILLCELL_X8 FILLER_60_17 ();
 FILLCELL_X2 FILLER_60_25 ();
 FILLCELL_X1 FILLER_60_27 ();
 FILLCELL_X32 FILLER_60_34 ();
 FILLCELL_X8 FILLER_60_66 ();
 FILLCELL_X4 FILLER_60_74 ();
 FILLCELL_X8 FILLER_60_95 ();
 FILLCELL_X32 FILLER_60_120 ();
 FILLCELL_X32 FILLER_60_152 ();
 FILLCELL_X8 FILLER_60_184 ();
 FILLCELL_X4 FILLER_60_192 ();
 FILLCELL_X1 FILLER_60_196 ();
 FILLCELL_X4 FILLER_60_218 ();
 FILLCELL_X2 FILLER_60_222 ();
 FILLCELL_X1 FILLER_60_224 ();
 FILLCELL_X8 FILLER_60_232 ();
 FILLCELL_X4 FILLER_60_240 ();
 FILLCELL_X2 FILLER_60_244 ();
 FILLCELL_X2 FILLER_60_255 ();
 FILLCELL_X4 FILLER_60_275 ();
 FILLCELL_X1 FILLER_60_279 ();
 FILLCELL_X8 FILLER_60_296 ();
 FILLCELL_X1 FILLER_60_343 ();
 FILLCELL_X2 FILLER_60_347 ();
 FILLCELL_X1 FILLER_60_349 ();
 FILLCELL_X8 FILLER_60_368 ();
 FILLCELL_X2 FILLER_60_376 ();
 FILLCELL_X2 FILLER_60_382 ();
 FILLCELL_X1 FILLER_60_384 ();
 FILLCELL_X1 FILLER_60_392 ();
 FILLCELL_X1 FILLER_60_409 ();
 FILLCELL_X2 FILLER_60_430 ();
 FILLCELL_X2 FILLER_60_446 ();
 FILLCELL_X1 FILLER_60_448 ();
 FILLCELL_X4 FILLER_60_459 ();
 FILLCELL_X1 FILLER_60_463 ();
 FILLCELL_X1 FILLER_60_473 ();
 FILLCELL_X1 FILLER_60_492 ();
 FILLCELL_X1 FILLER_60_527 ();
 FILLCELL_X1 FILLER_60_553 ();
 FILLCELL_X8 FILLER_60_564 ();
 FILLCELL_X1 FILLER_60_582 ();
 FILLCELL_X8 FILLER_60_611 ();
 FILLCELL_X4 FILLER_60_619 ();
 FILLCELL_X2 FILLER_60_623 ();
 FILLCELL_X4 FILLER_60_650 ();
 FILLCELL_X1 FILLER_60_654 ();
 FILLCELL_X2 FILLER_60_658 ();
 FILLCELL_X4 FILLER_60_665 ();
 FILLCELL_X4 FILLER_60_673 ();
 FILLCELL_X1 FILLER_60_677 ();
 FILLCELL_X4 FILLER_60_697 ();
 FILLCELL_X2 FILLER_60_701 ();
 FILLCELL_X16 FILLER_60_719 ();
 FILLCELL_X8 FILLER_60_735 ();
 FILLCELL_X2 FILLER_60_743 ();
 FILLCELL_X1 FILLER_60_745 ();
 FILLCELL_X16 FILLER_60_756 ();
 FILLCELL_X8 FILLER_60_772 ();
 FILLCELL_X2 FILLER_60_780 ();
 FILLCELL_X1 FILLER_60_782 ();
 FILLCELL_X16 FILLER_60_809 ();
 FILLCELL_X4 FILLER_60_825 ();
 FILLCELL_X2 FILLER_60_829 ();
 FILLCELL_X4 FILLER_60_883 ();
 FILLCELL_X4 FILLER_60_905 ();
 FILLCELL_X2 FILLER_60_909 ();
 FILLCELL_X8 FILLER_60_913 ();
 FILLCELL_X2 FILLER_60_921 ();
 FILLCELL_X16 FILLER_60_925 ();
 FILLCELL_X8 FILLER_60_941 ();
 FILLCELL_X1 FILLER_60_949 ();
 FILLCELL_X16 FILLER_60_963 ();
 FILLCELL_X2 FILLER_60_979 ();
 FILLCELL_X1 FILLER_60_981 ();
 FILLCELL_X16 FILLER_61_1 ();
 FILLCELL_X8 FILLER_61_17 ();
 FILLCELL_X4 FILLER_61_25 ();
 FILLCELL_X2 FILLER_61_29 ();
 FILLCELL_X1 FILLER_61_34 ();
 FILLCELL_X32 FILLER_61_38 ();
 FILLCELL_X8 FILLER_61_70 ();
 FILLCELL_X2 FILLER_61_78 ();
 FILLCELL_X8 FILLER_61_97 ();
 FILLCELL_X2 FILLER_61_125 ();
 FILLCELL_X1 FILLER_61_127 ();
 FILLCELL_X4 FILLER_61_148 ();
 FILLCELL_X1 FILLER_61_152 ();
 FILLCELL_X32 FILLER_61_170 ();
 FILLCELL_X16 FILLER_61_202 ();
 FILLCELL_X4 FILLER_61_218 ();
 FILLCELL_X2 FILLER_61_222 ();
 FILLCELL_X32 FILLER_61_227 ();
 FILLCELL_X16 FILLER_61_259 ();
 FILLCELL_X8 FILLER_61_275 ();
 FILLCELL_X1 FILLER_61_283 ();
 FILLCELL_X2 FILLER_61_364 ();
 FILLCELL_X1 FILLER_61_366 ();
 FILLCELL_X8 FILLER_61_377 ();
 FILLCELL_X2 FILLER_61_406 ();
 FILLCELL_X1 FILLER_61_408 ();
 FILLCELL_X4 FILLER_61_436 ();
 FILLCELL_X4 FILLER_61_522 ();
 FILLCELL_X1 FILLER_61_595 ();
 FILLCELL_X32 FILLER_61_605 ();
 FILLCELL_X32 FILLER_61_637 ();
 FILLCELL_X32 FILLER_61_669 ();
 FILLCELL_X2 FILLER_61_701 ();
 FILLCELL_X1 FILLER_61_703 ();
 FILLCELL_X16 FILLER_61_711 ();
 FILLCELL_X8 FILLER_61_727 ();
 FILLCELL_X2 FILLER_61_735 ();
 FILLCELL_X1 FILLER_61_737 ();
 FILLCELL_X8 FILLER_61_748 ();
 FILLCELL_X4 FILLER_61_756 ();
 FILLCELL_X2 FILLER_61_760 ();
 FILLCELL_X16 FILLER_61_764 ();
 FILLCELL_X2 FILLER_61_798 ();
 FILLCELL_X16 FILLER_61_802 ();
 FILLCELL_X4 FILLER_61_818 ();
 FILLCELL_X4 FILLER_61_824 ();
 FILLCELL_X2 FILLER_61_828 ();
 FILLCELL_X2 FILLER_61_832 ();
 FILLCELL_X16 FILLER_61_844 ();
 FILLCELL_X2 FILLER_61_860 ();
 FILLCELL_X2 FILLER_61_864 ();
 FILLCELL_X1 FILLER_61_866 ();
 FILLCELL_X4 FILLER_61_869 ();
 FILLCELL_X2 FILLER_61_873 ();
 FILLCELL_X1 FILLER_61_875 ();
 FILLCELL_X16 FILLER_61_878 ();
 FILLCELL_X2 FILLER_61_894 ();
 FILLCELL_X1 FILLER_61_896 ();
 FILLCELL_X8 FILLER_61_899 ();
 FILLCELL_X2 FILLER_61_907 ();
 FILLCELL_X8 FILLER_61_911 ();
 FILLCELL_X4 FILLER_61_919 ();
 FILLCELL_X2 FILLER_61_923 ();
 FILLCELL_X8 FILLER_61_927 ();
 FILLCELL_X4 FILLER_61_935 ();
 FILLCELL_X2 FILLER_61_939 ();
 FILLCELL_X8 FILLER_61_957 ();
 FILLCELL_X4 FILLER_61_965 ();
 FILLCELL_X2 FILLER_61_979 ();
 FILLCELL_X1 FILLER_61_981 ();
 FILLCELL_X32 FILLER_62_1 ();
 FILLCELL_X16 FILLER_62_33 ();
 FILLCELL_X8 FILLER_62_49 ();
 FILLCELL_X4 FILLER_62_57 ();
 FILLCELL_X4 FILLER_62_78 ();
 FILLCELL_X2 FILLER_62_82 ();
 FILLCELL_X1 FILLER_62_84 ();
 FILLCELL_X2 FILLER_62_88 ();
 FILLCELL_X1 FILLER_62_97 ();
 FILLCELL_X2 FILLER_62_101 ();
 FILLCELL_X2 FILLER_62_107 ();
 FILLCELL_X4 FILLER_62_116 ();
 FILLCELL_X4 FILLER_62_124 ();
 FILLCELL_X1 FILLER_62_128 ();
 FILLCELL_X4 FILLER_62_156 ();
 FILLCELL_X2 FILLER_62_160 ();
 FILLCELL_X1 FILLER_62_162 ();
 FILLCELL_X16 FILLER_62_168 ();
 FILLCELL_X8 FILLER_62_184 ();
 FILLCELL_X1 FILLER_62_212 ();
 FILLCELL_X1 FILLER_62_234 ();
 FILLCELL_X4 FILLER_62_239 ();
 FILLCELL_X1 FILLER_62_243 ();
 FILLCELL_X4 FILLER_62_247 ();
 FILLCELL_X2 FILLER_62_251 ();
 FILLCELL_X2 FILLER_62_257 ();
 FILLCELL_X1 FILLER_62_259 ();
 FILLCELL_X16 FILLER_62_263 ();
 FILLCELL_X32 FILLER_62_282 ();
 FILLCELL_X4 FILLER_62_314 ();
 FILLCELL_X1 FILLER_62_318 ();
 FILLCELL_X4 FILLER_62_347 ();
 FILLCELL_X1 FILLER_62_351 ();
 FILLCELL_X32 FILLER_62_361 ();
 FILLCELL_X4 FILLER_62_393 ();
 FILLCELL_X1 FILLER_62_397 ();
 FILLCELL_X8 FILLER_62_435 ();
 FILLCELL_X2 FILLER_62_443 ();
 FILLCELL_X1 FILLER_62_478 ();
 FILLCELL_X2 FILLER_62_497 ();
 FILLCELL_X2 FILLER_62_519 ();
 FILLCELL_X1 FILLER_62_525 ();
 FILLCELL_X2 FILLER_62_539 ();
 FILLCELL_X1 FILLER_62_541 ();
 FILLCELL_X32 FILLER_62_559 ();
 FILLCELL_X32 FILLER_62_591 ();
 FILLCELL_X8 FILLER_62_623 ();
 FILLCELL_X32 FILLER_62_632 ();
 FILLCELL_X32 FILLER_62_664 ();
 FILLCELL_X32 FILLER_62_696 ();
 FILLCELL_X1 FILLER_62_728 ();
 FILLCELL_X2 FILLER_62_745 ();
 FILLCELL_X32 FILLER_62_773 ();
 FILLCELL_X1 FILLER_62_805 ();
 FILLCELL_X8 FILLER_62_832 ();
 FILLCELL_X8 FILLER_62_878 ();
 FILLCELL_X4 FILLER_62_886 ();
 FILLCELL_X1 FILLER_62_890 ();
 FILLCELL_X4 FILLER_62_901 ();
 FILLCELL_X2 FILLER_62_905 ();
 FILLCELL_X1 FILLER_62_907 ();
 FILLCELL_X16 FILLER_62_924 ();
 FILLCELL_X8 FILLER_62_940 ();
 FILLCELL_X2 FILLER_62_948 ();
 FILLCELL_X8 FILLER_62_973 ();
 FILLCELL_X1 FILLER_62_981 ();
 FILLCELL_X4 FILLER_63_1 ();
 FILLCELL_X32 FILLER_63_8 ();
 FILLCELL_X16 FILLER_63_40 ();
 FILLCELL_X4 FILLER_63_56 ();
 FILLCELL_X2 FILLER_63_60 ();
 FILLCELL_X1 FILLER_63_62 ();
 FILLCELL_X2 FILLER_63_80 ();
 FILLCELL_X1 FILLER_63_82 ();
 FILLCELL_X1 FILLER_63_90 ();
 FILLCELL_X32 FILLER_63_95 ();
 FILLCELL_X2 FILLER_63_127 ();
 FILLCELL_X1 FILLER_63_129 ();
 FILLCELL_X8 FILLER_63_134 ();
 FILLCELL_X2 FILLER_63_142 ();
 FILLCELL_X16 FILLER_63_148 ();
 FILLCELL_X2 FILLER_63_164 ();
 FILLCELL_X1 FILLER_63_166 ();
 FILLCELL_X16 FILLER_63_172 ();
 FILLCELL_X8 FILLER_63_188 ();
 FILLCELL_X4 FILLER_63_196 ();
 FILLCELL_X2 FILLER_63_200 ();
 FILLCELL_X1 FILLER_63_202 ();
 FILLCELL_X8 FILLER_63_211 ();
 FILLCELL_X4 FILLER_63_219 ();
 FILLCELL_X1 FILLER_63_223 ();
 FILLCELL_X1 FILLER_63_228 ();
 FILLCELL_X2 FILLER_63_248 ();
 FILLCELL_X2 FILLER_63_269 ();
 FILLCELL_X32 FILLER_63_296 ();
 FILLCELL_X4 FILLER_63_328 ();
 FILLCELL_X2 FILLER_63_332 ();
 FILLCELL_X16 FILLER_63_339 ();
 FILLCELL_X1 FILLER_63_355 ();
 FILLCELL_X2 FILLER_63_379 ();
 FILLCELL_X1 FILLER_63_381 ();
 FILLCELL_X8 FILLER_63_401 ();
 FILLCELL_X4 FILLER_63_409 ();
 FILLCELL_X16 FILLER_63_417 ();
 FILLCELL_X8 FILLER_63_433 ();
 FILLCELL_X2 FILLER_63_441 ();
 FILLCELL_X32 FILLER_63_453 ();
 FILLCELL_X16 FILLER_63_485 ();
 FILLCELL_X4 FILLER_63_501 ();
 FILLCELL_X2 FILLER_63_505 ();
 FILLCELL_X1 FILLER_63_507 ();
 FILLCELL_X8 FILLER_63_518 ();
 FILLCELL_X4 FILLER_63_526 ();
 FILLCELL_X2 FILLER_63_530 ();
 FILLCELL_X1 FILLER_63_532 ();
 FILLCELL_X32 FILLER_63_542 ();
 FILLCELL_X32 FILLER_63_574 ();
 FILLCELL_X32 FILLER_63_606 ();
 FILLCELL_X32 FILLER_63_638 ();
 FILLCELL_X32 FILLER_63_670 ();
 FILLCELL_X32 FILLER_63_702 ();
 FILLCELL_X1 FILLER_63_734 ();
 FILLCELL_X2 FILLER_63_747 ();
 FILLCELL_X8 FILLER_63_759 ();
 FILLCELL_X8 FILLER_63_785 ();
 FILLCELL_X2 FILLER_63_793 ();
 FILLCELL_X1 FILLER_63_795 ();
 FILLCELL_X4 FILLER_63_830 ();
 FILLCELL_X2 FILLER_63_834 ();
 FILLCELL_X1 FILLER_63_836 ();
 FILLCELL_X4 FILLER_63_853 ();
 FILLCELL_X1 FILLER_63_857 ();
 FILLCELL_X4 FILLER_63_870 ();
 FILLCELL_X4 FILLER_63_876 ();
 FILLCELL_X1 FILLER_63_880 ();
 FILLCELL_X8 FILLER_63_901 ();
 FILLCELL_X2 FILLER_63_919 ();
 FILLCELL_X1 FILLER_63_921 ();
 FILLCELL_X8 FILLER_63_938 ();
 FILLCELL_X2 FILLER_63_946 ();
 FILLCELL_X1 FILLER_63_948 ();
 FILLCELL_X1 FILLER_63_965 ();
 FILLCELL_X2 FILLER_63_976 ();
 FILLCELL_X1 FILLER_63_978 ();
 FILLCELL_X8 FILLER_64_1 ();
 FILLCELL_X4 FILLER_64_9 ();
 FILLCELL_X2 FILLER_64_13 ();
 FILLCELL_X1 FILLER_64_15 ();
 FILLCELL_X32 FILLER_64_19 ();
 FILLCELL_X16 FILLER_64_51 ();
 FILLCELL_X4 FILLER_64_67 ();
 FILLCELL_X1 FILLER_64_71 ();
 FILLCELL_X8 FILLER_64_95 ();
 FILLCELL_X4 FILLER_64_103 ();
 FILLCELL_X1 FILLER_64_113 ();
 FILLCELL_X32 FILLER_64_138 ();
 FILLCELL_X2 FILLER_64_170 ();
 FILLCELL_X1 FILLER_64_172 ();
 FILLCELL_X1 FILLER_64_183 ();
 FILLCELL_X8 FILLER_64_198 ();
 FILLCELL_X1 FILLER_64_206 ();
 FILLCELL_X4 FILLER_64_209 ();
 FILLCELL_X2 FILLER_64_213 ();
 FILLCELL_X8 FILLER_64_218 ();
 FILLCELL_X4 FILLER_64_226 ();
 FILLCELL_X1 FILLER_64_230 ();
 FILLCELL_X16 FILLER_64_234 ();
 FILLCELL_X4 FILLER_64_269 ();
 FILLCELL_X1 FILLER_64_273 ();
 FILLCELL_X1 FILLER_64_279 ();
 FILLCELL_X32 FILLER_64_303 ();
 FILLCELL_X8 FILLER_64_335 ();
 FILLCELL_X4 FILLER_64_343 ();
 FILLCELL_X1 FILLER_64_347 ();
 FILLCELL_X8 FILLER_64_357 ();
 FILLCELL_X4 FILLER_64_365 ();
 FILLCELL_X1 FILLER_64_369 ();
 FILLCELL_X8 FILLER_64_374 ();
 FILLCELL_X1 FILLER_64_382 ();
 FILLCELL_X16 FILLER_64_389 ();
 FILLCELL_X4 FILLER_64_405 ();
 FILLCELL_X16 FILLER_64_431 ();
 FILLCELL_X1 FILLER_64_447 ();
 FILLCELL_X32 FILLER_64_464 ();
 FILLCELL_X8 FILLER_64_496 ();
 FILLCELL_X4 FILLER_64_504 ();
 FILLCELL_X32 FILLER_64_534 ();
 FILLCELL_X32 FILLER_64_566 ();
 FILLCELL_X32 FILLER_64_598 ();
 FILLCELL_X1 FILLER_64_630 ();
 FILLCELL_X32 FILLER_64_632 ();
 FILLCELL_X32 FILLER_64_664 ();
 FILLCELL_X32 FILLER_64_696 ();
 FILLCELL_X8 FILLER_64_728 ();
 FILLCELL_X4 FILLER_64_736 ();
 FILLCELL_X2 FILLER_64_740 ();
 FILLCELL_X1 FILLER_64_742 ();
 FILLCELL_X2 FILLER_64_745 ();
 FILLCELL_X1 FILLER_64_779 ();
 FILLCELL_X8 FILLER_64_796 ();
 FILLCELL_X1 FILLER_64_804 ();
 FILLCELL_X32 FILLER_64_807 ();
 FILLCELL_X32 FILLER_64_839 ();
 FILLCELL_X16 FILLER_64_871 ();
 FILLCELL_X1 FILLER_64_887 ();
 FILLCELL_X16 FILLER_64_900 ();
 FILLCELL_X16 FILLER_64_918 ();
 FILLCELL_X8 FILLER_64_934 ();
 FILLCELL_X4 FILLER_64_942 ();
 FILLCELL_X2 FILLER_64_958 ();
 FILLCELL_X1 FILLER_64_960 ();
 FILLCELL_X2 FILLER_64_964 ();
 FILLCELL_X1 FILLER_64_966 ();
 FILLCELL_X2 FILLER_64_973 ();
 FILLCELL_X1 FILLER_64_975 ();
 FILLCELL_X2 FILLER_64_979 ();
 FILLCELL_X1 FILLER_64_981 ();
 FILLCELL_X32 FILLER_65_1 ();
 FILLCELL_X16 FILLER_65_33 ();
 FILLCELL_X8 FILLER_65_49 ();
 FILLCELL_X2 FILLER_65_57 ();
 FILLCELL_X1 FILLER_65_59 ();
 FILLCELL_X16 FILLER_65_63 ();
 FILLCELL_X4 FILLER_65_79 ();
 FILLCELL_X1 FILLER_65_83 ();
 FILLCELL_X1 FILLER_65_114 ();
 FILLCELL_X2 FILLER_65_118 ();
 FILLCELL_X8 FILLER_65_123 ();
 FILLCELL_X4 FILLER_65_131 ();
 FILLCELL_X4 FILLER_65_138 ();
 FILLCELL_X2 FILLER_65_142 ();
 FILLCELL_X4 FILLER_65_147 ();
 FILLCELL_X1 FILLER_65_151 ();
 FILLCELL_X2 FILLER_65_155 ();
 FILLCELL_X4 FILLER_65_169 ();
 FILLCELL_X1 FILLER_65_173 ();
 FILLCELL_X2 FILLER_65_184 ();
 FILLCELL_X1 FILLER_65_186 ();
 FILLCELL_X4 FILLER_65_200 ();
 FILLCELL_X32 FILLER_65_227 ();
 FILLCELL_X1 FILLER_65_259 ();
 FILLCELL_X8 FILLER_65_272 ();
 FILLCELL_X2 FILLER_65_283 ();
 FILLCELL_X1 FILLER_65_312 ();
 FILLCELL_X4 FILLER_65_322 ();
 FILLCELL_X2 FILLER_65_326 ();
 FILLCELL_X1 FILLER_65_328 ();
 FILLCELL_X2 FILLER_65_373 ();
 FILLCELL_X1 FILLER_65_375 ();
 FILLCELL_X2 FILLER_65_381 ();
 FILLCELL_X8 FILLER_65_387 ();
 FILLCELL_X4 FILLER_65_395 ();
 FILLCELL_X2 FILLER_65_420 ();
 FILLCELL_X1 FILLER_65_422 ();
 FILLCELL_X16 FILLER_65_430 ();
 FILLCELL_X16 FILLER_65_452 ();
 FILLCELL_X1 FILLER_65_481 ();
 FILLCELL_X32 FILLER_65_485 ();
 FILLCELL_X32 FILLER_65_517 ();
 FILLCELL_X32 FILLER_65_549 ();
 FILLCELL_X32 FILLER_65_581 ();
 FILLCELL_X4 FILLER_65_613 ();
 FILLCELL_X4 FILLER_65_621 ();
 FILLCELL_X1 FILLER_65_625 ();
 FILLCELL_X2 FILLER_65_629 ();
 FILLCELL_X32 FILLER_65_636 ();
 FILLCELL_X32 FILLER_65_668 ();
 FILLCELL_X16 FILLER_65_700 ();
 FILLCELL_X8 FILLER_65_716 ();
 FILLCELL_X1 FILLER_65_724 ();
 FILLCELL_X1 FILLER_65_741 ();
 FILLCELL_X4 FILLER_65_752 ();
 FILLCELL_X2 FILLER_65_756 ();
 FILLCELL_X1 FILLER_65_758 ();
 FILLCELL_X16 FILLER_65_761 ();
 FILLCELL_X1 FILLER_65_777 ();
 FILLCELL_X4 FILLER_65_780 ();
 FILLCELL_X32 FILLER_65_800 ();
 FILLCELL_X16 FILLER_65_832 ();
 FILLCELL_X4 FILLER_65_848 ();
 FILLCELL_X1 FILLER_65_852 ();
 FILLCELL_X32 FILLER_65_879 ();
 FILLCELL_X4 FILLER_65_911 ();
 FILLCELL_X2 FILLER_65_915 ();
 FILLCELL_X4 FILLER_66_1 ();
 FILLCELL_X1 FILLER_66_5 ();
 FILLCELL_X16 FILLER_66_12 ();
 FILLCELL_X8 FILLER_66_31 ();
 FILLCELL_X4 FILLER_66_39 ();
 FILLCELL_X1 FILLER_66_43 ();
 FILLCELL_X8 FILLER_66_76 ();
 FILLCELL_X4 FILLER_66_84 ();
 FILLCELL_X2 FILLER_66_88 ();
 FILLCELL_X1 FILLER_66_90 ();
 FILLCELL_X4 FILLER_66_97 ();
 FILLCELL_X1 FILLER_66_101 ();
 FILLCELL_X2 FILLER_66_105 ();
 FILLCELL_X4 FILLER_66_113 ();
 FILLCELL_X1 FILLER_66_117 ();
 FILLCELL_X8 FILLER_66_123 ();
 FILLCELL_X4 FILLER_66_131 ();
 FILLCELL_X8 FILLER_66_143 ();
 FILLCELL_X4 FILLER_66_151 ();
 FILLCELL_X1 FILLER_66_155 ();
 FILLCELL_X2 FILLER_66_160 ();
 FILLCELL_X1 FILLER_66_162 ();
 FILLCELL_X1 FILLER_66_183 ();
 FILLCELL_X1 FILLER_66_197 ();
 FILLCELL_X8 FILLER_66_218 ();
 FILLCELL_X1 FILLER_66_226 ();
 FILLCELL_X4 FILLER_66_246 ();
 FILLCELL_X2 FILLER_66_250 ();
 FILLCELL_X1 FILLER_66_252 ();
 FILLCELL_X4 FILLER_66_256 ();
 FILLCELL_X16 FILLER_66_263 ();
 FILLCELL_X4 FILLER_66_279 ();
 FILLCELL_X2 FILLER_66_283 ();
 FILLCELL_X1 FILLER_66_285 ();
 FILLCELL_X16 FILLER_66_292 ();
 FILLCELL_X1 FILLER_66_315 ();
 FILLCELL_X8 FILLER_66_333 ();
 FILLCELL_X4 FILLER_66_341 ();
 FILLCELL_X1 FILLER_66_370 ();
 FILLCELL_X1 FILLER_66_386 ();
 FILLCELL_X1 FILLER_66_391 ();
 FILLCELL_X1 FILLER_66_399 ();
 FILLCELL_X2 FILLER_66_414 ();
 FILLCELL_X16 FILLER_66_423 ();
 FILLCELL_X4 FILLER_66_439 ();
 FILLCELL_X2 FILLER_66_443 ();
 FILLCELL_X1 FILLER_66_445 ();
 FILLCELL_X8 FILLER_66_452 ();
 FILLCELL_X4 FILLER_66_460 ();
 FILLCELL_X2 FILLER_66_464 ();
 FILLCELL_X1 FILLER_66_466 ();
 FILLCELL_X32 FILLER_66_491 ();
 FILLCELL_X8 FILLER_66_523 ();
 FILLCELL_X2 FILLER_66_531 ();
 FILLCELL_X32 FILLER_66_543 ();
 FILLCELL_X32 FILLER_66_575 ();
 FILLCELL_X4 FILLER_66_607 ();
 FILLCELL_X1 FILLER_66_611 ();
 FILLCELL_X8 FILLER_66_632 ();
 FILLCELL_X4 FILLER_66_640 ();
 FILLCELL_X32 FILLER_66_666 ();
 FILLCELL_X16 FILLER_66_698 ();
 FILLCELL_X2 FILLER_66_714 ();
 FILLCELL_X8 FILLER_66_732 ();
 FILLCELL_X4 FILLER_66_740 ();
 FILLCELL_X2 FILLER_66_744 ();
 FILLCELL_X1 FILLER_66_746 ();
 FILLCELL_X32 FILLER_66_749 ();
 FILLCELL_X8 FILLER_66_781 ();
 FILLCELL_X4 FILLER_66_789 ();
 FILLCELL_X2 FILLER_66_793 ();
 FILLCELL_X1 FILLER_66_815 ();
 FILLCELL_X16 FILLER_66_832 ();
 FILLCELL_X4 FILLER_66_864 ();
 FILLCELL_X2 FILLER_66_868 ();
 FILLCELL_X4 FILLER_66_886 ();
 FILLCELL_X2 FILLER_66_890 ();
 FILLCELL_X1 FILLER_66_892 ();
 FILLCELL_X16 FILLER_66_895 ();
 FILLCELL_X2 FILLER_66_911 ();
 FILLCELL_X1 FILLER_66_913 ();
 FILLCELL_X16 FILLER_66_932 ();
 FILLCELL_X8 FILLER_66_948 ();
 FILLCELL_X4 FILLER_66_972 ();
 FILLCELL_X1 FILLER_66_978 ();
 FILLCELL_X16 FILLER_67_1 ();
 FILLCELL_X4 FILLER_67_17 ();
 FILLCELL_X1 FILLER_67_21 ();
 FILLCELL_X16 FILLER_67_25 ();
 FILLCELL_X8 FILLER_67_41 ();
 FILLCELL_X4 FILLER_67_49 ();
 FILLCELL_X4 FILLER_67_74 ();
 FILLCELL_X1 FILLER_67_81 ();
 FILLCELL_X32 FILLER_67_86 ();
 FILLCELL_X16 FILLER_67_118 ();
 FILLCELL_X2 FILLER_67_165 ();
 FILLCELL_X1 FILLER_67_167 ();
 FILLCELL_X1 FILLER_67_178 ();
 FILLCELL_X16 FILLER_67_186 ();
 FILLCELL_X4 FILLER_67_202 ();
 FILLCELL_X2 FILLER_67_206 ();
 FILLCELL_X4 FILLER_67_241 ();
 FILLCELL_X1 FILLER_67_245 ();
 FILLCELL_X32 FILLER_67_256 ();
 FILLCELL_X8 FILLER_67_288 ();
 FILLCELL_X2 FILLER_67_296 ();
 FILLCELL_X1 FILLER_67_301 ();
 FILLCELL_X32 FILLER_67_321 ();
 FILLCELL_X4 FILLER_67_353 ();
 FILLCELL_X2 FILLER_67_357 ();
 FILLCELL_X1 FILLER_67_359 ();
 FILLCELL_X4 FILLER_67_364 ();
 FILLCELL_X2 FILLER_67_373 ();
 FILLCELL_X16 FILLER_67_409 ();
 FILLCELL_X1 FILLER_67_425 ();
 FILLCELL_X8 FILLER_67_436 ();
 FILLCELL_X2 FILLER_67_444 ();
 FILLCELL_X16 FILLER_67_468 ();
 FILLCELL_X16 FILLER_67_517 ();
 FILLCELL_X4 FILLER_67_533 ();
 FILLCELL_X32 FILLER_67_554 ();
 FILLCELL_X16 FILLER_67_586 ();
 FILLCELL_X8 FILLER_67_602 ();
 FILLCELL_X2 FILLER_67_610 ();
 FILLCELL_X8 FILLER_67_619 ();
 FILLCELL_X4 FILLER_67_627 ();
 FILLCELL_X2 FILLER_67_631 ();
 FILLCELL_X2 FILLER_67_663 ();
 FILLCELL_X32 FILLER_67_684 ();
 FILLCELL_X4 FILLER_67_716 ();
 FILLCELL_X2 FILLER_67_720 ();
 FILLCELL_X4 FILLER_67_728 ();
 FILLCELL_X8 FILLER_67_754 ();
 FILLCELL_X4 FILLER_67_762 ();
 FILLCELL_X2 FILLER_67_766 ();
 FILLCELL_X1 FILLER_67_768 ();
 FILLCELL_X2 FILLER_67_787 ();
 FILLCELL_X2 FILLER_67_791 ();
 FILLCELL_X8 FILLER_67_809 ();
 FILLCELL_X4 FILLER_67_817 ();
 FILLCELL_X8 FILLER_67_847 ();
 FILLCELL_X4 FILLER_67_855 ();
 FILLCELL_X2 FILLER_67_859 ();
 FILLCELL_X1 FILLER_67_861 ();
 FILLCELL_X1 FILLER_67_878 ();
 FILLCELL_X2 FILLER_67_889 ();
 FILLCELL_X1 FILLER_67_891 ();
 FILLCELL_X1 FILLER_67_894 ();
 FILLCELL_X8 FILLER_67_915 ();
 FILLCELL_X2 FILLER_67_923 ();
 FILLCELL_X4 FILLER_67_927 ();
 FILLCELL_X1 FILLER_67_931 ();
 FILLCELL_X4 FILLER_67_942 ();
 FILLCELL_X2 FILLER_67_946 ();
 FILLCELL_X1 FILLER_67_948 ();
 FILLCELL_X8 FILLER_67_969 ();
 FILLCELL_X4 FILLER_67_977 ();
 FILLCELL_X1 FILLER_67_981 ();
 FILLCELL_X32 FILLER_68_1 ();
 FILLCELL_X32 FILLER_68_33 ();
 FILLCELL_X4 FILLER_68_65 ();
 FILLCELL_X2 FILLER_68_69 ();
 FILLCELL_X32 FILLER_68_88 ();
 FILLCELL_X4 FILLER_68_120 ();
 FILLCELL_X2 FILLER_68_124 ();
 FILLCELL_X4 FILLER_68_131 ();
 FILLCELL_X2 FILLER_68_154 ();
 FILLCELL_X2 FILLER_68_168 ();
 FILLCELL_X2 FILLER_68_172 ();
 FILLCELL_X1 FILLER_68_174 ();
 FILLCELL_X1 FILLER_68_182 ();
 FILLCELL_X1 FILLER_68_197 ();
 FILLCELL_X1 FILLER_68_208 ();
 FILLCELL_X1 FILLER_68_216 ();
 FILLCELL_X2 FILLER_68_223 ();
 FILLCELL_X1 FILLER_68_225 ();
 FILLCELL_X4 FILLER_68_274 ();
 FILLCELL_X1 FILLER_68_278 ();
 FILLCELL_X1 FILLER_68_296 ();
 FILLCELL_X16 FILLER_68_316 ();
 FILLCELL_X2 FILLER_68_332 ();
 FILLCELL_X8 FILLER_68_343 ();
 FILLCELL_X4 FILLER_68_351 ();
 FILLCELL_X2 FILLER_68_355 ();
 FILLCELL_X1 FILLER_68_357 ();
 FILLCELL_X8 FILLER_68_361 ();
 FILLCELL_X2 FILLER_68_369 ();
 FILLCELL_X1 FILLER_68_371 ();
 FILLCELL_X2 FILLER_68_374 ();
 FILLCELL_X4 FILLER_68_389 ();
 FILLCELL_X2 FILLER_68_393 ();
 FILLCELL_X4 FILLER_68_419 ();
 FILLCELL_X1 FILLER_68_423 ();
 FILLCELL_X4 FILLER_68_443 ();
 FILLCELL_X2 FILLER_68_447 ();
 FILLCELL_X1 FILLER_68_449 ();
 FILLCELL_X8 FILLER_68_454 ();
 FILLCELL_X2 FILLER_68_462 ();
 FILLCELL_X1 FILLER_68_464 ();
 FILLCELL_X1 FILLER_68_491 ();
 FILLCELL_X2 FILLER_68_502 ();
 FILLCELL_X1 FILLER_68_504 ();
 FILLCELL_X4 FILLER_68_543 ();
 FILLCELL_X2 FILLER_68_547 ();
 FILLCELL_X32 FILLER_68_568 ();
 FILLCELL_X16 FILLER_68_600 ();
 FILLCELL_X2 FILLER_68_616 ();
 FILLCELL_X8 FILLER_68_621 ();
 FILLCELL_X2 FILLER_68_629 ();
 FILLCELL_X4 FILLER_68_632 ();
 FILLCELL_X4 FILLER_68_640 ();
 FILLCELL_X2 FILLER_68_644 ();
 FILLCELL_X8 FILLER_68_653 ();
 FILLCELL_X1 FILLER_68_661 ();
 FILLCELL_X1 FILLER_68_665 ();
 FILLCELL_X32 FILLER_68_670 ();
 FILLCELL_X8 FILLER_68_702 ();
 FILLCELL_X4 FILLER_68_710 ();
 FILLCELL_X2 FILLER_68_714 ();
 FILLCELL_X1 FILLER_68_716 ();
 FILLCELL_X2 FILLER_68_735 ();
 FILLCELL_X1 FILLER_68_737 ();
 FILLCELL_X2 FILLER_68_748 ();
 FILLCELL_X8 FILLER_68_782 ();
 FILLCELL_X4 FILLER_68_790 ();
 FILLCELL_X2 FILLER_68_794 ();
 FILLCELL_X8 FILLER_68_806 ();
 FILLCELL_X4 FILLER_68_814 ();
 FILLCELL_X2 FILLER_68_818 ();
 FILLCELL_X1 FILLER_68_823 ();
 FILLCELL_X8 FILLER_68_850 ();
 FILLCELL_X2 FILLER_68_858 ();
 FILLCELL_X1 FILLER_68_860 ();
 FILLCELL_X4 FILLER_68_887 ();
 FILLCELL_X2 FILLER_68_891 ();
 FILLCELL_X4 FILLER_68_905 ();
 FILLCELL_X1 FILLER_68_909 ();
 FILLCELL_X8 FILLER_68_940 ();
 FILLCELL_X2 FILLER_68_948 ();
 FILLCELL_X1 FILLER_68_950 ();
 FILLCELL_X2 FILLER_68_953 ();
 FILLCELL_X1 FILLER_68_955 ();
 FILLCELL_X8 FILLER_68_972 ();
 FILLCELL_X2 FILLER_68_980 ();
 FILLCELL_X8 FILLER_69_1 ();
 FILLCELL_X4 FILLER_69_9 ();
 FILLCELL_X16 FILLER_69_19 ();
 FILLCELL_X8 FILLER_69_35 ();
 FILLCELL_X2 FILLER_69_43 ();
 FILLCELL_X1 FILLER_69_45 ();
 FILLCELL_X32 FILLER_69_49 ();
 FILLCELL_X1 FILLER_69_81 ();
 FILLCELL_X8 FILLER_69_85 ();
 FILLCELL_X1 FILLER_69_98 ();
 FILLCELL_X2 FILLER_69_118 ();
 FILLCELL_X8 FILLER_69_139 ();
 FILLCELL_X4 FILLER_69_147 ();
 FILLCELL_X1 FILLER_69_151 ();
 FILLCELL_X8 FILLER_69_165 ();
 FILLCELL_X4 FILLER_69_173 ();
 FILLCELL_X2 FILLER_69_177 ();
 FILLCELL_X8 FILLER_69_190 ();
 FILLCELL_X1 FILLER_69_198 ();
 FILLCELL_X1 FILLER_69_223 ();
 FILLCELL_X8 FILLER_69_230 ();
 FILLCELL_X2 FILLER_69_238 ();
 FILLCELL_X8 FILLER_69_249 ();
 FILLCELL_X2 FILLER_69_257 ();
 FILLCELL_X1 FILLER_69_289 ();
 FILLCELL_X8 FILLER_69_319 ();
 FILLCELL_X4 FILLER_69_327 ();
 FILLCELL_X2 FILLER_69_331 ();
 FILLCELL_X1 FILLER_69_333 ();
 FILLCELL_X2 FILLER_69_351 ();
 FILLCELL_X16 FILLER_69_362 ();
 FILLCELL_X1 FILLER_69_378 ();
 FILLCELL_X2 FILLER_69_385 ();
 FILLCELL_X1 FILLER_69_387 ();
 FILLCELL_X4 FILLER_69_405 ();
 FILLCELL_X1 FILLER_69_409 ();
 FILLCELL_X8 FILLER_69_417 ();
 FILLCELL_X2 FILLER_69_425 ();
 FILLCELL_X1 FILLER_69_430 ();
 FILLCELL_X8 FILLER_69_435 ();
 FILLCELL_X4 FILLER_69_443 ();
 FILLCELL_X2 FILLER_69_447 ();
 FILLCELL_X8 FILLER_69_452 ();
 FILLCELL_X1 FILLER_69_460 ();
 FILLCELL_X1 FILLER_69_494 ();
 FILLCELL_X4 FILLER_69_509 ();
 FILLCELL_X32 FILLER_69_551 ();
 FILLCELL_X32 FILLER_69_583 ();
 FILLCELL_X16 FILLER_69_615 ();
 FILLCELL_X4 FILLER_69_631 ();
 FILLCELL_X32 FILLER_69_638 ();
 FILLCELL_X32 FILLER_69_670 ();
 FILLCELL_X32 FILLER_69_702 ();
 FILLCELL_X4 FILLER_69_734 ();
 FILLCELL_X2 FILLER_69_738 ();
 FILLCELL_X16 FILLER_69_742 ();
 FILLCELL_X4 FILLER_69_758 ();
 FILLCELL_X4 FILLER_69_794 ();
 FILLCELL_X8 FILLER_69_801 ();
 FILLCELL_X4 FILLER_69_809 ();
 FILLCELL_X1 FILLER_69_829 ();
 FILLCELL_X16 FILLER_69_865 ();
 FILLCELL_X4 FILLER_69_881 ();
 FILLCELL_X2 FILLER_69_885 ();
 FILLCELL_X8 FILLER_69_905 ();
 FILLCELL_X4 FILLER_69_913 ();
 FILLCELL_X2 FILLER_69_917 ();
 FILLCELL_X4 FILLER_69_929 ();
 FILLCELL_X1 FILLER_69_933 ();
 FILLCELL_X4 FILLER_69_950 ();
 FILLCELL_X2 FILLER_69_954 ();
 FILLCELL_X1 FILLER_69_956 ();
 FILLCELL_X8 FILLER_69_973 ();
 FILLCELL_X1 FILLER_69_981 ();
 FILLCELL_X16 FILLER_70_1 ();
 FILLCELL_X8 FILLER_70_17 ();
 FILLCELL_X2 FILLER_70_25 ();
 FILLCELL_X1 FILLER_70_27 ();
 FILLCELL_X8 FILLER_70_52 ();
 FILLCELL_X4 FILLER_70_60 ();
 FILLCELL_X4 FILLER_70_67 ();
 FILLCELL_X2 FILLER_70_71 ();
 FILLCELL_X8 FILLER_70_76 ();
 FILLCELL_X4 FILLER_70_84 ();
 FILLCELL_X1 FILLER_70_88 ();
 FILLCELL_X4 FILLER_70_95 ();
 FILLCELL_X2 FILLER_70_99 ();
 FILLCELL_X8 FILLER_70_120 ();
 FILLCELL_X8 FILLER_70_147 ();
 FILLCELL_X1 FILLER_70_166 ();
 FILLCELL_X4 FILLER_70_180 ();
 FILLCELL_X2 FILLER_70_184 ();
 FILLCELL_X1 FILLER_70_186 ();
 FILLCELL_X1 FILLER_70_224 ();
 FILLCELL_X1 FILLER_70_229 ();
 FILLCELL_X1 FILLER_70_256 ();
 FILLCELL_X1 FILLER_70_269 ();
 FILLCELL_X1 FILLER_70_277 ();
 FILLCELL_X8 FILLER_70_322 ();
 FILLCELL_X4 FILLER_70_330 ();
 FILLCELL_X2 FILLER_70_334 ();
 FILLCELL_X1 FILLER_70_336 ();
 FILLCELL_X2 FILLER_70_380 ();
 FILLCELL_X16 FILLER_70_401 ();
 FILLCELL_X8 FILLER_70_417 ();
 FILLCELL_X2 FILLER_70_425 ();
 FILLCELL_X1 FILLER_70_427 ();
 FILLCELL_X8 FILLER_70_452 ();
 FILLCELL_X4 FILLER_70_460 ();
 FILLCELL_X2 FILLER_70_464 ();
 FILLCELL_X1 FILLER_70_479 ();
 FILLCELL_X2 FILLER_70_500 ();
 FILLCELL_X1 FILLER_70_506 ();
 FILLCELL_X32 FILLER_70_540 ();
 FILLCELL_X32 FILLER_70_572 ();
 FILLCELL_X16 FILLER_70_604 ();
 FILLCELL_X8 FILLER_70_620 ();
 FILLCELL_X2 FILLER_70_628 ();
 FILLCELL_X1 FILLER_70_630 ();
 FILLCELL_X32 FILLER_70_632 ();
 FILLCELL_X32 FILLER_70_664 ();
 FILLCELL_X8 FILLER_70_696 ();
 FILLCELL_X4 FILLER_70_704 ();
 FILLCELL_X8 FILLER_70_724 ();
 FILLCELL_X1 FILLER_70_732 ();
 FILLCELL_X8 FILLER_70_749 ();
 FILLCELL_X4 FILLER_70_757 ();
 FILLCELL_X2 FILLER_70_761 ();
 FILLCELL_X1 FILLER_70_763 ();
 FILLCELL_X16 FILLER_70_766 ();
 FILLCELL_X8 FILLER_70_782 ();
 FILLCELL_X4 FILLER_70_792 ();
 FILLCELL_X16 FILLER_70_799 ();
 FILLCELL_X2 FILLER_70_815 ();
 FILLCELL_X1 FILLER_70_817 ();
 FILLCELL_X1 FILLER_70_820 ();
 FILLCELL_X8 FILLER_70_824 ();
 FILLCELL_X2 FILLER_70_832 ();
 FILLCELL_X1 FILLER_70_834 ();
 FILLCELL_X16 FILLER_70_845 ();
 FILLCELL_X16 FILLER_70_864 ();
 FILLCELL_X8 FILLER_70_880 ();
 FILLCELL_X4 FILLER_70_888 ();
 FILLCELL_X2 FILLER_70_892 ();
 FILLCELL_X1 FILLER_70_894 ();
 FILLCELL_X32 FILLER_70_913 ();
 FILLCELL_X8 FILLER_70_945 ();
 FILLCELL_X4 FILLER_70_953 ();
 FILLCELL_X8 FILLER_70_967 ();
 FILLCELL_X4 FILLER_70_975 ();
 FILLCELL_X2 FILLER_70_979 ();
 FILLCELL_X1 FILLER_70_981 ();
 FILLCELL_X16 FILLER_71_1 ();
 FILLCELL_X2 FILLER_71_17 ();
 FILLCELL_X1 FILLER_71_19 ();
 FILLCELL_X16 FILLER_71_28 ();
 FILLCELL_X2 FILLER_71_44 ();
 FILLCELL_X1 FILLER_71_46 ();
 FILLCELL_X8 FILLER_71_50 ();
 FILLCELL_X2 FILLER_71_58 ();
 FILLCELL_X16 FILLER_71_81 ();
 FILLCELL_X8 FILLER_71_97 ();
 FILLCELL_X2 FILLER_71_105 ();
 FILLCELL_X8 FILLER_71_126 ();
 FILLCELL_X4 FILLER_71_134 ();
 FILLCELL_X1 FILLER_71_138 ();
 FILLCELL_X2 FILLER_71_153 ();
 FILLCELL_X1 FILLER_71_155 ();
 FILLCELL_X16 FILLER_71_183 ();
 FILLCELL_X4 FILLER_71_199 ();
 FILLCELL_X1 FILLER_71_203 ();
 FILLCELL_X1 FILLER_71_214 ();
 FILLCELL_X4 FILLER_71_226 ();
 FILLCELL_X2 FILLER_71_230 ();
 FILLCELL_X4 FILLER_71_246 ();
 FILLCELL_X2 FILLER_71_250 ();
 FILLCELL_X1 FILLER_71_264 ();
 FILLCELL_X1 FILLER_71_268 ();
 FILLCELL_X8 FILLER_71_271 ();
 FILLCELL_X1 FILLER_71_283 ();
 FILLCELL_X1 FILLER_71_286 ();
 FILLCELL_X4 FILLER_71_290 ();
 FILLCELL_X16 FILLER_71_325 ();
 FILLCELL_X1 FILLER_71_341 ();
 FILLCELL_X2 FILLER_71_378 ();
 FILLCELL_X16 FILLER_71_383 ();
 FILLCELL_X16 FILLER_71_403 ();
 FILLCELL_X8 FILLER_71_419 ();
 FILLCELL_X2 FILLER_71_427 ();
 FILLCELL_X16 FILLER_71_446 ();
 FILLCELL_X4 FILLER_71_462 ();
 FILLCELL_X1 FILLER_71_466 ();
 FILLCELL_X1 FILLER_71_469 ();
 FILLCELL_X8 FILLER_71_495 ();
 FILLCELL_X4 FILLER_71_503 ();
 FILLCELL_X1 FILLER_71_507 ();
 FILLCELL_X1 FILLER_71_527 ();
 FILLCELL_X1 FILLER_71_540 ();
 FILLCELL_X1 FILLER_71_566 ();
 FILLCELL_X4 FILLER_71_577 ();
 FILLCELL_X2 FILLER_71_581 ();
 FILLCELL_X32 FILLER_71_589 ();
 FILLCELL_X32 FILLER_71_621 ();
 FILLCELL_X32 FILLER_71_653 ();
 FILLCELL_X16 FILLER_71_685 ();
 FILLCELL_X2 FILLER_71_701 ();
 FILLCELL_X1 FILLER_71_703 ();
 FILLCELL_X4 FILLER_71_726 ();
 FILLCELL_X2 FILLER_71_730 ();
 FILLCELL_X4 FILLER_71_754 ();
 FILLCELL_X1 FILLER_71_758 ();
 FILLCELL_X8 FILLER_71_771 ();
 FILLCELL_X4 FILLER_71_779 ();
 FILLCELL_X2 FILLER_71_793 ();
 FILLCELL_X4 FILLER_71_811 ();
 FILLCELL_X4 FILLER_71_825 ();
 FILLCELL_X2 FILLER_71_829 ();
 FILLCELL_X4 FILLER_71_857 ();
 FILLCELL_X1 FILLER_71_861 ();
 FILLCELL_X4 FILLER_71_865 ();
 FILLCELL_X8 FILLER_71_879 ();
 FILLCELL_X4 FILLER_71_903 ();
 FILLCELL_X1 FILLER_71_907 ();
 FILLCELL_X8 FILLER_71_922 ();
 FILLCELL_X2 FILLER_71_930 ();
 FILLCELL_X32 FILLER_71_942 ();
 FILLCELL_X8 FILLER_71_974 ();
 FILLCELL_X16 FILLER_72_1 ();
 FILLCELL_X8 FILLER_72_17 ();
 FILLCELL_X2 FILLER_72_25 ();
 FILLCELL_X32 FILLER_72_52 ();
 FILLCELL_X1 FILLER_72_84 ();
 FILLCELL_X8 FILLER_72_120 ();
 FILLCELL_X1 FILLER_72_128 ();
 FILLCELL_X4 FILLER_72_144 ();
 FILLCELL_X2 FILLER_72_148 ();
 FILLCELL_X1 FILLER_72_150 ();
 FILLCELL_X2 FILLER_72_171 ();
 FILLCELL_X16 FILLER_72_180 ();
 FILLCELL_X2 FILLER_72_196 ();
 FILLCELL_X1 FILLER_72_198 ();
 FILLCELL_X16 FILLER_72_201 ();
 FILLCELL_X4 FILLER_72_217 ();
 FILLCELL_X1 FILLER_72_221 ();
 FILLCELL_X16 FILLER_72_233 ();
 FILLCELL_X2 FILLER_72_249 ();
 FILLCELL_X4 FILLER_72_291 ();
 FILLCELL_X2 FILLER_72_295 ();
 FILLCELL_X2 FILLER_72_299 ();
 FILLCELL_X1 FILLER_72_301 ();
 FILLCELL_X2 FILLER_72_305 ();
 FILLCELL_X2 FILLER_72_317 ();
 FILLCELL_X1 FILLER_72_319 ();
 FILLCELL_X32 FILLER_72_323 ();
 FILLCELL_X4 FILLER_72_355 ();
 FILLCELL_X4 FILLER_72_367 ();
 FILLCELL_X2 FILLER_72_371 ();
 FILLCELL_X1 FILLER_72_373 ();
 FILLCELL_X2 FILLER_72_379 ();
 FILLCELL_X16 FILLER_72_398 ();
 FILLCELL_X8 FILLER_72_414 ();
 FILLCELL_X4 FILLER_72_422 ();
 FILLCELL_X16 FILLER_72_434 ();
 FILLCELL_X8 FILLER_72_450 ();
 FILLCELL_X2 FILLER_72_458 ();
 FILLCELL_X1 FILLER_72_494 ();
 FILLCELL_X4 FILLER_72_504 ();
 FILLCELL_X1 FILLER_72_508 ();
 FILLCELL_X4 FILLER_72_555 ();
 FILLCELL_X4 FILLER_72_602 ();
 FILLCELL_X2 FILLER_72_606 ();
 FILLCELL_X16 FILLER_72_615 ();
 FILLCELL_X32 FILLER_72_632 ();
 FILLCELL_X32 FILLER_72_664 ();
 FILLCELL_X8 FILLER_72_696 ();
 FILLCELL_X4 FILLER_72_704 ();
 FILLCELL_X2 FILLER_72_708 ();
 FILLCELL_X1 FILLER_72_710 ();
 FILLCELL_X8 FILLER_72_717 ();
 FILLCELL_X4 FILLER_72_725 ();
 FILLCELL_X2 FILLER_72_729 ();
 FILLCELL_X1 FILLER_72_731 ();
 FILLCELL_X32 FILLER_72_738 ();
 FILLCELL_X16 FILLER_72_770 ();
 FILLCELL_X4 FILLER_72_786 ();
 FILLCELL_X2 FILLER_72_790 ();
 FILLCELL_X2 FILLER_72_794 ();
 FILLCELL_X1 FILLER_72_796 ();
 FILLCELL_X1 FILLER_72_799 ();
 FILLCELL_X4 FILLER_72_802 ();
 FILLCELL_X2 FILLER_72_822 ();
 FILLCELL_X16 FILLER_72_840 ();
 FILLCELL_X4 FILLER_72_856 ();
 FILLCELL_X2 FILLER_72_876 ();
 FILLCELL_X1 FILLER_72_878 ();
 FILLCELL_X8 FILLER_72_895 ();
 FILLCELL_X4 FILLER_72_903 ();
 FILLCELL_X2 FILLER_72_919 ();
 FILLCELL_X8 FILLER_72_923 ();
 FILLCELL_X1 FILLER_72_931 ();
 FILLCELL_X1 FILLER_72_948 ();
 FILLCELL_X4 FILLER_72_975 ();
 FILLCELL_X2 FILLER_72_979 ();
 FILLCELL_X1 FILLER_72_981 ();
 FILLCELL_X4 FILLER_73_1 ();
 FILLCELL_X1 FILLER_73_5 ();
 FILLCELL_X8 FILLER_73_10 ();
 FILLCELL_X1 FILLER_73_18 ();
 FILLCELL_X8 FILLER_73_26 ();
 FILLCELL_X4 FILLER_73_34 ();
 FILLCELL_X2 FILLER_73_38 ();
 FILLCELL_X4 FILLER_73_44 ();
 FILLCELL_X1 FILLER_73_48 ();
 FILLCELL_X32 FILLER_73_52 ();
 FILLCELL_X4 FILLER_73_84 ();
 FILLCELL_X2 FILLER_73_88 ();
 FILLCELL_X16 FILLER_73_114 ();
 FILLCELL_X8 FILLER_73_130 ();
 FILLCELL_X1 FILLER_73_138 ();
 FILLCELL_X1 FILLER_73_157 ();
 FILLCELL_X16 FILLER_73_215 ();
 FILLCELL_X8 FILLER_73_231 ();
 FILLCELL_X1 FILLER_73_239 ();
 FILLCELL_X2 FILLER_73_242 ();
 FILLCELL_X16 FILLER_73_249 ();
 FILLCELL_X2 FILLER_73_265 ();
 FILLCELL_X1 FILLER_73_301 ();
 FILLCELL_X16 FILLER_73_320 ();
 FILLCELL_X1 FILLER_73_336 ();
 FILLCELL_X2 FILLER_73_341 ();
 FILLCELL_X1 FILLER_73_343 ();
 FILLCELL_X8 FILLER_73_379 ();
 FILLCELL_X4 FILLER_73_387 ();
 FILLCELL_X2 FILLER_73_391 ();
 FILLCELL_X1 FILLER_73_393 ();
 FILLCELL_X16 FILLER_73_399 ();
 FILLCELL_X8 FILLER_73_415 ();
 FILLCELL_X32 FILLER_73_427 ();
 FILLCELL_X8 FILLER_73_459 ();
 FILLCELL_X2 FILLER_73_467 ();
 FILLCELL_X1 FILLER_73_469 ();
 FILLCELL_X1 FILLER_73_490 ();
 FILLCELL_X8 FILLER_73_498 ();
 FILLCELL_X2 FILLER_73_506 ();
 FILLCELL_X1 FILLER_73_508 ();
 FILLCELL_X2 FILLER_73_516 ();
 FILLCELL_X1 FILLER_73_518 ();
 FILLCELL_X2 FILLER_73_546 ();
 FILLCELL_X1 FILLER_73_548 ();
 FILLCELL_X1 FILLER_73_584 ();
 FILLCELL_X32 FILLER_73_595 ();
 FILLCELL_X2 FILLER_73_627 ();
 FILLCELL_X1 FILLER_73_629 ();
 FILLCELL_X32 FILLER_73_637 ();
 FILLCELL_X32 FILLER_73_669 ();
 FILLCELL_X16 FILLER_73_701 ();
 FILLCELL_X8 FILLER_73_717 ();
 FILLCELL_X4 FILLER_73_725 ();
 FILLCELL_X2 FILLER_73_729 ();
 FILLCELL_X1 FILLER_73_731 ();
 FILLCELL_X8 FILLER_73_742 ();
 FILLCELL_X2 FILLER_73_750 ();
 FILLCELL_X1 FILLER_73_752 ();
 FILLCELL_X8 FILLER_73_769 ();
 FILLCELL_X4 FILLER_73_777 ();
 FILLCELL_X1 FILLER_73_781 ();
 FILLCELL_X16 FILLER_73_800 ();
 FILLCELL_X2 FILLER_73_816 ();
 FILLCELL_X8 FILLER_73_834 ();
 FILLCELL_X2 FILLER_73_842 ();
 FILLCELL_X32 FILLER_73_846 ();
 FILLCELL_X32 FILLER_73_878 ();
 FILLCELL_X16 FILLER_73_910 ();
 FILLCELL_X4 FILLER_73_926 ();
 FILLCELL_X1 FILLER_73_930 ();
 FILLCELL_X4 FILLER_73_941 ();
 FILLCELL_X2 FILLER_73_945 ();
 FILLCELL_X1 FILLER_73_954 ();
 FILLCELL_X2 FILLER_73_957 ();
 FILLCELL_X1 FILLER_73_981 ();
 FILLCELL_X2 FILLER_74_1 ();
 FILLCELL_X16 FILLER_74_7 ();
 FILLCELL_X2 FILLER_74_23 ();
 FILLCELL_X1 FILLER_74_25 ();
 FILLCELL_X4 FILLER_74_30 ();
 FILLCELL_X8 FILLER_74_55 ();
 FILLCELL_X4 FILLER_74_63 ();
 FILLCELL_X2 FILLER_74_67 ();
 FILLCELL_X1 FILLER_74_69 ();
 FILLCELL_X4 FILLER_74_73 ();
 FILLCELL_X2 FILLER_74_77 ();
 FILLCELL_X4 FILLER_74_109 ();
 FILLCELL_X2 FILLER_74_113 ();
 FILLCELL_X1 FILLER_74_115 ();
 FILLCELL_X1 FILLER_74_136 ();
 FILLCELL_X2 FILLER_74_162 ();
 FILLCELL_X1 FILLER_74_174 ();
 FILLCELL_X2 FILLER_74_227 ();
 FILLCELL_X1 FILLER_74_229 ();
 FILLCELL_X16 FILLER_74_249 ();
 FILLCELL_X2 FILLER_74_265 ();
 FILLCELL_X2 FILLER_74_279 ();
 FILLCELL_X1 FILLER_74_281 ();
 FILLCELL_X1 FILLER_74_291 ();
 FILLCELL_X1 FILLER_74_297 ();
 FILLCELL_X1 FILLER_74_302 ();
 FILLCELL_X16 FILLER_74_319 ();
 FILLCELL_X8 FILLER_74_335 ();
 FILLCELL_X1 FILLER_74_362 ();
 FILLCELL_X4 FILLER_74_367 ();
 FILLCELL_X4 FILLER_74_395 ();
 FILLCELL_X1 FILLER_74_399 ();
 FILLCELL_X2 FILLER_74_417 ();
 FILLCELL_X2 FILLER_74_444 ();
 FILLCELL_X8 FILLER_74_463 ();
 FILLCELL_X4 FILLER_74_471 ();
 FILLCELL_X2 FILLER_74_475 ();
 FILLCELL_X1 FILLER_74_483 ();
 FILLCELL_X4 FILLER_74_514 ();
 FILLCELL_X1 FILLER_74_518 ();
 FILLCELL_X4 FILLER_74_540 ();
 FILLCELL_X2 FILLER_74_544 ();
 FILLCELL_X1 FILLER_74_546 ();
 FILLCELL_X4 FILLER_74_557 ();
 FILLCELL_X32 FILLER_74_597 ();
 FILLCELL_X2 FILLER_74_629 ();
 FILLCELL_X32 FILLER_74_632 ();
 FILLCELL_X32 FILLER_74_664 ();
 FILLCELL_X16 FILLER_74_696 ();
 FILLCELL_X8 FILLER_74_712 ();
 FILLCELL_X4 FILLER_74_720 ();
 FILLCELL_X1 FILLER_74_724 ();
 FILLCELL_X1 FILLER_74_731 ();
 FILLCELL_X4 FILLER_74_746 ();
 FILLCELL_X1 FILLER_74_750 ();
 FILLCELL_X16 FILLER_74_755 ();
 FILLCELL_X1 FILLER_74_771 ();
 FILLCELL_X2 FILLER_74_790 ();
 FILLCELL_X32 FILLER_74_794 ();
 FILLCELL_X32 FILLER_74_826 ();
 FILLCELL_X4 FILLER_74_858 ();
 FILLCELL_X2 FILLER_74_862 ();
 FILLCELL_X1 FILLER_74_867 ();
 FILLCELL_X4 FILLER_74_883 ();
 FILLCELL_X1 FILLER_74_887 ();
 FILLCELL_X4 FILLER_74_904 ();
 FILLCELL_X2 FILLER_74_908 ();
 FILLCELL_X1 FILLER_74_910 ();
 FILLCELL_X2 FILLER_74_921 ();
 FILLCELL_X1 FILLER_74_933 ();
 FILLCELL_X16 FILLER_74_946 ();
 FILLCELL_X1 FILLER_74_962 ();
 FILLCELL_X8 FILLER_74_968 ();
 FILLCELL_X4 FILLER_74_976 ();
 FILLCELL_X2 FILLER_74_980 ();
 FILLCELL_X8 FILLER_75_1 ();
 FILLCELL_X8 FILLER_75_13 ();
 FILLCELL_X4 FILLER_75_21 ();
 FILLCELL_X2 FILLER_75_25 ();
 FILLCELL_X4 FILLER_75_31 ();
 FILLCELL_X2 FILLER_75_35 ();
 FILLCELL_X1 FILLER_75_37 ();
 FILLCELL_X16 FILLER_75_42 ();
 FILLCELL_X8 FILLER_75_58 ();
 FILLCELL_X1 FILLER_75_66 ();
 FILLCELL_X32 FILLER_75_111 ();
 FILLCELL_X1 FILLER_75_143 ();
 FILLCELL_X4 FILLER_75_172 ();
 FILLCELL_X1 FILLER_75_219 ();
 FILLCELL_X8 FILLER_75_229 ();
 FILLCELL_X1 FILLER_75_237 ();
 FILLCELL_X4 FILLER_75_248 ();
 FILLCELL_X16 FILLER_75_258 ();
 FILLCELL_X8 FILLER_75_274 ();
 FILLCELL_X4 FILLER_75_282 ();
 FILLCELL_X16 FILLER_75_300 ();
 FILLCELL_X4 FILLER_75_316 ();
 FILLCELL_X1 FILLER_75_320 ();
 FILLCELL_X8 FILLER_75_347 ();
 FILLCELL_X4 FILLER_75_355 ();
 FILLCELL_X8 FILLER_75_363 ();
 FILLCELL_X4 FILLER_75_371 ();
 FILLCELL_X2 FILLER_75_375 ();
 FILLCELL_X1 FILLER_75_377 ();
 FILLCELL_X4 FILLER_75_387 ();
 FILLCELL_X2 FILLER_75_401 ();
 FILLCELL_X1 FILLER_75_403 ();
 FILLCELL_X2 FILLER_75_451 ();
 FILLCELL_X1 FILLER_75_453 ();
 FILLCELL_X2 FILLER_75_474 ();
 FILLCELL_X1 FILLER_75_488 ();
 FILLCELL_X32 FILLER_75_498 ();
 FILLCELL_X1 FILLER_75_530 ();
 FILLCELL_X32 FILLER_75_538 ();
 FILLCELL_X4 FILLER_75_570 ();
 FILLCELL_X2 FILLER_75_574 ();
 FILLCELL_X1 FILLER_75_576 ();
 FILLCELL_X32 FILLER_75_603 ();
 FILLCELL_X16 FILLER_75_635 ();
 FILLCELL_X8 FILLER_75_651 ();
 FILLCELL_X2 FILLER_75_659 ();
 FILLCELL_X16 FILLER_75_711 ();
 FILLCELL_X2 FILLER_75_789 ();
 FILLCELL_X1 FILLER_75_791 ();
 FILLCELL_X4 FILLER_75_818 ();
 FILLCELL_X2 FILLER_75_838 ();
 FILLCELL_X1 FILLER_75_840 ();
 FILLCELL_X4 FILLER_75_860 ();
 FILLCELL_X2 FILLER_75_864 ();
 FILLCELL_X1 FILLER_75_866 ();
 FILLCELL_X4 FILLER_75_870 ();
 FILLCELL_X1 FILLER_75_874 ();
 FILLCELL_X8 FILLER_75_878 ();
 FILLCELL_X2 FILLER_75_886 ();
 FILLCELL_X1 FILLER_75_888 ();
 FILLCELL_X1 FILLER_75_891 ();
 FILLCELL_X1 FILLER_75_908 ();
 FILLCELL_X8 FILLER_75_927 ();
 FILLCELL_X1 FILLER_75_935 ();
 FILLCELL_X1 FILLER_75_946 ();
 FILLCELL_X2 FILLER_75_963 ();
 FILLCELL_X8 FILLER_75_967 ();
 FILLCELL_X4 FILLER_75_975 ();
 FILLCELL_X2 FILLER_75_979 ();
 FILLCELL_X1 FILLER_75_981 ();
 FILLCELL_X8 FILLER_76_1 ();
 FILLCELL_X2 FILLER_76_9 ();
 FILLCELL_X1 FILLER_76_11 ();
 FILLCELL_X4 FILLER_76_16 ();
 FILLCELL_X2 FILLER_76_24 ();
 FILLCELL_X32 FILLER_76_30 ();
 FILLCELL_X4 FILLER_76_62 ();
 FILLCELL_X2 FILLER_76_66 ();
 FILLCELL_X1 FILLER_76_68 ();
 FILLCELL_X1 FILLER_76_77 ();
 FILLCELL_X2 FILLER_76_108 ();
 FILLCELL_X1 FILLER_76_110 ();
 FILLCELL_X8 FILLER_76_130 ();
 FILLCELL_X4 FILLER_76_138 ();
 FILLCELL_X2 FILLER_76_142 ();
 FILLCELL_X2 FILLER_76_191 ();
 FILLCELL_X1 FILLER_76_226 ();
 FILLCELL_X2 FILLER_76_237 ();
 FILLCELL_X2 FILLER_76_252 ();
 FILLCELL_X2 FILLER_76_271 ();
 FILLCELL_X1 FILLER_76_273 ();
 FILLCELL_X2 FILLER_76_285 ();
 FILLCELL_X1 FILLER_76_307 ();
 FILLCELL_X8 FILLER_76_342 ();
 FILLCELL_X4 FILLER_76_350 ();
 FILLCELL_X2 FILLER_76_354 ();
 FILLCELL_X4 FILLER_76_388 ();
 FILLCELL_X2 FILLER_76_392 ();
 FILLCELL_X1 FILLER_76_394 ();
 FILLCELL_X2 FILLER_76_398 ();
 FILLCELL_X4 FILLER_76_422 ();
 FILLCELL_X1 FILLER_76_426 ();
 FILLCELL_X4 FILLER_76_437 ();
 FILLCELL_X1 FILLER_76_441 ();
 FILLCELL_X4 FILLER_76_446 ();
 FILLCELL_X2 FILLER_76_450 ();
 FILLCELL_X1 FILLER_76_469 ();
 FILLCELL_X32 FILLER_76_508 ();
 FILLCELL_X16 FILLER_76_540 ();
 FILLCELL_X4 FILLER_76_556 ();
 FILLCELL_X2 FILLER_76_560 ();
 FILLCELL_X1 FILLER_76_572 ();
 FILLCELL_X1 FILLER_76_575 ();
 FILLCELL_X2 FILLER_76_589 ();
 FILLCELL_X2 FILLER_76_601 ();
 FILLCELL_X16 FILLER_76_611 ();
 FILLCELL_X4 FILLER_76_627 ();
 FILLCELL_X16 FILLER_76_632 ();
 FILLCELL_X4 FILLER_76_648 ();
 FILLCELL_X1 FILLER_76_652 ();
 FILLCELL_X4 FILLER_76_675 ();
 FILLCELL_X2 FILLER_76_679 ();
 FILLCELL_X16 FILLER_76_684 ();
 FILLCELL_X8 FILLER_76_700 ();
 FILLCELL_X4 FILLER_76_708 ();
 FILLCELL_X2 FILLER_76_712 ();
 FILLCELL_X1 FILLER_76_714 ();
 FILLCELL_X8 FILLER_76_721 ();
 FILLCELL_X2 FILLER_76_729 ();
 FILLCELL_X1 FILLER_76_731 ();
 FILLCELL_X8 FILLER_76_754 ();
 FILLCELL_X1 FILLER_76_762 ();
 FILLCELL_X8 FILLER_76_765 ();
 FILLCELL_X8 FILLER_76_789 ();
 FILLCELL_X1 FILLER_76_797 ();
 FILLCELL_X4 FILLER_76_832 ();
 FILLCELL_X16 FILLER_76_862 ();
 FILLCELL_X8 FILLER_76_878 ();
 FILLCELL_X1 FILLER_76_886 ();
 FILLCELL_X2 FILLER_76_897 ();
 FILLCELL_X8 FILLER_76_917 ();
 FILLCELL_X2 FILLER_76_927 ();
 FILLCELL_X32 FILLER_76_939 ();
 FILLCELL_X8 FILLER_76_971 ();
 FILLCELL_X2 FILLER_76_979 ();
 FILLCELL_X1 FILLER_76_981 ();
 FILLCELL_X16 FILLER_77_4 ();
 FILLCELL_X1 FILLER_77_20 ();
 FILLCELL_X4 FILLER_77_24 ();
 FILLCELL_X2 FILLER_77_28 ();
 FILLCELL_X8 FILLER_77_57 ();
 FILLCELL_X2 FILLER_77_65 ();
 FILLCELL_X8 FILLER_77_86 ();
 FILLCELL_X4 FILLER_77_94 ();
 FILLCELL_X2 FILLER_77_98 ();
 FILLCELL_X2 FILLER_77_111 ();
 FILLCELL_X16 FILLER_77_133 ();
 FILLCELL_X8 FILLER_77_149 ();
 FILLCELL_X4 FILLER_77_157 ();
 FILLCELL_X1 FILLER_77_166 ();
 FILLCELL_X1 FILLER_77_177 ();
 FILLCELL_X1 FILLER_77_188 ();
 FILLCELL_X2 FILLER_77_221 ();
 FILLCELL_X2 FILLER_77_230 ();
 FILLCELL_X2 FILLER_77_237 ();
 FILLCELL_X1 FILLER_77_239 ();
 FILLCELL_X2 FILLER_77_253 ();
 FILLCELL_X1 FILLER_77_255 ();
 FILLCELL_X2 FILLER_77_273 ();
 FILLCELL_X1 FILLER_77_275 ();
 FILLCELL_X2 FILLER_77_286 ();
 FILLCELL_X16 FILLER_77_301 ();
 FILLCELL_X4 FILLER_77_317 ();
 FILLCELL_X4 FILLER_77_326 ();
 FILLCELL_X1 FILLER_77_330 ();
 FILLCELL_X16 FILLER_77_344 ();
 FILLCELL_X8 FILLER_77_360 ();
 FILLCELL_X1 FILLER_77_368 ();
 FILLCELL_X8 FILLER_77_390 ();
 FILLCELL_X2 FILLER_77_398 ();
 FILLCELL_X2 FILLER_77_407 ();
 FILLCELL_X8 FILLER_77_418 ();
 FILLCELL_X2 FILLER_77_426 ();
 FILLCELL_X8 FILLER_77_444 ();
 FILLCELL_X2 FILLER_77_452 ();
 FILLCELL_X8 FILLER_77_471 ();
 FILLCELL_X4 FILLER_77_479 ();
 FILLCELL_X1 FILLER_77_483 ();
 FILLCELL_X4 FILLER_77_509 ();
 FILLCELL_X2 FILLER_77_538 ();
 FILLCELL_X1 FILLER_77_540 ();
 FILLCELL_X16 FILLER_77_545 ();
 FILLCELL_X1 FILLER_77_561 ();
 FILLCELL_X2 FILLER_77_592 ();
 FILLCELL_X1 FILLER_77_594 ();
 FILLCELL_X2 FILLER_77_618 ();
 FILLCELL_X1 FILLER_77_620 ();
 FILLCELL_X8 FILLER_77_640 ();
 FILLCELL_X4 FILLER_77_648 ();
 FILLCELL_X1 FILLER_77_652 ();
 FILLCELL_X1 FILLER_77_656 ();
 FILLCELL_X8 FILLER_77_661 ();
 FILLCELL_X8 FILLER_77_673 ();
 FILLCELL_X1 FILLER_77_681 ();
 FILLCELL_X8 FILLER_77_704 ();
 FILLCELL_X1 FILLER_77_712 ();
 FILLCELL_X2 FILLER_77_731 ();
 FILLCELL_X16 FILLER_77_739 ();
 FILLCELL_X4 FILLER_77_755 ();
 FILLCELL_X1 FILLER_77_759 ();
 FILLCELL_X8 FILLER_77_766 ();
 FILLCELL_X4 FILLER_77_774 ();
 FILLCELL_X2 FILLER_77_778 ();
 FILLCELL_X1 FILLER_77_780 ();
 FILLCELL_X32 FILLER_77_799 ();
 FILLCELL_X8 FILLER_77_831 ();
 FILLCELL_X8 FILLER_77_844 ();
 FILLCELL_X2 FILLER_77_852 ();
 FILLCELL_X1 FILLER_77_854 ();
 FILLCELL_X2 FILLER_77_873 ();
 FILLCELL_X4 FILLER_77_883 ();
 FILLCELL_X2 FILLER_77_887 ();
 FILLCELL_X1 FILLER_77_892 ();
 FILLCELL_X2 FILLER_77_896 ();
 FILLCELL_X8 FILLER_77_908 ();
 FILLCELL_X16 FILLER_77_918 ();
 FILLCELL_X4 FILLER_77_934 ();
 FILLCELL_X16 FILLER_77_956 ();
 FILLCELL_X8 FILLER_77_972 ();
 FILLCELL_X2 FILLER_77_980 ();
 FILLCELL_X4 FILLER_78_1 ();
 FILLCELL_X2 FILLER_78_5 ();
 FILLCELL_X16 FILLER_78_11 ();
 FILLCELL_X1 FILLER_78_27 ();
 FILLCELL_X4 FILLER_78_49 ();
 FILLCELL_X2 FILLER_78_53 ();
 FILLCELL_X4 FILLER_78_59 ();
 FILLCELL_X2 FILLER_78_63 ();
 FILLCELL_X16 FILLER_78_68 ();
 FILLCELL_X8 FILLER_78_84 ();
 FILLCELL_X4 FILLER_78_92 ();
 FILLCELL_X16 FILLER_78_118 ();
 FILLCELL_X8 FILLER_78_134 ();
 FILLCELL_X4 FILLER_78_181 ();
 FILLCELL_X2 FILLER_78_202 ();
 FILLCELL_X8 FILLER_78_217 ();
 FILLCELL_X1 FILLER_78_225 ();
 FILLCELL_X32 FILLER_78_236 ();
 FILLCELL_X4 FILLER_78_268 ();
 FILLCELL_X2 FILLER_78_272 ();
 FILLCELL_X1 FILLER_78_274 ();
 FILLCELL_X2 FILLER_78_282 ();
 FILLCELL_X1 FILLER_78_284 ();
 FILLCELL_X2 FILLER_78_302 ();
 FILLCELL_X2 FILLER_78_321 ();
 FILLCELL_X1 FILLER_78_323 ();
 FILLCELL_X16 FILLER_78_346 ();
 FILLCELL_X4 FILLER_78_362 ();
 FILLCELL_X2 FILLER_78_366 ();
 FILLCELL_X16 FILLER_78_387 ();
 FILLCELL_X4 FILLER_78_403 ();
 FILLCELL_X2 FILLER_78_407 ();
 FILLCELL_X1 FILLER_78_409 ();
 FILLCELL_X16 FILLER_78_412 ();
 FILLCELL_X1 FILLER_78_428 ();
 FILLCELL_X4 FILLER_78_457 ();
 FILLCELL_X1 FILLER_78_461 ();
 FILLCELL_X8 FILLER_78_467 ();
 FILLCELL_X4 FILLER_78_475 ();
 FILLCELL_X1 FILLER_78_502 ();
 FILLCELL_X2 FILLER_78_543 ();
 FILLCELL_X1 FILLER_78_562 ();
 FILLCELL_X1 FILLER_78_586 ();
 FILLCELL_X16 FILLER_78_614 ();
 FILLCELL_X1 FILLER_78_630 ();
 FILLCELL_X16 FILLER_78_632 ();
 FILLCELL_X2 FILLER_78_648 ();
 FILLCELL_X1 FILLER_78_650 ();
 FILLCELL_X2 FILLER_78_656 ();
 FILLCELL_X1 FILLER_78_658 ();
 FILLCELL_X16 FILLER_78_662 ();
 FILLCELL_X4 FILLER_78_678 ();
 FILLCELL_X2 FILLER_78_682 ();
 FILLCELL_X32 FILLER_78_688 ();
 FILLCELL_X8 FILLER_78_720 ();
 FILLCELL_X1 FILLER_78_728 ();
 FILLCELL_X2 FILLER_78_735 ();
 FILLCELL_X16 FILLER_78_761 ();
 FILLCELL_X2 FILLER_78_777 ();
 FILLCELL_X8 FILLER_78_795 ();
 FILLCELL_X8 FILLER_78_809 ();
 FILLCELL_X2 FILLER_78_817 ();
 FILLCELL_X1 FILLER_78_819 ();
 FILLCELL_X4 FILLER_78_841 ();
 FILLCELL_X2 FILLER_78_845 ();
 FILLCELL_X2 FILLER_78_850 ();
 FILLCELL_X1 FILLER_78_852 ();
 FILLCELL_X2 FILLER_78_857 ();
 FILLCELL_X1 FILLER_78_862 ();
 FILLCELL_X2 FILLER_78_891 ();
 FILLCELL_X1 FILLER_78_893 ();
 FILLCELL_X16 FILLER_78_913 ();
 FILLCELL_X4 FILLER_78_929 ();
 FILLCELL_X1 FILLER_78_933 ();
 FILLCELL_X16 FILLER_78_936 ();
 FILLCELL_X1 FILLER_78_952 ();
 FILLCELL_X16 FILLER_78_955 ();
 FILLCELL_X8 FILLER_78_971 ();
 FILLCELL_X2 FILLER_78_979 ();
 FILLCELL_X1 FILLER_78_981 ();
 FILLCELL_X16 FILLER_79_1 ();
 FILLCELL_X4 FILLER_79_17 ();
 FILLCELL_X1 FILLER_79_21 ();
 FILLCELL_X32 FILLER_79_33 ();
 FILLCELL_X4 FILLER_79_65 ();
 FILLCELL_X2 FILLER_79_69 ();
 FILLCELL_X32 FILLER_79_85 ();
 FILLCELL_X16 FILLER_79_117 ();
 FILLCELL_X2 FILLER_79_133 ();
 FILLCELL_X1 FILLER_79_135 ();
 FILLCELL_X2 FILLER_79_168 ();
 FILLCELL_X1 FILLER_79_170 ();
 FILLCELL_X2 FILLER_79_178 ();
 FILLCELL_X1 FILLER_79_180 ();
 FILLCELL_X16 FILLER_79_198 ();
 FILLCELL_X4 FILLER_79_214 ();
 FILLCELL_X1 FILLER_79_218 ();
 FILLCELL_X8 FILLER_79_236 ();
 FILLCELL_X4 FILLER_79_244 ();
 FILLCELL_X1 FILLER_79_248 ();
 FILLCELL_X16 FILLER_79_252 ();
 FILLCELL_X4 FILLER_79_268 ();
 FILLCELL_X2 FILLER_79_272 ();
 FILLCELL_X1 FILLER_79_274 ();
 FILLCELL_X4 FILLER_79_288 ();
 FILLCELL_X4 FILLER_79_301 ();
 FILLCELL_X2 FILLER_79_305 ();
 FILLCELL_X8 FILLER_79_312 ();
 FILLCELL_X4 FILLER_79_320 ();
 FILLCELL_X2 FILLER_79_324 ();
 FILLCELL_X4 FILLER_79_346 ();
 FILLCELL_X16 FILLER_79_359 ();
 FILLCELL_X2 FILLER_79_375 ();
 FILLCELL_X8 FILLER_79_389 ();
 FILLCELL_X16 FILLER_79_420 ();
 FILLCELL_X1 FILLER_79_436 ();
 FILLCELL_X1 FILLER_79_450 ();
 FILLCELL_X2 FILLER_79_458 ();
 FILLCELL_X2 FILLER_79_463 ();
 FILLCELL_X1 FILLER_79_495 ();
 FILLCELL_X1 FILLER_79_536 ();
 FILLCELL_X4 FILLER_79_556 ();
 FILLCELL_X2 FILLER_79_560 ();
 FILLCELL_X1 FILLER_79_562 ();
 FILLCELL_X2 FILLER_79_566 ();
 FILLCELL_X4 FILLER_79_577 ();
 FILLCELL_X2 FILLER_79_591 ();
 FILLCELL_X32 FILLER_79_611 ();
 FILLCELL_X8 FILLER_79_643 ();
 FILLCELL_X4 FILLER_79_651 ();
 FILLCELL_X1 FILLER_79_655 ();
 FILLCELL_X32 FILLER_79_664 ();
 FILLCELL_X8 FILLER_79_702 ();
 FILLCELL_X4 FILLER_79_710 ();
 FILLCELL_X2 FILLER_79_714 ();
 FILLCELL_X8 FILLER_79_734 ();
 FILLCELL_X2 FILLER_79_742 ();
 FILLCELL_X2 FILLER_79_750 ();
 FILLCELL_X1 FILLER_79_752 ();
 FILLCELL_X4 FILLER_79_779 ();
 FILLCELL_X2 FILLER_79_783 ();
 FILLCELL_X1 FILLER_79_785 ();
 FILLCELL_X8 FILLER_79_788 ();
 FILLCELL_X2 FILLER_79_796 ();
 FILLCELL_X1 FILLER_79_798 ();
 FILLCELL_X4 FILLER_79_835 ();
 FILLCELL_X1 FILLER_79_839 ();
 FILLCELL_X16 FILLER_79_856 ();
 FILLCELL_X2 FILLER_79_872 ();
 FILLCELL_X1 FILLER_79_874 ();
 FILLCELL_X4 FILLER_79_880 ();
 FILLCELL_X2 FILLER_79_884 ();
 FILLCELL_X16 FILLER_79_891 ();
 FILLCELL_X4 FILLER_79_907 ();
 FILLCELL_X2 FILLER_79_911 ();
 FILLCELL_X1 FILLER_79_913 ();
 FILLCELL_X32 FILLER_79_948 ();
 FILLCELL_X2 FILLER_79_980 ();
 FILLCELL_X8 FILLER_80_1 ();
 FILLCELL_X2 FILLER_80_9 ();
 FILLCELL_X1 FILLER_80_11 ();
 FILLCELL_X8 FILLER_80_16 ();
 FILLCELL_X1 FILLER_80_24 ();
 FILLCELL_X4 FILLER_80_33 ();
 FILLCELL_X8 FILLER_80_41 ();
 FILLCELL_X4 FILLER_80_49 ();
 FILLCELL_X2 FILLER_80_53 ();
 FILLCELL_X1 FILLER_80_79 ();
 FILLCELL_X4 FILLER_80_85 ();
 FILLCELL_X1 FILLER_80_89 ();
 FILLCELL_X4 FILLER_80_113 ();
 FILLCELL_X2 FILLER_80_117 ();
 FILLCELL_X1 FILLER_80_119 ();
 FILLCELL_X1 FILLER_80_139 ();
 FILLCELL_X8 FILLER_80_154 ();
 FILLCELL_X1 FILLER_80_162 ();
 FILLCELL_X2 FILLER_80_166 ();
 FILLCELL_X8 FILLER_80_188 ();
 FILLCELL_X2 FILLER_80_196 ();
 FILLCELL_X1 FILLER_80_198 ();
 FILLCELL_X2 FILLER_80_238 ();
 FILLCELL_X1 FILLER_80_240 ();
 FILLCELL_X2 FILLER_80_258 ();
 FILLCELL_X16 FILLER_80_269 ();
 FILLCELL_X1 FILLER_80_285 ();
 FILLCELL_X8 FILLER_80_299 ();
 FILLCELL_X1 FILLER_80_307 ();
 FILLCELL_X4 FILLER_80_336 ();
 FILLCELL_X1 FILLER_80_340 ();
 FILLCELL_X2 FILLER_80_350 ();
 FILLCELL_X1 FILLER_80_352 ();
 FILLCELL_X1 FILLER_80_377 ();
 FILLCELL_X4 FILLER_80_394 ();
 FILLCELL_X2 FILLER_80_398 ();
 FILLCELL_X1 FILLER_80_414 ();
 FILLCELL_X8 FILLER_80_442 ();
 FILLCELL_X2 FILLER_80_450 ();
 FILLCELL_X1 FILLER_80_501 ();
 FILLCELL_X1 FILLER_80_512 ();
 FILLCELL_X4 FILLER_80_529 ();
 FILLCELL_X2 FILLER_80_533 ();
 FILLCELL_X1 FILLER_80_535 ();
 FILLCELL_X8 FILLER_80_552 ();
 FILLCELL_X1 FILLER_80_560 ();
 FILLCELL_X2 FILLER_80_584 ();
 FILLCELL_X4 FILLER_80_593 ();
 FILLCELL_X4 FILLER_80_606 ();
 FILLCELL_X1 FILLER_80_610 ();
 FILLCELL_X1 FILLER_80_630 ();
 FILLCELL_X4 FILLER_80_632 ();
 FILLCELL_X2 FILLER_80_636 ();
 FILLCELL_X1 FILLER_80_638 ();
 FILLCELL_X1 FILLER_80_658 ();
 FILLCELL_X2 FILLER_80_662 ();
 FILLCELL_X1 FILLER_80_664 ();
 FILLCELL_X8 FILLER_80_684 ();
 FILLCELL_X4 FILLER_80_692 ();
 FILLCELL_X2 FILLER_80_696 ();
 FILLCELL_X16 FILLER_80_715 ();
 FILLCELL_X4 FILLER_80_731 ();
 FILLCELL_X2 FILLER_80_735 ();
 FILLCELL_X1 FILLER_80_737 ();
 FILLCELL_X2 FILLER_80_748 ();
 FILLCELL_X1 FILLER_80_750 ();
 FILLCELL_X2 FILLER_80_760 ();
 FILLCELL_X8 FILLER_80_798 ();
 FILLCELL_X1 FILLER_80_806 ();
 FILLCELL_X1 FILLER_80_825 ();
 FILLCELL_X4 FILLER_80_829 ();
 FILLCELL_X2 FILLER_80_833 ();
 FILLCELL_X1 FILLER_80_835 ();
 FILLCELL_X2 FILLER_80_838 ();
 FILLCELL_X1 FILLER_80_840 ();
 FILLCELL_X4 FILLER_80_843 ();
 FILLCELL_X2 FILLER_80_847 ();
 FILLCELL_X1 FILLER_80_849 ();
 FILLCELL_X2 FILLER_80_852 ();
 FILLCELL_X1 FILLER_80_854 ();
 FILLCELL_X16 FILLER_80_868 ();
 FILLCELL_X8 FILLER_80_884 ();
 FILLCELL_X2 FILLER_80_892 ();
 FILLCELL_X1 FILLER_80_894 ();
 FILLCELL_X4 FILLER_80_898 ();
 FILLCELL_X1 FILLER_80_902 ();
 FILLCELL_X2 FILLER_80_913 ();
 FILLCELL_X1 FILLER_80_915 ();
 FILLCELL_X8 FILLER_80_926 ();
 FILLCELL_X2 FILLER_80_934 ();
 FILLCELL_X1 FILLER_80_936 ();
 FILLCELL_X32 FILLER_80_947 ();
 FILLCELL_X2 FILLER_80_979 ();
 FILLCELL_X1 FILLER_80_981 ();
 FILLCELL_X16 FILLER_81_1 ();
 FILLCELL_X4 FILLER_81_37 ();
 FILLCELL_X2 FILLER_81_41 ();
 FILLCELL_X1 FILLER_81_43 ();
 FILLCELL_X16 FILLER_81_48 ();
 FILLCELL_X8 FILLER_81_64 ();
 FILLCELL_X1 FILLER_81_72 ();
 FILLCELL_X2 FILLER_81_103 ();
 FILLCELL_X1 FILLER_81_135 ();
 FILLCELL_X1 FILLER_81_152 ();
 FILLCELL_X8 FILLER_81_169 ();
 FILLCELL_X2 FILLER_81_177 ();
 FILLCELL_X4 FILLER_81_182 ();
 FILLCELL_X2 FILLER_81_186 ();
 FILLCELL_X1 FILLER_81_188 ();
 FILLCELL_X4 FILLER_81_192 ();
 FILLCELL_X1 FILLER_81_203 ();
 FILLCELL_X4 FILLER_81_254 ();
 FILLCELL_X2 FILLER_81_263 ();
 FILLCELL_X1 FILLER_81_265 ();
 FILLCELL_X4 FILLER_81_270 ();
 FILLCELL_X16 FILLER_81_279 ();
 FILLCELL_X2 FILLER_81_295 ();
 FILLCELL_X2 FILLER_81_300 ();
 FILLCELL_X1 FILLER_81_302 ();
 FILLCELL_X1 FILLER_81_310 ();
 FILLCELL_X16 FILLER_81_330 ();
 FILLCELL_X2 FILLER_81_346 ();
 FILLCELL_X16 FILLER_81_355 ();
 FILLCELL_X4 FILLER_81_371 ();
 FILLCELL_X2 FILLER_81_375 ();
 FILLCELL_X8 FILLER_81_379 ();
 FILLCELL_X4 FILLER_81_387 ();
 FILLCELL_X1 FILLER_81_403 ();
 FILLCELL_X1 FILLER_81_442 ();
 FILLCELL_X1 FILLER_81_448 ();
 FILLCELL_X4 FILLER_81_452 ();
 FILLCELL_X16 FILLER_81_483 ();
 FILLCELL_X1 FILLER_81_499 ();
 FILLCELL_X8 FILLER_81_520 ();
 FILLCELL_X2 FILLER_81_528 ();
 FILLCELL_X1 FILLER_81_530 ();
 FILLCELL_X2 FILLER_81_540 ();
 FILLCELL_X8 FILLER_81_549 ();
 FILLCELL_X2 FILLER_81_557 ();
 FILLCELL_X1 FILLER_81_559 ();
 FILLCELL_X4 FILLER_81_570 ();
 FILLCELL_X4 FILLER_81_576 ();
 FILLCELL_X1 FILLER_81_580 ();
 FILLCELL_X2 FILLER_81_586 ();
 FILLCELL_X1 FILLER_81_588 ();
 FILLCELL_X16 FILLER_81_596 ();
 FILLCELL_X8 FILLER_81_612 ();
 FILLCELL_X8 FILLER_81_657 ();
 FILLCELL_X2 FILLER_81_665 ();
 FILLCELL_X16 FILLER_81_682 ();
 FILLCELL_X1 FILLER_81_698 ();
 FILLCELL_X2 FILLER_81_716 ();
 FILLCELL_X4 FILLER_81_723 ();
 FILLCELL_X1 FILLER_81_727 ();
 FILLCELL_X8 FILLER_81_730 ();
 FILLCELL_X4 FILLER_81_738 ();
 FILLCELL_X2 FILLER_81_742 ();
 FILLCELL_X1 FILLER_81_744 ();
 FILLCELL_X2 FILLER_81_751 ();
 FILLCELL_X1 FILLER_81_753 ();
 FILLCELL_X8 FILLER_81_757 ();
 FILLCELL_X8 FILLER_81_774 ();
 FILLCELL_X4 FILLER_81_782 ();
 FILLCELL_X2 FILLER_81_786 ();
 FILLCELL_X1 FILLER_81_788 ();
 FILLCELL_X8 FILLER_81_798 ();
 FILLCELL_X1 FILLER_81_806 ();
 FILLCELL_X4 FILLER_81_816 ();
 FILLCELL_X2 FILLER_81_820 ();
 FILLCELL_X1 FILLER_81_822 ();
 FILLCELL_X2 FILLER_81_839 ();
 FILLCELL_X16 FILLER_81_843 ();
 FILLCELL_X4 FILLER_81_859 ();
 FILLCELL_X1 FILLER_81_863 ();
 FILLCELL_X8 FILLER_81_873 ();
 FILLCELL_X4 FILLER_81_881 ();
 FILLCELL_X2 FILLER_81_885 ();
 FILLCELL_X1 FILLER_81_887 ();
 FILLCELL_X1 FILLER_81_894 ();
 FILLCELL_X8 FILLER_81_918 ();
 FILLCELL_X4 FILLER_81_926 ();
 FILLCELL_X2 FILLER_81_930 ();
 FILLCELL_X1 FILLER_81_932 ();
 FILLCELL_X16 FILLER_81_951 ();
 FILLCELL_X8 FILLER_81_967 ();
 FILLCELL_X4 FILLER_81_975 ();
 FILLCELL_X2 FILLER_81_979 ();
 FILLCELL_X1 FILLER_81_981 ();
 FILLCELL_X2 FILLER_82_1 ();
 FILLCELL_X2 FILLER_82_24 ();
 FILLCELL_X16 FILLER_82_50 ();
 FILLCELL_X8 FILLER_82_66 ();
 FILLCELL_X2 FILLER_82_74 ();
 FILLCELL_X2 FILLER_82_93 ();
 FILLCELL_X2 FILLER_82_108 ();
 FILLCELL_X8 FILLER_82_118 ();
 FILLCELL_X4 FILLER_82_126 ();
 FILLCELL_X2 FILLER_82_130 ();
 FILLCELL_X4 FILLER_82_136 ();
 FILLCELL_X2 FILLER_82_140 ();
 FILLCELL_X2 FILLER_82_145 ();
 FILLCELL_X8 FILLER_82_166 ();
 FILLCELL_X2 FILLER_82_174 ();
 FILLCELL_X4 FILLER_82_179 ();
 FILLCELL_X2 FILLER_82_183 ();
 FILLCELL_X1 FILLER_82_185 ();
 FILLCELL_X2 FILLER_82_189 ();
 FILLCELL_X8 FILLER_82_211 ();
 FILLCELL_X1 FILLER_82_222 ();
 FILLCELL_X4 FILLER_82_242 ();
 FILLCELL_X1 FILLER_82_246 ();
 FILLCELL_X8 FILLER_82_275 ();
 FILLCELL_X4 FILLER_82_283 ();
 FILLCELL_X2 FILLER_82_287 ();
 FILLCELL_X2 FILLER_82_297 ();
 FILLCELL_X1 FILLER_82_299 ();
 FILLCELL_X2 FILLER_82_314 ();
 FILLCELL_X1 FILLER_82_316 ();
 FILLCELL_X1 FILLER_82_323 ();
 FILLCELL_X2 FILLER_82_328 ();
 FILLCELL_X16 FILLER_82_379 ();
 FILLCELL_X4 FILLER_82_395 ();
 FILLCELL_X2 FILLER_82_437 ();
 FILLCELL_X4 FILLER_82_456 ();
 FILLCELL_X2 FILLER_82_460 ();
 FILLCELL_X1 FILLER_82_462 ();
 FILLCELL_X8 FILLER_82_480 ();
 FILLCELL_X1 FILLER_82_488 ();
 FILLCELL_X1 FILLER_82_520 ();
 FILLCELL_X2 FILLER_82_539 ();
 FILLCELL_X8 FILLER_82_548 ();
 FILLCELL_X2 FILLER_82_582 ();
 FILLCELL_X8 FILLER_82_589 ();
 FILLCELL_X2 FILLER_82_597 ();
 FILLCELL_X1 FILLER_82_599 ();
 FILLCELL_X8 FILLER_82_609 ();
 FILLCELL_X2 FILLER_82_628 ();
 FILLCELL_X1 FILLER_82_630 ();
 FILLCELL_X1 FILLER_82_643 ();
 FILLCELL_X1 FILLER_82_702 ();
 FILLCELL_X4 FILLER_82_711 ();
 FILLCELL_X8 FILLER_82_732 ();
 FILLCELL_X4 FILLER_82_740 ();
 FILLCELL_X1 FILLER_82_744 ();
 FILLCELL_X16 FILLER_82_774 ();
 FILLCELL_X1 FILLER_82_790 ();
 FILLCELL_X8 FILLER_82_797 ();
 FILLCELL_X2 FILLER_82_805 ();
 FILLCELL_X2 FILLER_82_813 ();
 FILLCELL_X1 FILLER_82_820 ();
 FILLCELL_X2 FILLER_82_824 ();
 FILLCELL_X4 FILLER_82_852 ();
 FILLCELL_X16 FILLER_82_861 ();
 FILLCELL_X8 FILLER_82_877 ();
 FILLCELL_X4 FILLER_82_885 ();
 FILLCELL_X2 FILLER_82_889 ();
 FILLCELL_X1 FILLER_82_891 ();
 FILLCELL_X32 FILLER_82_898 ();
 FILLCELL_X32 FILLER_82_930 ();
 FILLCELL_X16 FILLER_82_962 ();
 FILLCELL_X4 FILLER_82_978 ();
 FILLCELL_X4 FILLER_83_4 ();
 FILLCELL_X4 FILLER_83_14 ();
 FILLCELL_X2 FILLER_83_24 ();
 FILLCELL_X8 FILLER_83_31 ();
 FILLCELL_X32 FILLER_83_46 ();
 FILLCELL_X4 FILLER_83_83 ();
 FILLCELL_X2 FILLER_83_87 ();
 FILLCELL_X16 FILLER_83_131 ();
 FILLCELL_X1 FILLER_83_147 ();
 FILLCELL_X16 FILLER_83_157 ();
 FILLCELL_X2 FILLER_83_173 ();
 FILLCELL_X1 FILLER_83_175 ();
 FILLCELL_X16 FILLER_83_190 ();
 FILLCELL_X2 FILLER_83_213 ();
 FILLCELL_X1 FILLER_83_215 ();
 FILLCELL_X8 FILLER_83_234 ();
 FILLCELL_X1 FILLER_83_242 ();
 FILLCELL_X16 FILLER_83_256 ();
 FILLCELL_X4 FILLER_83_272 ();
 FILLCELL_X2 FILLER_83_276 ();
 FILLCELL_X1 FILLER_83_278 ();
 FILLCELL_X32 FILLER_83_305 ();
 FILLCELL_X8 FILLER_83_337 ();
 FILLCELL_X4 FILLER_83_345 ();
 FILLCELL_X1 FILLER_83_349 ();
 FILLCELL_X4 FILLER_83_359 ();
 FILLCELL_X2 FILLER_83_376 ();
 FILLCELL_X2 FILLER_83_385 ();
 FILLCELL_X1 FILLER_83_387 ();
 FILLCELL_X8 FILLER_83_481 ();
 FILLCELL_X4 FILLER_83_489 ();
 FILLCELL_X1 FILLER_83_493 ();
 FILLCELL_X2 FILLER_83_511 ();
 FILLCELL_X2 FILLER_83_530 ();
 FILLCELL_X1 FILLER_83_577 ();
 FILLCELL_X2 FILLER_83_597 ();
 FILLCELL_X2 FILLER_83_623 ();
 FILLCELL_X4 FILLER_83_674 ();
 FILLCELL_X1 FILLER_83_678 ();
 FILLCELL_X16 FILLER_83_703 ();
 FILLCELL_X4 FILLER_83_719 ();
 FILLCELL_X1 FILLER_83_723 ();
 FILLCELL_X4 FILLER_83_733 ();
 FILLCELL_X1 FILLER_83_737 ();
 FILLCELL_X8 FILLER_83_747 ();
 FILLCELL_X1 FILLER_83_755 ();
 FILLCELL_X2 FILLER_83_759 ();
 FILLCELL_X1 FILLER_83_761 ();
 FILLCELL_X8 FILLER_83_765 ();
 FILLCELL_X8 FILLER_83_775 ();
 FILLCELL_X4 FILLER_83_783 ();
 FILLCELL_X2 FILLER_83_787 ();
 FILLCELL_X8 FILLER_83_811 ();
 FILLCELL_X2 FILLER_83_819 ();
 FILLCELL_X16 FILLER_83_823 ();
 FILLCELL_X4 FILLER_83_839 ();
 FILLCELL_X1 FILLER_83_843 ();
 FILLCELL_X32 FILLER_83_849 ();
 FILLCELL_X32 FILLER_83_881 ();
 FILLCELL_X32 FILLER_83_913 ();
 FILLCELL_X32 FILLER_83_945 ();
 FILLCELL_X4 FILLER_83_977 ();
 FILLCELL_X1 FILLER_83_981 ();
 FILLCELL_X4 FILLER_84_1 ();
 FILLCELL_X32 FILLER_84_29 ();
 FILLCELL_X8 FILLER_84_61 ();
 FILLCELL_X1 FILLER_84_112 ();
 FILLCELL_X4 FILLER_84_124 ();
 FILLCELL_X4 FILLER_84_139 ();
 FILLCELL_X1 FILLER_84_143 ();
 FILLCELL_X8 FILLER_84_163 ();
 FILLCELL_X4 FILLER_84_171 ();
 FILLCELL_X1 FILLER_84_175 ();
 FILLCELL_X16 FILLER_84_192 ();
 FILLCELL_X8 FILLER_84_208 ();
 FILLCELL_X4 FILLER_84_216 ();
 FILLCELL_X2 FILLER_84_220 ();
 FILLCELL_X1 FILLER_84_222 ();
 FILLCELL_X16 FILLER_84_232 ();
 FILLCELL_X2 FILLER_84_248 ();
 FILLCELL_X1 FILLER_84_250 ();
 FILLCELL_X16 FILLER_84_270 ();
 FILLCELL_X1 FILLER_84_286 ();
 FILLCELL_X4 FILLER_84_292 ();
 FILLCELL_X2 FILLER_84_296 ();
 FILLCELL_X32 FILLER_84_303 ();
 FILLCELL_X16 FILLER_84_335 ();
 FILLCELL_X2 FILLER_84_351 ();
 FILLCELL_X8 FILLER_84_380 ();
 FILLCELL_X4 FILLER_84_388 ();
 FILLCELL_X2 FILLER_84_392 ();
 FILLCELL_X1 FILLER_84_394 ();
 FILLCELL_X4 FILLER_84_420 ();
 FILLCELL_X4 FILLER_84_429 ();
 FILLCELL_X1 FILLER_84_446 ();
 FILLCELL_X8 FILLER_84_454 ();
 FILLCELL_X1 FILLER_84_462 ();
 FILLCELL_X4 FILLER_84_470 ();
 FILLCELL_X2 FILLER_84_474 ();
 FILLCELL_X8 FILLER_84_487 ();
 FILLCELL_X4 FILLER_84_495 ();
 FILLCELL_X2 FILLER_84_499 ();
 FILLCELL_X4 FILLER_84_507 ();
 FILLCELL_X2 FILLER_84_511 ();
 FILLCELL_X1 FILLER_84_513 ();
 FILLCELL_X8 FILLER_84_539 ();
 FILLCELL_X4 FILLER_84_547 ();
 FILLCELL_X1 FILLER_84_551 ();
 FILLCELL_X4 FILLER_84_569 ();
 FILLCELL_X2 FILLER_84_573 ();
 FILLCELL_X1 FILLER_84_575 ();
 FILLCELL_X8 FILLER_84_595 ();
 FILLCELL_X2 FILLER_84_603 ();
 FILLCELL_X4 FILLER_84_624 ();
 FILLCELL_X2 FILLER_84_628 ();
 FILLCELL_X1 FILLER_84_630 ();
 FILLCELL_X4 FILLER_84_632 ();
 FILLCELL_X1 FILLER_84_655 ();
 FILLCELL_X1 FILLER_84_675 ();
 FILLCELL_X8 FILLER_84_687 ();
 FILLCELL_X2 FILLER_84_695 ();
 FILLCELL_X1 FILLER_84_697 ();
 FILLCELL_X16 FILLER_84_700 ();
 FILLCELL_X8 FILLER_84_716 ();
 FILLCELL_X2 FILLER_84_724 ();
 FILLCELL_X1 FILLER_84_726 ();
 FILLCELL_X2 FILLER_84_737 ();
 FILLCELL_X16 FILLER_84_765 ();
 FILLCELL_X1 FILLER_84_781 ();
 FILLCELL_X1 FILLER_84_800 ();
 FILLCELL_X1 FILLER_84_803 ();
 FILLCELL_X1 FILLER_84_809 ();
 FILLCELL_X2 FILLER_84_826 ();
 FILLCELL_X32 FILLER_84_830 ();
 FILLCELL_X32 FILLER_84_862 ();
 FILLCELL_X32 FILLER_84_894 ();
 FILLCELL_X32 FILLER_84_926 ();
 FILLCELL_X16 FILLER_84_958 ();
 FILLCELL_X8 FILLER_84_974 ();
 FILLCELL_X2 FILLER_85_4 ();
 FILLCELL_X2 FILLER_85_30 ();
 FILLCELL_X8 FILLER_85_52 ();
 FILLCELL_X4 FILLER_85_60 ();
 FILLCELL_X2 FILLER_85_64 ();
 FILLCELL_X1 FILLER_85_66 ();
 FILLCELL_X1 FILLER_85_89 ();
 FILLCELL_X8 FILLER_85_93 ();
 FILLCELL_X4 FILLER_85_101 ();
 FILLCELL_X2 FILLER_85_105 ();
 FILLCELL_X8 FILLER_85_145 ();
 FILLCELL_X1 FILLER_85_153 ();
 FILLCELL_X4 FILLER_85_170 ();
 FILLCELL_X2 FILLER_85_174 ();
 FILLCELL_X1 FILLER_85_176 ();
 FILLCELL_X4 FILLER_85_194 ();
 FILLCELL_X2 FILLER_85_198 ();
 FILLCELL_X2 FILLER_85_209 ();
 FILLCELL_X1 FILLER_85_211 ();
 FILLCELL_X2 FILLER_85_218 ();
 FILLCELL_X1 FILLER_85_220 ();
 FILLCELL_X2 FILLER_85_238 ();
 FILLCELL_X1 FILLER_85_240 ();
 FILLCELL_X8 FILLER_85_264 ();
 FILLCELL_X4 FILLER_85_272 ();
 FILLCELL_X8 FILLER_85_280 ();
 FILLCELL_X8 FILLER_85_293 ();
 FILLCELL_X4 FILLER_85_301 ();
 FILLCELL_X2 FILLER_85_305 ();
 FILLCELL_X1 FILLER_85_307 ();
 FILLCELL_X1 FILLER_85_321 ();
 FILLCELL_X4 FILLER_85_348 ();
 FILLCELL_X2 FILLER_85_352 ();
 FILLCELL_X1 FILLER_85_354 ();
 FILLCELL_X2 FILLER_85_362 ();
 FILLCELL_X1 FILLER_85_364 ();
 FILLCELL_X2 FILLER_85_367 ();
 FILLCELL_X1 FILLER_85_382 ();
 FILLCELL_X2 FILLER_85_392 ();
 FILLCELL_X1 FILLER_85_394 ();
 FILLCELL_X8 FILLER_85_400 ();
 FILLCELL_X4 FILLER_85_408 ();
 FILLCELL_X2 FILLER_85_412 ();
 FILLCELL_X1 FILLER_85_414 ();
 FILLCELL_X4 FILLER_85_449 ();
 FILLCELL_X1 FILLER_85_453 ();
 FILLCELL_X2 FILLER_85_472 ();
 FILLCELL_X1 FILLER_85_474 ();
 FILLCELL_X8 FILLER_85_521 ();
 FILLCELL_X2 FILLER_85_535 ();
 FILLCELL_X8 FILLER_85_542 ();
 FILLCELL_X4 FILLER_85_550 ();
 FILLCELL_X32 FILLER_85_582 ();
 FILLCELL_X4 FILLER_85_614 ();
 FILLCELL_X1 FILLER_85_618 ();
 FILLCELL_X2 FILLER_85_630 ();
 FILLCELL_X1 FILLER_85_632 ();
 FILLCELL_X4 FILLER_85_658 ();
 FILLCELL_X2 FILLER_85_693 ();
 FILLCELL_X1 FILLER_85_695 ();
 FILLCELL_X8 FILLER_85_702 ();
 FILLCELL_X4 FILLER_85_710 ();
 FILLCELL_X2 FILLER_85_714 ();
 FILLCELL_X1 FILLER_85_716 ();
 FILLCELL_X1 FILLER_85_734 ();
 FILLCELL_X4 FILLER_85_750 ();
 FILLCELL_X2 FILLER_85_754 ();
 FILLCELL_X4 FILLER_85_759 ();
 FILLCELL_X2 FILLER_85_763 ();
 FILLCELL_X8 FILLER_85_797 ();
 FILLCELL_X1 FILLER_85_829 ();
 FILLCELL_X32 FILLER_85_835 ();
 FILLCELL_X32 FILLER_85_867 ();
 FILLCELL_X32 FILLER_85_899 ();
 FILLCELL_X32 FILLER_85_931 ();
 FILLCELL_X16 FILLER_85_963 ();
 FILLCELL_X2 FILLER_85_979 ();
 FILLCELL_X1 FILLER_85_981 ();
 FILLCELL_X2 FILLER_86_1 ();
 FILLCELL_X1 FILLER_86_3 ();
 FILLCELL_X2 FILLER_86_7 ();
 FILLCELL_X8 FILLER_86_12 ();
 FILLCELL_X1 FILLER_86_20 ();
 FILLCELL_X8 FILLER_86_24 ();
 FILLCELL_X2 FILLER_86_32 ();
 FILLCELL_X32 FILLER_86_54 ();
 FILLCELL_X32 FILLER_86_86 ();
 FILLCELL_X16 FILLER_86_118 ();
 FILLCELL_X1 FILLER_86_134 ();
 FILLCELL_X4 FILLER_86_152 ();
 FILLCELL_X1 FILLER_86_156 ();
 FILLCELL_X16 FILLER_86_176 ();
 FILLCELL_X4 FILLER_86_192 ();
 FILLCELL_X2 FILLER_86_196 ();
 FILLCELL_X4 FILLER_86_217 ();
 FILLCELL_X2 FILLER_86_221 ();
 FILLCELL_X4 FILLER_86_232 ();
 FILLCELL_X4 FILLER_86_268 ();
 FILLCELL_X1 FILLER_86_272 ();
 FILLCELL_X8 FILLER_86_290 ();
 FILLCELL_X1 FILLER_86_298 ();
 FILLCELL_X4 FILLER_86_304 ();
 FILLCELL_X1 FILLER_86_308 ();
 FILLCELL_X1 FILLER_86_320 ();
 FILLCELL_X1 FILLER_86_324 ();
 FILLCELL_X32 FILLER_86_328 ();
 FILLCELL_X4 FILLER_86_360 ();
 FILLCELL_X2 FILLER_86_364 ();
 FILLCELL_X2 FILLER_86_380 ();
 FILLCELL_X1 FILLER_86_382 ();
 FILLCELL_X1 FILLER_86_386 ();
 FILLCELL_X2 FILLER_86_390 ();
 FILLCELL_X2 FILLER_86_418 ();
 FILLCELL_X8 FILLER_86_472 ();
 FILLCELL_X2 FILLER_86_489 ();
 FILLCELL_X1 FILLER_86_491 ();
 FILLCELL_X8 FILLER_86_502 ();
 FILLCELL_X4 FILLER_86_510 ();
 FILLCELL_X1 FILLER_86_514 ();
 FILLCELL_X4 FILLER_86_518 ();
 FILLCELL_X1 FILLER_86_522 ();
 FILLCELL_X4 FILLER_86_542 ();
 FILLCELL_X4 FILLER_86_549 ();
 FILLCELL_X1 FILLER_86_553 ();
 FILLCELL_X4 FILLER_86_567 ();
 FILLCELL_X32 FILLER_86_580 ();
 FILLCELL_X4 FILLER_86_650 ();
 FILLCELL_X2 FILLER_86_654 ();
 FILLCELL_X8 FILLER_86_673 ();
 FILLCELL_X1 FILLER_86_681 ();
 FILLCELL_X8 FILLER_86_685 ();
 FILLCELL_X2 FILLER_86_693 ();
 FILLCELL_X1 FILLER_86_714 ();
 FILLCELL_X1 FILLER_86_724 ();
 FILLCELL_X2 FILLER_86_731 ();
 FILLCELL_X1 FILLER_86_743 ();
 FILLCELL_X16 FILLER_86_770 ();
 FILLCELL_X4 FILLER_86_789 ();
 FILLCELL_X1 FILLER_86_793 ();
 FILLCELL_X1 FILLER_86_804 ();
 FILLCELL_X4 FILLER_86_814 ();
 FILLCELL_X1 FILLER_86_818 ();
 FILLCELL_X8 FILLER_86_822 ();
 FILLCELL_X4 FILLER_86_830 ();
 FILLCELL_X2 FILLER_86_834 ();
 FILLCELL_X1 FILLER_86_836 ();
 FILLCELL_X2 FILLER_86_846 ();
 FILLCELL_X1 FILLER_86_860 ();
 FILLCELL_X8 FILLER_86_871 ();
 FILLCELL_X2 FILLER_86_879 ();
 FILLCELL_X16 FILLER_86_899 ();
 FILLCELL_X32 FILLER_86_938 ();
 FILLCELL_X8 FILLER_86_970 ();
 FILLCELL_X4 FILLER_86_978 ();
 FILLCELL_X2 FILLER_87_1 ();
 FILLCELL_X1 FILLER_87_3 ();
 FILLCELL_X1 FILLER_87_21 ();
 FILLCELL_X8 FILLER_87_26 ();
 FILLCELL_X2 FILLER_87_34 ();
 FILLCELL_X1 FILLER_87_36 ();
 FILLCELL_X8 FILLER_87_41 ();
 FILLCELL_X4 FILLER_87_49 ();
 FILLCELL_X1 FILLER_87_53 ();
 FILLCELL_X16 FILLER_87_67 ();
 FILLCELL_X8 FILLER_87_83 ();
 FILLCELL_X4 FILLER_87_91 ();
 FILLCELL_X2 FILLER_87_95 ();
 FILLCELL_X16 FILLER_87_108 ();
 FILLCELL_X8 FILLER_87_124 ();
 FILLCELL_X4 FILLER_87_132 ();
 FILLCELL_X16 FILLER_87_155 ();
 FILLCELL_X8 FILLER_87_171 ();
 FILLCELL_X1 FILLER_87_179 ();
 FILLCELL_X8 FILLER_87_198 ();
 FILLCELL_X4 FILLER_87_206 ();
 FILLCELL_X2 FILLER_87_210 ();
 FILLCELL_X1 FILLER_87_212 ();
 FILLCELL_X8 FILLER_87_216 ();
 FILLCELL_X2 FILLER_87_224 ();
 FILLCELL_X1 FILLER_87_229 ();
 FILLCELL_X8 FILLER_87_249 ();
 FILLCELL_X32 FILLER_87_260 ();
 FILLCELL_X1 FILLER_87_292 ();
 FILLCELL_X2 FILLER_87_312 ();
 FILLCELL_X1 FILLER_87_314 ();
 FILLCELL_X16 FILLER_87_330 ();
 FILLCELL_X4 FILLER_87_346 ();
 FILLCELL_X2 FILLER_87_350 ();
 FILLCELL_X4 FILLER_87_359 ();
 FILLCELL_X1 FILLER_87_363 ();
 FILLCELL_X1 FILLER_87_383 ();
 FILLCELL_X8 FILLER_87_395 ();
 FILLCELL_X4 FILLER_87_403 ();
 FILLCELL_X8 FILLER_87_429 ();
 FILLCELL_X2 FILLER_87_437 ();
 FILLCELL_X1 FILLER_87_439 ();
 FILLCELL_X2 FILLER_87_456 ();
 FILLCELL_X2 FILLER_87_467 ();
 FILLCELL_X1 FILLER_87_469 ();
 FILLCELL_X4 FILLER_87_490 ();
 FILLCELL_X2 FILLER_87_494 ();
 FILLCELL_X1 FILLER_87_496 ();
 FILLCELL_X2 FILLER_87_504 ();
 FILLCELL_X1 FILLER_87_513 ();
 FILLCELL_X8 FILLER_87_521 ();
 FILLCELL_X4 FILLER_87_529 ();
 FILLCELL_X4 FILLER_87_550 ();
 FILLCELL_X1 FILLER_87_554 ();
 FILLCELL_X4 FILLER_87_565 ();
 FILLCELL_X8 FILLER_87_603 ();
 FILLCELL_X1 FILLER_87_611 ();
 FILLCELL_X1 FILLER_87_623 ();
 FILLCELL_X32 FILLER_87_665 ();
 FILLCELL_X1 FILLER_87_697 ();
 FILLCELL_X8 FILLER_87_700 ();
 FILLCELL_X2 FILLER_87_708 ();
 FILLCELL_X1 FILLER_87_713 ();
 FILLCELL_X1 FILLER_87_717 ();
 FILLCELL_X2 FILLER_87_727 ();
 FILLCELL_X1 FILLER_87_741 ();
 FILLCELL_X8 FILLER_87_745 ();
 FILLCELL_X2 FILLER_87_753 ();
 FILLCELL_X8 FILLER_87_773 ();
 FILLCELL_X4 FILLER_87_781 ();
 FILLCELL_X4 FILLER_87_790 ();
 FILLCELL_X2 FILLER_87_794 ();
 FILLCELL_X1 FILLER_87_796 ();
 FILLCELL_X8 FILLER_87_806 ();
 FILLCELL_X4 FILLER_87_814 ();
 FILLCELL_X2 FILLER_87_818 ();
 FILLCELL_X1 FILLER_87_820 ();
 FILLCELL_X16 FILLER_87_823 ();
 FILLCELL_X4 FILLER_87_839 ();
 FILLCELL_X2 FILLER_87_843 ();
 FILLCELL_X1 FILLER_87_845 ();
 FILLCELL_X4 FILLER_87_878 ();
 FILLCELL_X4 FILLER_87_916 ();
 FILLCELL_X32 FILLER_87_936 ();
 FILLCELL_X8 FILLER_87_968 ();
 FILLCELL_X4 FILLER_87_976 ();
 FILLCELL_X2 FILLER_87_980 ();
 FILLCELL_X4 FILLER_88_1 ();
 FILLCELL_X16 FILLER_88_8 ();
 FILLCELL_X8 FILLER_88_24 ();
 FILLCELL_X2 FILLER_88_52 ();
 FILLCELL_X16 FILLER_88_67 ();
 FILLCELL_X2 FILLER_88_83 ();
 FILLCELL_X1 FILLER_88_85 ();
 FILLCELL_X32 FILLER_88_118 ();
 FILLCELL_X16 FILLER_88_150 ();
 FILLCELL_X4 FILLER_88_207 ();
 FILLCELL_X16 FILLER_88_228 ();
 FILLCELL_X8 FILLER_88_244 ();
 FILLCELL_X1 FILLER_88_270 ();
 FILLCELL_X1 FILLER_88_289 ();
 FILLCELL_X1 FILLER_88_295 ();
 FILLCELL_X1 FILLER_88_314 ();
 FILLCELL_X8 FILLER_88_332 ();
 FILLCELL_X4 FILLER_88_340 ();
 FILLCELL_X2 FILLER_88_344 ();
 FILLCELL_X4 FILLER_88_377 ();
 FILLCELL_X2 FILLER_88_381 ();
 FILLCELL_X8 FILLER_88_397 ();
 FILLCELL_X1 FILLER_88_405 ();
 FILLCELL_X4 FILLER_88_425 ();
 FILLCELL_X1 FILLER_88_444 ();
 FILLCELL_X1 FILLER_88_484 ();
 FILLCELL_X4 FILLER_88_498 ();
 FILLCELL_X4 FILLER_88_531 ();
 FILLCELL_X1 FILLER_88_535 ();
 FILLCELL_X2 FILLER_88_542 ();
 FILLCELL_X1 FILLER_88_544 ();
 FILLCELL_X4 FILLER_88_554 ();
 FILLCELL_X1 FILLER_88_558 ();
 FILLCELL_X4 FILLER_88_566 ();
 FILLCELL_X1 FILLER_88_570 ();
 FILLCELL_X1 FILLER_88_577 ();
 FILLCELL_X1 FILLER_88_600 ();
 FILLCELL_X4 FILLER_88_650 ();
 FILLCELL_X1 FILLER_88_654 ();
 FILLCELL_X4 FILLER_88_664 ();
 FILLCELL_X1 FILLER_88_668 ();
 FILLCELL_X16 FILLER_88_678 ();
 FILLCELL_X2 FILLER_88_717 ();
 FILLCELL_X8 FILLER_88_722 ();
 FILLCELL_X2 FILLER_88_730 ();
 FILLCELL_X1 FILLER_88_732 ();
 FILLCELL_X2 FILLER_88_736 ();
 FILLCELL_X4 FILLER_88_756 ();
 FILLCELL_X2 FILLER_88_760 ();
 FILLCELL_X1 FILLER_88_762 ();
 FILLCELL_X8 FILLER_88_781 ();
 FILLCELL_X4 FILLER_88_789 ();
 FILLCELL_X8 FILLER_88_800 ();
 FILLCELL_X1 FILLER_88_808 ();
 FILLCELL_X4 FILLER_88_828 ();
 FILLCELL_X1 FILLER_88_859 ();
 FILLCELL_X4 FILLER_88_862 ();
 FILLCELL_X2 FILLER_88_866 ();
 FILLCELL_X16 FILLER_88_870 ();
 FILLCELL_X2 FILLER_88_886 ();
 FILLCELL_X1 FILLER_88_888 ();
 FILLCELL_X8 FILLER_88_905 ();
 FILLCELL_X4 FILLER_88_913 ();
 FILLCELL_X1 FILLER_88_917 ();
 FILLCELL_X4 FILLER_88_920 ();
 FILLCELL_X2 FILLER_88_924 ();
 FILLCELL_X4 FILLER_88_930 ();
 FILLCELL_X1 FILLER_88_934 ();
 FILLCELL_X16 FILLER_88_955 ();
 FILLCELL_X8 FILLER_88_971 ();
 FILLCELL_X2 FILLER_88_979 ();
 FILLCELL_X1 FILLER_88_981 ();
 FILLCELL_X1 FILLER_89_24 ();
 FILLCELL_X4 FILLER_89_32 ();
 FILLCELL_X1 FILLER_89_36 ();
 FILLCELL_X8 FILLER_89_45 ();
 FILLCELL_X4 FILLER_89_53 ();
 FILLCELL_X2 FILLER_89_57 ();
 FILLCELL_X8 FILLER_89_65 ();
 FILLCELL_X4 FILLER_89_73 ();
 FILLCELL_X1 FILLER_89_77 ();
 FILLCELL_X4 FILLER_89_112 ();
 FILLCELL_X2 FILLER_89_116 ();
 FILLCELL_X16 FILLER_89_129 ();
 FILLCELL_X1 FILLER_89_145 ();
 FILLCELL_X8 FILLER_89_155 ();
 FILLCELL_X1 FILLER_89_163 ();
 FILLCELL_X32 FILLER_89_170 ();
 FILLCELL_X8 FILLER_89_202 ();
 FILLCELL_X16 FILLER_89_229 ();
 FILLCELL_X1 FILLER_89_245 ();
 FILLCELL_X1 FILLER_89_260 ();
 FILLCELL_X16 FILLER_89_330 ();
 FILLCELL_X4 FILLER_89_346 ();
 FILLCELL_X1 FILLER_89_350 ();
 FILLCELL_X4 FILLER_89_369 ();
 FILLCELL_X1 FILLER_89_373 ();
 FILLCELL_X1 FILLER_89_400 ();
 FILLCELL_X8 FILLER_89_403 ();
 FILLCELL_X8 FILLER_89_421 ();
 FILLCELL_X4 FILLER_89_429 ();
 FILLCELL_X2 FILLER_89_433 ();
 FILLCELL_X16 FILLER_89_454 ();
 FILLCELL_X4 FILLER_89_470 ();
 FILLCELL_X1 FILLER_89_474 ();
 FILLCELL_X1 FILLER_89_501 ();
 FILLCELL_X2 FILLER_89_543 ();
 FILLCELL_X1 FILLER_89_545 ();
 FILLCELL_X4 FILLER_89_565 ();
 FILLCELL_X2 FILLER_89_569 ();
 FILLCELL_X1 FILLER_89_571 ();
 FILLCELL_X4 FILLER_89_575 ();
 FILLCELL_X2 FILLER_89_579 ();
 FILLCELL_X1 FILLER_89_581 ();
 FILLCELL_X8 FILLER_89_601 ();
 FILLCELL_X4 FILLER_89_609 ();
 FILLCELL_X2 FILLER_89_613 ();
 FILLCELL_X1 FILLER_89_615 ();
 FILLCELL_X4 FILLER_89_652 ();
 FILLCELL_X1 FILLER_89_656 ();
 FILLCELL_X16 FILLER_89_694 ();
 FILLCELL_X2 FILLER_89_710 ();
 FILLCELL_X1 FILLER_89_712 ();
 FILLCELL_X8 FILLER_89_719 ();
 FILLCELL_X4 FILLER_89_727 ();
 FILLCELL_X1 FILLER_89_731 ();
 FILLCELL_X4 FILLER_89_735 ();
 FILLCELL_X4 FILLER_89_747 ();
 FILLCELL_X2 FILLER_89_760 ();
 FILLCELL_X8 FILLER_89_784 ();
 FILLCELL_X4 FILLER_89_792 ();
 FILLCELL_X1 FILLER_89_796 ();
 FILLCELL_X32 FILLER_89_802 ();
 FILLCELL_X4 FILLER_89_834 ();
 FILLCELL_X1 FILLER_89_838 ();
 FILLCELL_X4 FILLER_89_841 ();
 FILLCELL_X1 FILLER_89_845 ();
 FILLCELL_X2 FILLER_89_848 ();
 FILLCELL_X8 FILLER_89_866 ();
 FILLCELL_X4 FILLER_89_874 ();
 FILLCELL_X1 FILLER_89_878 ();
 FILLCELL_X16 FILLER_89_881 ();
 FILLCELL_X2 FILLER_89_897 ();
 FILLCELL_X1 FILLER_89_901 ();
 FILLCELL_X8 FILLER_89_904 ();
 FILLCELL_X2 FILLER_89_912 ();
 FILLCELL_X2 FILLER_89_916 ();
 FILLCELL_X32 FILLER_89_936 ();
 FILLCELL_X8 FILLER_89_968 ();
 FILLCELL_X4 FILLER_89_976 ();
 FILLCELL_X2 FILLER_89_980 ();
 FILLCELL_X1 FILLER_90_28 ();
 FILLCELL_X4 FILLER_90_32 ();
 FILLCELL_X1 FILLER_90_39 ();
 FILLCELL_X16 FILLER_90_63 ();
 FILLCELL_X4 FILLER_90_79 ();
 FILLCELL_X1 FILLER_90_83 ();
 FILLCELL_X2 FILLER_90_112 ();
 FILLCELL_X1 FILLER_90_114 ();
 FILLCELL_X8 FILLER_90_134 ();
 FILLCELL_X2 FILLER_90_142 ();
 FILLCELL_X1 FILLER_90_144 ();
 FILLCELL_X4 FILLER_90_179 ();
 FILLCELL_X1 FILLER_90_183 ();
 FILLCELL_X32 FILLER_90_201 ();
 FILLCELL_X4 FILLER_90_233 ();
 FILLCELL_X1 FILLER_90_237 ();
 FILLCELL_X4 FILLER_90_257 ();
 FILLCELL_X2 FILLER_90_261 ();
 FILLCELL_X8 FILLER_90_289 ();
 FILLCELL_X1 FILLER_90_297 ();
 FILLCELL_X2 FILLER_90_322 ();
 FILLCELL_X4 FILLER_90_343 ();
 FILLCELL_X1 FILLER_90_347 ();
 FILLCELL_X8 FILLER_90_357 ();
 FILLCELL_X2 FILLER_90_365 ();
 FILLCELL_X1 FILLER_90_367 ();
 FILLCELL_X8 FILLER_90_377 ();
 FILLCELL_X8 FILLER_90_394 ();
 FILLCELL_X4 FILLER_90_402 ();
 FILLCELL_X2 FILLER_90_406 ();
 FILLCELL_X1 FILLER_90_408 ();
 FILLCELL_X8 FILLER_90_428 ();
 FILLCELL_X2 FILLER_90_436 ();
 FILLCELL_X32 FILLER_90_462 ();
 FILLCELL_X16 FILLER_90_494 ();
 FILLCELL_X8 FILLER_90_510 ();
 FILLCELL_X4 FILLER_90_518 ();
 FILLCELL_X2 FILLER_90_522 ();
 FILLCELL_X2 FILLER_90_531 ();
 FILLCELL_X32 FILLER_90_552 ();
 FILLCELL_X16 FILLER_90_584 ();
 FILLCELL_X8 FILLER_90_600 ();
 FILLCELL_X8 FILLER_90_616 ();
 FILLCELL_X4 FILLER_90_624 ();
 FILLCELL_X2 FILLER_90_628 ();
 FILLCELL_X1 FILLER_90_630 ();
 FILLCELL_X4 FILLER_90_666 ();
 FILLCELL_X2 FILLER_90_670 ();
 FILLCELL_X1 FILLER_90_672 ();
 FILLCELL_X4 FILLER_90_699 ();
 FILLCELL_X2 FILLER_90_720 ();
 FILLCELL_X1 FILLER_90_729 ();
 FILLCELL_X4 FILLER_90_736 ();
 FILLCELL_X2 FILLER_90_740 ();
 FILLCELL_X1 FILLER_90_769 ();
 FILLCELL_X1 FILLER_90_779 ();
 FILLCELL_X2 FILLER_90_783 ();
 FILLCELL_X1 FILLER_90_785 ();
 FILLCELL_X4 FILLER_90_807 ();
 FILLCELL_X2 FILLER_90_811 ();
 FILLCELL_X1 FILLER_90_813 ();
 FILLCELL_X1 FILLER_90_830 ();
 FILLCELL_X4 FILLER_90_833 ();
 FILLCELL_X1 FILLER_90_849 ();
 FILLCELL_X16 FILLER_90_852 ();
 FILLCELL_X2 FILLER_90_868 ();
 FILLCELL_X1 FILLER_90_870 ();
 FILLCELL_X4 FILLER_90_877 ();
 FILLCELL_X1 FILLER_90_881 ();
 FILLCELL_X4 FILLER_90_888 ();
 FILLCELL_X2 FILLER_90_892 ();
 FILLCELL_X8 FILLER_90_910 ();
 FILLCELL_X1 FILLER_90_918 ();
 FILLCELL_X2 FILLER_90_929 ();
 FILLCELL_X1 FILLER_90_933 ();
 FILLCELL_X2 FILLER_90_944 ();
 FILLCELL_X32 FILLER_90_948 ();
 FILLCELL_X2 FILLER_90_980 ();
 FILLCELL_X16 FILLER_91_1 ();
 FILLCELL_X2 FILLER_91_17 ();
 FILLCELL_X2 FILLER_91_36 ();
 FILLCELL_X1 FILLER_91_42 ();
 FILLCELL_X1 FILLER_91_47 ();
 FILLCELL_X16 FILLER_91_51 ();
 FILLCELL_X4 FILLER_91_67 ();
 FILLCELL_X1 FILLER_91_71 ();
 FILLCELL_X8 FILLER_91_114 ();
 FILLCELL_X2 FILLER_91_122 ();
 FILLCELL_X8 FILLER_91_131 ();
 FILLCELL_X2 FILLER_91_139 ();
 FILLCELL_X1 FILLER_91_141 ();
 FILLCELL_X16 FILLER_91_163 ();
 FILLCELL_X4 FILLER_91_179 ();
 FILLCELL_X32 FILLER_91_200 ();
 FILLCELL_X8 FILLER_91_232 ();
 FILLCELL_X4 FILLER_91_240 ();
 FILLCELL_X1 FILLER_91_244 ();
 FILLCELL_X8 FILLER_91_252 ();
 FILLCELL_X2 FILLER_91_260 ();
 FILLCELL_X4 FILLER_91_269 ();
 FILLCELL_X2 FILLER_91_273 ();
 FILLCELL_X4 FILLER_91_286 ();
 FILLCELL_X1 FILLER_91_295 ();
 FILLCELL_X2 FILLER_91_307 ();
 FILLCELL_X16 FILLER_91_319 ();
 FILLCELL_X4 FILLER_91_335 ();
 FILLCELL_X2 FILLER_91_339 ();
 FILLCELL_X8 FILLER_91_357 ();
 FILLCELL_X4 FILLER_91_365 ();
 FILLCELL_X2 FILLER_91_387 ();
 FILLCELL_X2 FILLER_91_405 ();
 FILLCELL_X1 FILLER_91_458 ();
 FILLCELL_X8 FILLER_91_478 ();
 FILLCELL_X4 FILLER_91_486 ();
 FILLCELL_X1 FILLER_91_490 ();
 FILLCELL_X16 FILLER_91_497 ();
 FILLCELL_X8 FILLER_91_513 ();
 FILLCELL_X2 FILLER_91_521 ();
 FILLCELL_X1 FILLER_91_523 ();
 FILLCELL_X16 FILLER_91_535 ();
 FILLCELL_X4 FILLER_91_551 ();
 FILLCELL_X1 FILLER_91_555 ();
 FILLCELL_X4 FILLER_91_575 ();
 FILLCELL_X2 FILLER_91_584 ();
 FILLCELL_X1 FILLER_91_586 ();
 FILLCELL_X1 FILLER_91_600 ();
 FILLCELL_X1 FILLER_91_606 ();
 FILLCELL_X4 FILLER_91_627 ();
 FILLCELL_X2 FILLER_91_631 ();
 FILLCELL_X8 FILLER_91_691 ();
 FILLCELL_X2 FILLER_91_699 ();
 FILLCELL_X8 FILLER_91_718 ();
 FILLCELL_X1 FILLER_91_726 ();
 FILLCELL_X2 FILLER_91_733 ();
 FILLCELL_X16 FILLER_91_741 ();
 FILLCELL_X4 FILLER_91_757 ();
 FILLCELL_X4 FILLER_91_767 ();
 FILLCELL_X2 FILLER_91_771 ();
 FILLCELL_X2 FILLER_91_810 ();
 FILLCELL_X2 FILLER_91_824 ();
 FILLCELL_X1 FILLER_91_826 ();
 FILLCELL_X2 FILLER_91_845 ();
 FILLCELL_X1 FILLER_91_847 ();
 FILLCELL_X4 FILLER_91_864 ();
 FILLCELL_X1 FILLER_91_868 ();
 FILLCELL_X8 FILLER_91_891 ();
 FILLCELL_X2 FILLER_91_899 ();
 FILLCELL_X4 FILLER_91_937 ();
 FILLCELL_X2 FILLER_91_944 ();
 FILLCELL_X1 FILLER_91_946 ();
 FILLCELL_X16 FILLER_91_957 ();
 FILLCELL_X8 FILLER_91_973 ();
 FILLCELL_X1 FILLER_91_981 ();
 FILLCELL_X4 FILLER_92_1 ();
 FILLCELL_X16 FILLER_92_22 ();
 FILLCELL_X8 FILLER_92_38 ();
 FILLCELL_X1 FILLER_92_46 ();
 FILLCELL_X8 FILLER_92_52 ();
 FILLCELL_X2 FILLER_92_60 ();
 FILLCELL_X8 FILLER_92_66 ();
 FILLCELL_X4 FILLER_92_74 ();
 FILLCELL_X1 FILLER_92_78 ();
 FILLCELL_X2 FILLER_92_101 ();
 FILLCELL_X4 FILLER_92_117 ();
 FILLCELL_X1 FILLER_92_121 ();
 FILLCELL_X8 FILLER_92_136 ();
 FILLCELL_X1 FILLER_92_165 ();
 FILLCELL_X4 FILLER_92_173 ();
 FILLCELL_X4 FILLER_92_190 ();
 FILLCELL_X1 FILLER_92_194 ();
 FILLCELL_X16 FILLER_92_202 ();
 FILLCELL_X8 FILLER_92_218 ();
 FILLCELL_X4 FILLER_92_226 ();
 FILLCELL_X2 FILLER_92_239 ();
 FILLCELL_X8 FILLER_92_262 ();
 FILLCELL_X4 FILLER_92_270 ();
 FILLCELL_X1 FILLER_92_274 ();
 FILLCELL_X8 FILLER_92_283 ();
 FILLCELL_X1 FILLER_92_291 ();
 FILLCELL_X8 FILLER_92_299 ();
 FILLCELL_X4 FILLER_92_307 ();
 FILLCELL_X2 FILLER_92_311 ();
 FILLCELL_X32 FILLER_92_320 ();
 FILLCELL_X8 FILLER_92_352 ();
 FILLCELL_X2 FILLER_92_360 ();
 FILLCELL_X1 FILLER_92_362 ();
 FILLCELL_X8 FILLER_92_366 ();
 FILLCELL_X4 FILLER_92_374 ();
 FILLCELL_X2 FILLER_92_378 ();
 FILLCELL_X1 FILLER_92_400 ();
 FILLCELL_X1 FILLER_92_423 ();
 FILLCELL_X4 FILLER_92_428 ();
 FILLCELL_X2 FILLER_92_432 ();
 FILLCELL_X1 FILLER_92_441 ();
 FILLCELL_X16 FILLER_92_456 ();
 FILLCELL_X8 FILLER_92_472 ();
 FILLCELL_X4 FILLER_92_480 ();
 FILLCELL_X2 FILLER_92_484 ();
 FILLCELL_X1 FILLER_92_486 ();
 FILLCELL_X8 FILLER_92_511 ();
 FILLCELL_X2 FILLER_92_519 ();
 FILLCELL_X1 FILLER_92_521 ();
 FILLCELL_X8 FILLER_92_541 ();
 FILLCELL_X4 FILLER_92_549 ();
 FILLCELL_X2 FILLER_92_553 ();
 FILLCELL_X1 FILLER_92_555 ();
 FILLCELL_X4 FILLER_92_578 ();
 FILLCELL_X8 FILLER_92_601 ();
 FILLCELL_X2 FILLER_92_609 ();
 FILLCELL_X1 FILLER_92_611 ();
 FILLCELL_X16 FILLER_92_632 ();
 FILLCELL_X4 FILLER_92_648 ();
 FILLCELL_X16 FILLER_92_702 ();
 FILLCELL_X1 FILLER_92_718 ();
 FILLCELL_X8 FILLER_92_721 ();
 FILLCELL_X1 FILLER_92_729 ();
 FILLCELL_X4 FILLER_92_732 ();
 FILLCELL_X2 FILLER_92_736 ();
 FILLCELL_X4 FILLER_92_756 ();
 FILLCELL_X1 FILLER_92_760 ();
 FILLCELL_X8 FILLER_92_767 ();
 FILLCELL_X4 FILLER_92_775 ();
 FILLCELL_X2 FILLER_92_785 ();
 FILLCELL_X1 FILLER_92_799 ();
 FILLCELL_X16 FILLER_92_858 ();
 FILLCELL_X1 FILLER_92_874 ();
 FILLCELL_X1 FILLER_92_891 ();
 FILLCELL_X1 FILLER_92_902 ();
 FILLCELL_X1 FILLER_92_919 ();
 FILLCELL_X4 FILLER_92_933 ();
 FILLCELL_X16 FILLER_92_957 ();
 FILLCELL_X8 FILLER_92_973 ();
 FILLCELL_X1 FILLER_92_981 ();
 FILLCELL_X2 FILLER_93_1 ();
 FILLCELL_X8 FILLER_93_23 ();
 FILLCELL_X1 FILLER_93_31 ();
 FILLCELL_X4 FILLER_93_35 ();
 FILLCELL_X1 FILLER_93_39 ();
 FILLCELL_X8 FILLER_93_43 ();
 FILLCELL_X4 FILLER_93_51 ();
 FILLCELL_X2 FILLER_93_55 ();
 FILLCELL_X1 FILLER_93_63 ();
 FILLCELL_X1 FILLER_93_84 ();
 FILLCELL_X4 FILLER_93_114 ();
 FILLCELL_X2 FILLER_93_118 ();
 FILLCELL_X1 FILLER_93_127 ();
 FILLCELL_X2 FILLER_93_135 ();
 FILLCELL_X2 FILLER_93_144 ();
 FILLCELL_X2 FILLER_93_155 ();
 FILLCELL_X1 FILLER_93_157 ();
 FILLCELL_X4 FILLER_93_180 ();
 FILLCELL_X2 FILLER_93_184 ();
 FILLCELL_X1 FILLER_93_186 ();
 FILLCELL_X1 FILLER_93_201 ();
 FILLCELL_X2 FILLER_93_209 ();
 FILLCELL_X4 FILLER_93_220 ();
 FILLCELL_X2 FILLER_93_224 ();
 FILLCELL_X16 FILLER_93_233 ();
 FILLCELL_X8 FILLER_93_249 ();
 FILLCELL_X8 FILLER_93_283 ();
 FILLCELL_X4 FILLER_93_291 ();
 FILLCELL_X1 FILLER_93_340 ();
 FILLCELL_X1 FILLER_93_348 ();
 FILLCELL_X1 FILLER_93_354 ();
 FILLCELL_X1 FILLER_93_360 ();
 FILLCELL_X4 FILLER_93_377 ();
 FILLCELL_X2 FILLER_93_381 ();
 FILLCELL_X4 FILLER_93_392 ();
 FILLCELL_X2 FILLER_93_396 ();
 FILLCELL_X4 FILLER_93_403 ();
 FILLCELL_X2 FILLER_93_407 ();
 FILLCELL_X1 FILLER_93_420 ();
 FILLCELL_X2 FILLER_93_451 ();
 FILLCELL_X32 FILLER_93_460 ();
 FILLCELL_X2 FILLER_93_497 ();
 FILLCELL_X16 FILLER_93_506 ();
 FILLCELL_X4 FILLER_93_522 ();
 FILLCELL_X8 FILLER_93_545 ();
 FILLCELL_X4 FILLER_93_553 ();
 FILLCELL_X2 FILLER_93_557 ();
 FILLCELL_X1 FILLER_93_584 ();
 FILLCELL_X2 FILLER_93_598 ();
 FILLCELL_X1 FILLER_93_600 ();
 FILLCELL_X2 FILLER_93_612 ();
 FILLCELL_X1 FILLER_93_614 ();
 FILLCELL_X4 FILLER_93_626 ();
 FILLCELL_X2 FILLER_93_630 ();
 FILLCELL_X16 FILLER_93_641 ();
 FILLCELL_X4 FILLER_93_657 ();
 FILLCELL_X2 FILLER_93_661 ();
 FILLCELL_X2 FILLER_93_685 ();
 FILLCELL_X16 FILLER_93_694 ();
 FILLCELL_X8 FILLER_93_710 ();
 FILLCELL_X2 FILLER_93_718 ();
 FILLCELL_X4 FILLER_93_730 ();
 FILLCELL_X2 FILLER_93_734 ();
 FILLCELL_X4 FILLER_93_742 ();
 FILLCELL_X2 FILLER_93_746 ();
 FILLCELL_X1 FILLER_93_748 ();
 FILLCELL_X16 FILLER_93_760 ();
 FILLCELL_X4 FILLER_93_776 ();
 FILLCELL_X2 FILLER_93_780 ();
 FILLCELL_X32 FILLER_93_785 ();
 FILLCELL_X8 FILLER_93_817 ();
 FILLCELL_X32 FILLER_93_831 ();
 FILLCELL_X32 FILLER_93_889 ();
 FILLCELL_X32 FILLER_93_921 ();
 FILLCELL_X16 FILLER_93_953 ();
 FILLCELL_X8 FILLER_93_969 ();
 FILLCELL_X4 FILLER_93_977 ();
 FILLCELL_X1 FILLER_93_981 ();
 FILLCELL_X1 FILLER_94_1 ();
 FILLCELL_X2 FILLER_94_5 ();
 FILLCELL_X1 FILLER_94_7 ();
 FILLCELL_X2 FILLER_94_11 ();
 FILLCELL_X1 FILLER_94_13 ();
 FILLCELL_X8 FILLER_94_25 ();
 FILLCELL_X1 FILLER_94_33 ();
 FILLCELL_X4 FILLER_94_56 ();
 FILLCELL_X2 FILLER_94_60 ();
 FILLCELL_X1 FILLER_94_62 ();
 FILLCELL_X8 FILLER_94_67 ();
 FILLCELL_X4 FILLER_94_75 ();
 FILLCELL_X1 FILLER_94_105 ();
 FILLCELL_X4 FILLER_94_120 ();
 FILLCELL_X1 FILLER_94_124 ();
 FILLCELL_X8 FILLER_94_132 ();
 FILLCELL_X1 FILLER_94_140 ();
 FILLCELL_X32 FILLER_94_162 ();
 FILLCELL_X1 FILLER_94_208 ();
 FILLCELL_X4 FILLER_94_229 ();
 FILLCELL_X16 FILLER_94_247 ();
 FILLCELL_X4 FILLER_94_263 ();
 FILLCELL_X2 FILLER_94_267 ();
 FILLCELL_X1 FILLER_94_269 ();
 FILLCELL_X32 FILLER_94_291 ();
 FILLCELL_X1 FILLER_94_323 ();
 FILLCELL_X4 FILLER_94_359 ();
 FILLCELL_X2 FILLER_94_363 ();
 FILLCELL_X1 FILLER_94_394 ();
 FILLCELL_X4 FILLER_94_400 ();
 FILLCELL_X4 FILLER_94_411 ();
 FILLCELL_X8 FILLER_94_418 ();
 FILLCELL_X1 FILLER_94_426 ();
 FILLCELL_X8 FILLER_94_434 ();
 FILLCELL_X4 FILLER_94_442 ();
 FILLCELL_X2 FILLER_94_457 ();
 FILLCELL_X2 FILLER_94_485 ();
 FILLCELL_X1 FILLER_94_487 ();
 FILLCELL_X8 FILLER_94_513 ();
 FILLCELL_X1 FILLER_94_521 ();
 FILLCELL_X1 FILLER_94_528 ();
 FILLCELL_X8 FILLER_94_541 ();
 FILLCELL_X2 FILLER_94_549 ();
 FILLCELL_X1 FILLER_94_551 ();
 FILLCELL_X4 FILLER_94_607 ();
 FILLCELL_X1 FILLER_94_611 ();
 FILLCELL_X2 FILLER_94_632 ();
 FILLCELL_X1 FILLER_94_634 ();
 FILLCELL_X4 FILLER_94_646 ();
 FILLCELL_X2 FILLER_94_650 ();
 FILLCELL_X8 FILLER_94_663 ();
 FILLCELL_X2 FILLER_94_671 ();
 FILLCELL_X1 FILLER_94_673 ();
 FILLCELL_X16 FILLER_94_695 ();
 FILLCELL_X1 FILLER_94_711 ();
 FILLCELL_X2 FILLER_94_741 ();
 FILLCELL_X1 FILLER_94_743 ();
 FILLCELL_X2 FILLER_94_747 ();
 FILLCELL_X1 FILLER_94_749 ();
 FILLCELL_X4 FILLER_94_766 ();
 FILLCELL_X2 FILLER_94_773 ();
 FILLCELL_X1 FILLER_94_775 ();
 FILLCELL_X4 FILLER_94_792 ();
 FILLCELL_X2 FILLER_94_796 ();
 FILLCELL_X1 FILLER_94_798 ();
 FILLCELL_X2 FILLER_94_801 ();
 FILLCELL_X32 FILLER_94_806 ();
 FILLCELL_X32 FILLER_94_838 ();
 FILLCELL_X4 FILLER_94_870 ();
 FILLCELL_X2 FILLER_94_874 ();
 FILLCELL_X1 FILLER_94_886 ();
 FILLCELL_X8 FILLER_94_905 ();
 FILLCELL_X4 FILLER_94_913 ();
 FILLCELL_X1 FILLER_94_917 ();
 FILLCELL_X4 FILLER_94_928 ();
 FILLCELL_X32 FILLER_94_948 ();
 FILLCELL_X2 FILLER_94_980 ();
 FILLCELL_X16 FILLER_95_1 ();
 FILLCELL_X2 FILLER_95_17 ();
 FILLCELL_X8 FILLER_95_25 ();
 FILLCELL_X4 FILLER_95_33 ();
 FILLCELL_X1 FILLER_95_37 ();
 FILLCELL_X2 FILLER_95_47 ();
 FILLCELL_X1 FILLER_95_49 ();
 FILLCELL_X4 FILLER_95_53 ();
 FILLCELL_X16 FILLER_95_60 ();
 FILLCELL_X4 FILLER_95_76 ();
 FILLCELL_X32 FILLER_95_85 ();
 FILLCELL_X32 FILLER_95_117 ();
 FILLCELL_X1 FILLER_95_149 ();
 FILLCELL_X2 FILLER_95_173 ();
 FILLCELL_X1 FILLER_95_175 ();
 FILLCELL_X16 FILLER_95_190 ();
 FILLCELL_X8 FILLER_95_206 ();
 FILLCELL_X4 FILLER_95_214 ();
 FILLCELL_X2 FILLER_95_218 ();
 FILLCELL_X1 FILLER_95_250 ();
 FILLCELL_X4 FILLER_95_267 ();
 FILLCELL_X2 FILLER_95_271 ();
 FILLCELL_X1 FILLER_95_273 ();
 FILLCELL_X2 FILLER_95_297 ();
 FILLCELL_X32 FILLER_95_304 ();
 FILLCELL_X2 FILLER_95_336 ();
 FILLCELL_X1 FILLER_95_338 ();
 FILLCELL_X2 FILLER_95_348 ();
 FILLCELL_X4 FILLER_95_355 ();
 FILLCELL_X1 FILLER_95_359 ();
 FILLCELL_X8 FILLER_95_367 ();
 FILLCELL_X1 FILLER_95_375 ();
 FILLCELL_X2 FILLER_95_388 ();
 FILLCELL_X4 FILLER_95_397 ();
 FILLCELL_X1 FILLER_95_401 ();
 FILLCELL_X2 FILLER_95_409 ();
 FILLCELL_X2 FILLER_95_415 ();
 FILLCELL_X1 FILLER_95_427 ();
 FILLCELL_X2 FILLER_95_444 ();
 FILLCELL_X1 FILLER_95_446 ();
 FILLCELL_X8 FILLER_95_461 ();
 FILLCELL_X1 FILLER_95_469 ();
 FILLCELL_X8 FILLER_95_489 ();
 FILLCELL_X1 FILLER_95_497 ();
 FILLCELL_X8 FILLER_95_540 ();
 FILLCELL_X4 FILLER_95_548 ();
 FILLCELL_X1 FILLER_95_552 ();
 FILLCELL_X16 FILLER_95_582 ();
 FILLCELL_X4 FILLER_95_626 ();
 FILLCELL_X8 FILLER_95_691 ();
 FILLCELL_X4 FILLER_95_699 ();
 FILLCELL_X1 FILLER_95_703 ();
 FILLCELL_X8 FILLER_95_711 ();
 FILLCELL_X4 FILLER_95_719 ();
 FILLCELL_X2 FILLER_95_723 ();
 FILLCELL_X1 FILLER_95_725 ();
 FILLCELL_X1 FILLER_95_734 ();
 FILLCELL_X4 FILLER_95_740 ();
 FILLCELL_X2 FILLER_95_744 ();
 FILLCELL_X1 FILLER_95_746 ();
 FILLCELL_X2 FILLER_95_749 ();
 FILLCELL_X8 FILLER_95_769 ();
 FILLCELL_X8 FILLER_95_781 ();
 FILLCELL_X1 FILLER_95_789 ();
 FILLCELL_X8 FILLER_95_816 ();
 FILLCELL_X4 FILLER_95_824 ();
 FILLCELL_X1 FILLER_95_828 ();
 FILLCELL_X1 FILLER_95_837 ();
 FILLCELL_X1 FILLER_95_856 ();
 FILLCELL_X2 FILLER_95_873 ();
 FILLCELL_X2 FILLER_95_877 ();
 FILLCELL_X2 FILLER_95_895 ();
 FILLCELL_X4 FILLER_95_926 ();
 FILLCELL_X1 FILLER_95_930 ();
 FILLCELL_X4 FILLER_95_933 ();
 FILLCELL_X2 FILLER_95_947 ();
 FILLCELL_X16 FILLER_95_951 ();
 FILLCELL_X8 FILLER_95_967 ();
 FILLCELL_X4 FILLER_95_975 ();
 FILLCELL_X2 FILLER_95_979 ();
 FILLCELL_X1 FILLER_95_981 ();
 FILLCELL_X2 FILLER_96_4 ();
 FILLCELL_X1 FILLER_96_6 ();
 FILLCELL_X8 FILLER_96_62 ();
 FILLCELL_X4 FILLER_96_70 ();
 FILLCELL_X2 FILLER_96_74 ();
 FILLCELL_X8 FILLER_96_108 ();
 FILLCELL_X2 FILLER_96_116 ();
 FILLCELL_X1 FILLER_96_118 ();
 FILLCELL_X16 FILLER_96_133 ();
 FILLCELL_X1 FILLER_96_149 ();
 FILLCELL_X2 FILLER_96_157 ();
 FILLCELL_X1 FILLER_96_159 ();
 FILLCELL_X4 FILLER_96_167 ();
 FILLCELL_X2 FILLER_96_171 ();
 FILLCELL_X2 FILLER_96_186 ();
 FILLCELL_X1 FILLER_96_188 ();
 FILLCELL_X4 FILLER_96_196 ();
 FILLCELL_X2 FILLER_96_200 ();
 FILLCELL_X8 FILLER_96_215 ();
 FILLCELL_X1 FILLER_96_223 ();
 FILLCELL_X4 FILLER_96_238 ();
 FILLCELL_X2 FILLER_96_242 ();
 FILLCELL_X1 FILLER_96_251 ();
 FILLCELL_X8 FILLER_96_259 ();
 FILLCELL_X1 FILLER_96_267 ();
 FILLCELL_X2 FILLER_96_281 ();
 FILLCELL_X1 FILLER_96_305 ();
 FILLCELL_X8 FILLER_96_323 ();
 FILLCELL_X1 FILLER_96_331 ();
 FILLCELL_X2 FILLER_96_339 ();
 FILLCELL_X16 FILLER_96_348 ();
 FILLCELL_X8 FILLER_96_364 ();
 FILLCELL_X4 FILLER_96_372 ();
 FILLCELL_X2 FILLER_96_376 ();
 FILLCELL_X1 FILLER_96_378 ();
 FILLCELL_X4 FILLER_96_396 ();
 FILLCELL_X2 FILLER_96_400 ();
 FILLCELL_X1 FILLER_96_402 ();
 FILLCELL_X4 FILLER_96_422 ();
 FILLCELL_X2 FILLER_96_426 ();
 FILLCELL_X1 FILLER_96_428 ();
 FILLCELL_X16 FILLER_96_458 ();
 FILLCELL_X4 FILLER_96_480 ();
 FILLCELL_X16 FILLER_96_489 ();
 FILLCELL_X4 FILLER_96_505 ();
 FILLCELL_X2 FILLER_96_509 ();
 FILLCELL_X1 FILLER_96_511 ();
 FILLCELL_X8 FILLER_96_517 ();
 FILLCELL_X4 FILLER_96_525 ();
 FILLCELL_X32 FILLER_96_536 ();
 FILLCELL_X8 FILLER_96_568 ();
 FILLCELL_X4 FILLER_96_576 ();
 FILLCELL_X1 FILLER_96_580 ();
 FILLCELL_X8 FILLER_96_588 ();
 FILLCELL_X1 FILLER_96_596 ();
 FILLCELL_X4 FILLER_96_617 ();
 FILLCELL_X1 FILLER_96_621 ();
 FILLCELL_X4 FILLER_96_632 ();
 FILLCELL_X1 FILLER_96_636 ();
 FILLCELL_X4 FILLER_96_673 ();
 FILLCELL_X2 FILLER_96_677 ();
 FILLCELL_X1 FILLER_96_679 ();
 FILLCELL_X16 FILLER_96_716 ();
 FILLCELL_X8 FILLER_96_732 ();
 FILLCELL_X4 FILLER_96_740 ();
 FILLCELL_X2 FILLER_96_744 ();
 FILLCELL_X1 FILLER_96_746 ();
 FILLCELL_X2 FILLER_96_759 ();
 FILLCELL_X2 FILLER_96_777 ();
 FILLCELL_X8 FILLER_96_795 ();
 FILLCELL_X1 FILLER_96_803 ();
 FILLCELL_X1 FILLER_96_839 ();
 FILLCELL_X4 FILLER_96_858 ();
 FILLCELL_X2 FILLER_96_862 ();
 FILLCELL_X16 FILLER_96_880 ();
 FILLCELL_X2 FILLER_96_896 ();
 FILLCELL_X1 FILLER_96_898 ();
 FILLCELL_X8 FILLER_96_901 ();
 FILLCELL_X4 FILLER_96_909 ();
 FILLCELL_X2 FILLER_96_913 ();
 FILLCELL_X1 FILLER_96_915 ();
 FILLCELL_X4 FILLER_96_918 ();
 FILLCELL_X8 FILLER_96_941 ();
 FILLCELL_X8 FILLER_96_967 ();
 FILLCELL_X4 FILLER_96_975 ();
 FILLCELL_X2 FILLER_96_979 ();
 FILLCELL_X1 FILLER_96_981 ();
 FILLCELL_X8 FILLER_97_27 ();
 FILLCELL_X4 FILLER_97_35 ();
 FILLCELL_X2 FILLER_97_39 ();
 FILLCELL_X1 FILLER_97_41 ();
 FILLCELL_X8 FILLER_97_45 ();
 FILLCELL_X4 FILLER_97_53 ();
 FILLCELL_X2 FILLER_97_60 ();
 FILLCELL_X1 FILLER_97_62 ();
 FILLCELL_X8 FILLER_97_66 ();
 FILLCELL_X4 FILLER_97_74 ();
 FILLCELL_X2 FILLER_97_78 ();
 FILLCELL_X1 FILLER_97_80 ();
 FILLCELL_X4 FILLER_97_119 ();
 FILLCELL_X4 FILLER_97_166 ();
 FILLCELL_X2 FILLER_97_170 ();
 FILLCELL_X32 FILLER_97_193 ();
 FILLCELL_X8 FILLER_97_225 ();
 FILLCELL_X4 FILLER_97_233 ();
 FILLCELL_X2 FILLER_97_237 ();
 FILLCELL_X16 FILLER_97_255 ();
 FILLCELL_X2 FILLER_97_271 ();
 FILLCELL_X4 FILLER_97_280 ();
 FILLCELL_X16 FILLER_97_288 ();
 FILLCELL_X4 FILLER_97_311 ();
 FILLCELL_X2 FILLER_97_315 ();
 FILLCELL_X1 FILLER_97_317 ();
 FILLCELL_X4 FILLER_97_339 ();
 FILLCELL_X2 FILLER_97_343 ();
 FILLCELL_X1 FILLER_97_345 ();
 FILLCELL_X2 FILLER_97_353 ();
 FILLCELL_X4 FILLER_97_362 ();
 FILLCELL_X2 FILLER_97_366 ();
 FILLCELL_X1 FILLER_97_368 ();
 FILLCELL_X1 FILLER_97_380 ();
 FILLCELL_X4 FILLER_97_388 ();
 FILLCELL_X2 FILLER_97_392 ();
 FILLCELL_X1 FILLER_97_394 ();
 FILLCELL_X8 FILLER_97_402 ();
 FILLCELL_X4 FILLER_97_410 ();
 FILLCELL_X8 FILLER_97_430 ();
 FILLCELL_X16 FILLER_97_457 ();
 FILLCELL_X4 FILLER_97_473 ();
 FILLCELL_X2 FILLER_97_477 ();
 FILLCELL_X1 FILLER_97_479 ();
 FILLCELL_X8 FILLER_97_494 ();
 FILLCELL_X1 FILLER_97_502 ();
 FILLCELL_X16 FILLER_97_541 ();
 FILLCELL_X2 FILLER_97_557 ();
 FILLCELL_X2 FILLER_97_570 ();
 FILLCELL_X1 FILLER_97_586 ();
 FILLCELL_X2 FILLER_97_656 ();
 FILLCELL_X1 FILLER_97_658 ();
 FILLCELL_X2 FILLER_97_679 ();
 FILLCELL_X1 FILLER_97_681 ();
 FILLCELL_X16 FILLER_97_701 ();
 FILLCELL_X8 FILLER_97_717 ();
 FILLCELL_X2 FILLER_97_734 ();
 FILLCELL_X1 FILLER_97_736 ();
 FILLCELL_X1 FILLER_97_742 ();
 FILLCELL_X2 FILLER_97_775 ();
 FILLCELL_X8 FILLER_97_783 ();
 FILLCELL_X4 FILLER_97_791 ();
 FILLCELL_X1 FILLER_97_795 ();
 FILLCELL_X8 FILLER_97_798 ();
 FILLCELL_X4 FILLER_97_806 ();
 FILLCELL_X2 FILLER_97_810 ();
 FILLCELL_X8 FILLER_97_828 ();
 FILLCELL_X2 FILLER_97_836 ();
 FILLCELL_X4 FILLER_97_840 ();
 FILLCELL_X1 FILLER_97_844 ();
 FILLCELL_X8 FILLER_97_861 ();
 FILLCELL_X1 FILLER_97_869 ();
 FILLCELL_X16 FILLER_97_912 ();
 FILLCELL_X1 FILLER_97_928 ();
 FILLCELL_X8 FILLER_97_971 ();
 FILLCELL_X2 FILLER_97_979 ();
 FILLCELL_X1 FILLER_97_981 ();
 FILLCELL_X4 FILLER_98_1 ();
 FILLCELL_X2 FILLER_98_5 ();
 FILLCELL_X8 FILLER_98_10 ();
 FILLCELL_X2 FILLER_98_18 ();
 FILLCELL_X1 FILLER_98_23 ();
 FILLCELL_X1 FILLER_98_28 ();
 FILLCELL_X8 FILLER_98_50 ();
 FILLCELL_X16 FILLER_98_67 ();
 FILLCELL_X2 FILLER_98_83 ();
 FILLCELL_X1 FILLER_98_102 ();
 FILLCELL_X16 FILLER_98_122 ();
 FILLCELL_X8 FILLER_98_138 ();
 FILLCELL_X2 FILLER_98_146 ();
 FILLCELL_X1 FILLER_98_148 ();
 FILLCELL_X4 FILLER_98_170 ();
 FILLCELL_X2 FILLER_98_174 ();
 FILLCELL_X1 FILLER_98_176 ();
 FILLCELL_X1 FILLER_98_190 ();
 FILLCELL_X4 FILLER_98_200 ();
 FILLCELL_X8 FILLER_98_234 ();
 FILLCELL_X2 FILLER_98_242 ();
 FILLCELL_X1 FILLER_98_251 ();
 FILLCELL_X8 FILLER_98_259 ();
 FILLCELL_X2 FILLER_98_267 ();
 FILLCELL_X32 FILLER_98_316 ();
 FILLCELL_X16 FILLER_98_348 ();
 FILLCELL_X2 FILLER_98_378 ();
 FILLCELL_X8 FILLER_98_387 ();
 FILLCELL_X4 FILLER_98_409 ();
 FILLCELL_X2 FILLER_98_413 ();
 FILLCELL_X4 FILLER_98_429 ();
 FILLCELL_X2 FILLER_98_433 ();
 FILLCELL_X8 FILLER_98_440 ();
 FILLCELL_X2 FILLER_98_448 ();
 FILLCELL_X4 FILLER_98_471 ();
 FILLCELL_X2 FILLER_98_475 ();
 FILLCELL_X1 FILLER_98_477 ();
 FILLCELL_X8 FILLER_98_501 ();
 FILLCELL_X4 FILLER_98_509 ();
 FILLCELL_X2 FILLER_98_513 ();
 FILLCELL_X2 FILLER_98_534 ();
 FILLCELL_X1 FILLER_98_536 ();
 FILLCELL_X2 FILLER_98_546 ();
 FILLCELL_X1 FILLER_98_548 ();
 FILLCELL_X8 FILLER_98_575 ();
 FILLCELL_X8 FILLER_98_592 ();
 FILLCELL_X4 FILLER_98_600 ();
 FILLCELL_X2 FILLER_98_604 ();
 FILLCELL_X2 FILLER_98_613 ();
 FILLCELL_X1 FILLER_98_615 ();
 FILLCELL_X2 FILLER_98_629 ();
 FILLCELL_X4 FILLER_98_632 ();
 FILLCELL_X4 FILLER_98_643 ();
 FILLCELL_X2 FILLER_98_647 ();
 FILLCELL_X1 FILLER_98_649 ();
 FILLCELL_X4 FILLER_98_657 ();
 FILLCELL_X1 FILLER_98_661 ();
 FILLCELL_X16 FILLER_98_691 ();
 FILLCELL_X8 FILLER_98_707 ();
 FILLCELL_X4 FILLER_98_715 ();
 FILLCELL_X8 FILLER_98_738 ();
 FILLCELL_X4 FILLER_98_752 ();
 FILLCELL_X4 FILLER_98_788 ();
 FILLCELL_X1 FILLER_98_792 ();
 FILLCELL_X2 FILLER_98_809 ();
 FILLCELL_X1 FILLER_98_811 ();
 FILLCELL_X16 FILLER_98_814 ();
 FILLCELL_X4 FILLER_98_830 ();
 FILLCELL_X2 FILLER_98_834 ();
 FILLCELL_X8 FILLER_98_852 ();
 FILLCELL_X2 FILLER_98_860 ();
 FILLCELL_X1 FILLER_98_862 ();
 FILLCELL_X4 FILLER_98_881 ();
 FILLCELL_X1 FILLER_98_885 ();
 FILLCELL_X4 FILLER_98_888 ();
 FILLCELL_X2 FILLER_98_892 ();
 FILLCELL_X4 FILLER_98_910 ();
 FILLCELL_X2 FILLER_98_914 ();
 FILLCELL_X1 FILLER_98_916 ();
 FILLCELL_X8 FILLER_98_927 ();
 FILLCELL_X2 FILLER_98_935 ();
 FILLCELL_X4 FILLER_98_959 ();
 FILLCELL_X8 FILLER_98_967 ();
 FILLCELL_X4 FILLER_98_975 ();
 FILLCELL_X2 FILLER_98_979 ();
 FILLCELL_X1 FILLER_98_981 ();
 FILLCELL_X1 FILLER_99_1 ();
 FILLCELL_X1 FILLER_99_5 ();
 FILLCELL_X1 FILLER_99_23 ();
 FILLCELL_X1 FILLER_99_27 ();
 FILLCELL_X16 FILLER_99_32 ();
 FILLCELL_X8 FILLER_99_48 ();
 FILLCELL_X2 FILLER_99_56 ();
 FILLCELL_X1 FILLER_99_61 ();
 FILLCELL_X4 FILLER_99_65 ();
 FILLCELL_X2 FILLER_99_69 ();
 FILLCELL_X1 FILLER_99_71 ();
 FILLCELL_X16 FILLER_99_77 ();
 FILLCELL_X4 FILLER_99_93 ();
 FILLCELL_X1 FILLER_99_97 ();
 FILLCELL_X1 FILLER_99_111 ();
 FILLCELL_X16 FILLER_99_128 ();
 FILLCELL_X4 FILLER_99_147 ();
 FILLCELL_X32 FILLER_99_165 ();
 FILLCELL_X4 FILLER_99_197 ();
 FILLCELL_X2 FILLER_99_201 ();
 FILLCELL_X1 FILLER_99_203 ();
 FILLCELL_X16 FILLER_99_225 ();
 FILLCELL_X4 FILLER_99_241 ();
 FILLCELL_X2 FILLER_99_245 ();
 FILLCELL_X1 FILLER_99_247 ();
 FILLCELL_X8 FILLER_99_262 ();
 FILLCELL_X2 FILLER_99_270 ();
 FILLCELL_X1 FILLER_99_272 ();
 FILLCELL_X2 FILLER_99_289 ();
 FILLCELL_X2 FILLER_99_298 ();
 FILLCELL_X4 FILLER_99_319 ();
 FILLCELL_X16 FILLER_99_330 ();
 FILLCELL_X4 FILLER_99_346 ();
 FILLCELL_X2 FILLER_99_350 ();
 FILLCELL_X2 FILLER_99_359 ();
 FILLCELL_X1 FILLER_99_361 ();
 FILLCELL_X2 FILLER_99_382 ();
 FILLCELL_X4 FILLER_99_411 ();
 FILLCELL_X2 FILLER_99_415 ();
 FILLCELL_X16 FILLER_99_424 ();
 FILLCELL_X4 FILLER_99_440 ();
 FILLCELL_X4 FILLER_99_465 ();
 FILLCELL_X1 FILLER_99_469 ();
 FILLCELL_X4 FILLER_99_499 ();
 FILLCELL_X1 FILLER_99_510 ();
 FILLCELL_X16 FILLER_99_520 ();
 FILLCELL_X4 FILLER_99_536 ();
 FILLCELL_X2 FILLER_99_540 ();
 FILLCELL_X16 FILLER_99_549 ();
 FILLCELL_X2 FILLER_99_565 ();
 FILLCELL_X8 FILLER_99_574 ();
 FILLCELL_X2 FILLER_99_591 ();
 FILLCELL_X1 FILLER_99_593 ();
 FILLCELL_X2 FILLER_99_603 ();
 FILLCELL_X16 FILLER_99_612 ();
 FILLCELL_X2 FILLER_99_628 ();
 FILLCELL_X1 FILLER_99_630 ();
 FILLCELL_X4 FILLER_99_645 ();
 FILLCELL_X2 FILLER_99_649 ();
 FILLCELL_X1 FILLER_99_651 ();
 FILLCELL_X4 FILLER_99_666 ();
 FILLCELL_X2 FILLER_99_700 ();
 FILLCELL_X16 FILLER_99_705 ();
 FILLCELL_X2 FILLER_99_721 ();
 FILLCELL_X1 FILLER_99_723 ();
 FILLCELL_X16 FILLER_99_728 ();
 FILLCELL_X8 FILLER_99_744 ();
 FILLCELL_X4 FILLER_99_752 ();
 FILLCELL_X2 FILLER_99_756 ();
 FILLCELL_X2 FILLER_99_763 ();
 FILLCELL_X2 FILLER_99_767 ();
 FILLCELL_X8 FILLER_99_771 ();
 FILLCELL_X4 FILLER_99_779 ();
 FILLCELL_X8 FILLER_99_788 ();
 FILLCELL_X4 FILLER_99_796 ();
 FILLCELL_X2 FILLER_99_800 ();
 FILLCELL_X16 FILLER_99_818 ();
 FILLCELL_X4 FILLER_99_836 ();
 FILLCELL_X2 FILLER_99_840 ();
 FILLCELL_X2 FILLER_99_844 ();
 FILLCELL_X8 FILLER_99_866 ();
 FILLCELL_X2 FILLER_99_874 ();
 FILLCELL_X4 FILLER_99_886 ();
 FILLCELL_X2 FILLER_99_890 ();
 FILLCELL_X4 FILLER_99_902 ();
 FILLCELL_X2 FILLER_99_906 ();
 FILLCELL_X1 FILLER_99_940 ();
 FILLCELL_X1 FILLER_99_951 ();
 FILLCELL_X8 FILLER_99_968 ();
 FILLCELL_X4 FILLER_99_976 ();
 FILLCELL_X2 FILLER_99_980 ();
 FILLCELL_X4 FILLER_100_1 ();
 FILLCELL_X1 FILLER_100_5 ();
 FILLCELL_X2 FILLER_100_9 ();
 FILLCELL_X4 FILLER_100_52 ();
 FILLCELL_X2 FILLER_100_56 ();
 FILLCELL_X1 FILLER_100_58 ();
 FILLCELL_X1 FILLER_100_85 ();
 FILLCELL_X4 FILLER_100_90 ();
 FILLCELL_X2 FILLER_100_94 ();
 FILLCELL_X1 FILLER_100_96 ();
 FILLCELL_X1 FILLER_100_103 ();
 FILLCELL_X4 FILLER_100_117 ();
 FILLCELL_X4 FILLER_100_140 ();
 FILLCELL_X8 FILLER_100_150 ();
 FILLCELL_X4 FILLER_100_158 ();
 FILLCELL_X1 FILLER_100_162 ();
 FILLCELL_X1 FILLER_100_198 ();
 FILLCELL_X8 FILLER_100_206 ();
 FILLCELL_X4 FILLER_100_214 ();
 FILLCELL_X2 FILLER_100_218 ();
 FILLCELL_X1 FILLER_100_220 ();
 FILLCELL_X4 FILLER_100_228 ();
 FILLCELL_X2 FILLER_100_232 ();
 FILLCELL_X1 FILLER_100_234 ();
 FILLCELL_X4 FILLER_100_248 ();
 FILLCELL_X1 FILLER_100_252 ();
 FILLCELL_X2 FILLER_100_256 ();
 FILLCELL_X1 FILLER_100_258 ();
 FILLCELL_X32 FILLER_100_266 ();
 FILLCELL_X16 FILLER_100_298 ();
 FILLCELL_X2 FILLER_100_314 ();
 FILLCELL_X1 FILLER_100_316 ();
 FILLCELL_X8 FILLER_100_340 ();
 FILLCELL_X4 FILLER_100_348 ();
 FILLCELL_X1 FILLER_100_352 ();
 FILLCELL_X2 FILLER_100_381 ();
 FILLCELL_X8 FILLER_100_403 ();
 FILLCELL_X16 FILLER_100_425 ();
 FILLCELL_X2 FILLER_100_441 ();
 FILLCELL_X2 FILLER_100_459 ();
 FILLCELL_X1 FILLER_100_461 ();
 FILLCELL_X8 FILLER_100_465 ();
 FILLCELL_X4 FILLER_100_473 ();
 FILLCELL_X1 FILLER_100_477 ();
 FILLCELL_X8 FILLER_100_485 ();
 FILLCELL_X4 FILLER_100_517 ();
 FILLCELL_X2 FILLER_100_521 ();
 FILLCELL_X2 FILLER_100_532 ();
 FILLCELL_X1 FILLER_100_534 ();
 FILLCELL_X2 FILLER_100_542 ();
 FILLCELL_X8 FILLER_100_551 ();
 FILLCELL_X1 FILLER_100_559 ();
 FILLCELL_X2 FILLER_100_566 ();
 FILLCELL_X4 FILLER_100_575 ();
 FILLCELL_X1 FILLER_100_579 ();
 FILLCELL_X4 FILLER_100_587 ();
 FILLCELL_X2 FILLER_100_591 ();
 FILLCELL_X1 FILLER_100_593 ();
 FILLCELL_X2 FILLER_100_601 ();
 FILLCELL_X4 FILLER_100_610 ();
 FILLCELL_X2 FILLER_100_614 ();
 FILLCELL_X8 FILLER_100_623 ();
 FILLCELL_X4 FILLER_100_639 ();
 FILLCELL_X1 FILLER_100_643 ();
 FILLCELL_X8 FILLER_100_651 ();
 FILLCELL_X4 FILLER_100_659 ();
 FILLCELL_X1 FILLER_100_663 ();
 FILLCELL_X2 FILLER_100_678 ();
 FILLCELL_X32 FILLER_100_701 ();
 FILLCELL_X16 FILLER_100_733 ();
 FILLCELL_X4 FILLER_100_751 ();
 FILLCELL_X1 FILLER_100_755 ();
 FILLCELL_X8 FILLER_100_793 ();
 FILLCELL_X2 FILLER_100_801 ();
 FILLCELL_X1 FILLER_100_803 ();
 FILLCELL_X32 FILLER_100_822 ();
 FILLCELL_X16 FILLER_100_854 ();
 FILLCELL_X8 FILLER_100_870 ();
 FILLCELL_X4 FILLER_100_878 ();
 FILLCELL_X16 FILLER_100_884 ();
 FILLCELL_X8 FILLER_100_900 ();
 FILLCELL_X16 FILLER_100_918 ();
 FILLCELL_X16 FILLER_100_936 ();
 FILLCELL_X4 FILLER_100_952 ();
 FILLCELL_X2 FILLER_100_956 ();
 FILLCELL_X1 FILLER_100_958 ();
 FILLCELL_X1 FILLER_100_961 ();
 FILLCELL_X8 FILLER_100_972 ();
 FILLCELL_X2 FILLER_100_980 ();
 FILLCELL_X4 FILLER_101_1 ();
 FILLCELL_X2 FILLER_101_5 ();
 FILLCELL_X1 FILLER_101_7 ();
 FILLCELL_X1 FILLER_101_17 ();
 FILLCELL_X8 FILLER_101_25 ();
 FILLCELL_X1 FILLER_101_33 ();
 FILLCELL_X1 FILLER_101_37 ();
 FILLCELL_X4 FILLER_101_42 ();
 FILLCELL_X2 FILLER_101_49 ();
 FILLCELL_X1 FILLER_101_51 ();
 FILLCELL_X1 FILLER_101_72 ();
 FILLCELL_X16 FILLER_101_77 ();
 FILLCELL_X1 FILLER_101_93 ();
 FILLCELL_X1 FILLER_101_111 ();
 FILLCELL_X8 FILLER_101_161 ();
 FILLCELL_X2 FILLER_101_169 ();
 FILLCELL_X1 FILLER_101_171 ();
 FILLCELL_X16 FILLER_101_181 ();
 FILLCELL_X1 FILLER_101_197 ();
 FILLCELL_X8 FILLER_101_219 ();
 FILLCELL_X4 FILLER_101_227 ();
 FILLCELL_X4 FILLER_101_252 ();
 FILLCELL_X8 FILLER_101_265 ();
 FILLCELL_X2 FILLER_101_273 ();
 FILLCELL_X1 FILLER_101_275 ();
 FILLCELL_X4 FILLER_101_285 ();
 FILLCELL_X2 FILLER_101_289 ();
 FILLCELL_X8 FILLER_101_298 ();
 FILLCELL_X1 FILLER_101_306 ();
 FILLCELL_X8 FILLER_101_310 ();
 FILLCELL_X1 FILLER_101_318 ();
 FILLCELL_X2 FILLER_101_366 ();
 FILLCELL_X2 FILLER_101_396 ();
 FILLCELL_X4 FILLER_101_419 ();
 FILLCELL_X4 FILLER_101_433 ();
 FILLCELL_X1 FILLER_101_437 ();
 FILLCELL_X8 FILLER_101_452 ();
 FILLCELL_X16 FILLER_101_467 ();
 FILLCELL_X8 FILLER_101_483 ();
 FILLCELL_X4 FILLER_101_491 ();
 FILLCELL_X8 FILLER_101_522 ();
 FILLCELL_X4 FILLER_101_530 ();
 FILLCELL_X1 FILLER_101_534 ();
 FILLCELL_X16 FILLER_101_580 ();
 FILLCELL_X1 FILLER_101_596 ();
 FILLCELL_X16 FILLER_101_611 ();
 FILLCELL_X4 FILLER_101_627 ();
 FILLCELL_X1 FILLER_101_631 ();
 FILLCELL_X1 FILLER_101_646 ();
 FILLCELL_X4 FILLER_101_665 ();
 FILLCELL_X16 FILLER_101_676 ();
 FILLCELL_X1 FILLER_101_692 ();
 FILLCELL_X4 FILLER_101_706 ();
 FILLCELL_X16 FILLER_101_734 ();
 FILLCELL_X8 FILLER_101_750 ();
 FILLCELL_X4 FILLER_101_758 ();
 FILLCELL_X1 FILLER_101_762 ();
 FILLCELL_X2 FILLER_101_780 ();
 FILLCELL_X1 FILLER_101_782 ();
 FILLCELL_X2 FILLER_101_786 ();
 FILLCELL_X1 FILLER_101_788 ();
 FILLCELL_X2 FILLER_101_796 ();
 FILLCELL_X1 FILLER_101_798 ();
 FILLCELL_X16 FILLER_101_815 ();
 FILLCELL_X2 FILLER_101_831 ();
 FILLCELL_X1 FILLER_101_833 ();
 FILLCELL_X8 FILLER_101_850 ();
 FILLCELL_X4 FILLER_101_858 ();
 FILLCELL_X32 FILLER_101_878 ();
 FILLCELL_X8 FILLER_101_910 ();
 FILLCELL_X2 FILLER_101_928 ();
 FILLCELL_X16 FILLER_101_962 ();
 FILLCELL_X4 FILLER_101_978 ();
 FILLCELL_X16 FILLER_102_1 ();
 FILLCELL_X8 FILLER_102_34 ();
 FILLCELL_X2 FILLER_102_42 ();
 FILLCELL_X2 FILLER_102_47 ();
 FILLCELL_X4 FILLER_102_66 ();
 FILLCELL_X16 FILLER_102_74 ();
 FILLCELL_X8 FILLER_102_90 ();
 FILLCELL_X1 FILLER_102_98 ();
 FILLCELL_X4 FILLER_102_104 ();
 FILLCELL_X2 FILLER_102_108 ();
 FILLCELL_X1 FILLER_102_110 ();
 FILLCELL_X8 FILLER_102_123 ();
 FILLCELL_X4 FILLER_102_131 ();
 FILLCELL_X16 FILLER_102_164 ();
 FILLCELL_X4 FILLER_102_180 ();
 FILLCELL_X2 FILLER_102_198 ();
 FILLCELL_X1 FILLER_102_200 ();
 FILLCELL_X2 FILLER_102_204 ();
 FILLCELL_X1 FILLER_102_206 ();
 FILLCELL_X2 FILLER_102_214 ();
 FILLCELL_X1 FILLER_102_216 ();
 FILLCELL_X8 FILLER_102_224 ();
 FILLCELL_X4 FILLER_102_232 ();
 FILLCELL_X1 FILLER_102_236 ();
 FILLCELL_X4 FILLER_102_258 ();
 FILLCELL_X2 FILLER_102_262 ();
 FILLCELL_X4 FILLER_102_271 ();
 FILLCELL_X1 FILLER_102_275 ();
 FILLCELL_X1 FILLER_102_295 ();
 FILLCELL_X8 FILLER_102_306 ();
 FILLCELL_X4 FILLER_102_314 ();
 FILLCELL_X2 FILLER_102_318 ();
 FILLCELL_X1 FILLER_102_327 ();
 FILLCELL_X1 FILLER_102_335 ();
 FILLCELL_X1 FILLER_102_349 ();
 FILLCELL_X1 FILLER_102_409 ();
 FILLCELL_X2 FILLER_102_424 ();
 FILLCELL_X1 FILLER_102_426 ();
 FILLCELL_X4 FILLER_102_441 ();
 FILLCELL_X2 FILLER_102_445 ();
 FILLCELL_X2 FILLER_102_460 ();
 FILLCELL_X4 FILLER_102_489 ();
 FILLCELL_X2 FILLER_102_493 ();
 FILLCELL_X1 FILLER_102_495 ();
 FILLCELL_X2 FILLER_102_503 ();
 FILLCELL_X1 FILLER_102_505 ();
 FILLCELL_X32 FILLER_102_516 ();
 FILLCELL_X4 FILLER_102_548 ();
 FILLCELL_X16 FILLER_102_565 ();
 FILLCELL_X8 FILLER_102_581 ();
 FILLCELL_X4 FILLER_102_589 ();
 FILLCELL_X1 FILLER_102_593 ();
 FILLCELL_X4 FILLER_102_619 ();
 FILLCELL_X1 FILLER_102_623 ();
 FILLCELL_X4 FILLER_102_632 ();
 FILLCELL_X1 FILLER_102_636 ();
 FILLCELL_X8 FILLER_102_659 ();
 FILLCELL_X2 FILLER_102_667 ();
 FILLCELL_X1 FILLER_102_669 ();
 FILLCELL_X2 FILLER_102_680 ();
 FILLCELL_X1 FILLER_102_696 ();
 FILLCELL_X8 FILLER_102_707 ();
 FILLCELL_X4 FILLER_102_715 ();
 FILLCELL_X2 FILLER_102_723 ();
 FILLCELL_X1 FILLER_102_725 ();
 FILLCELL_X16 FILLER_102_729 ();
 FILLCELL_X8 FILLER_102_745 ();
 FILLCELL_X4 FILLER_102_753 ();
 FILLCELL_X2 FILLER_102_772 ();
 FILLCELL_X4 FILLER_102_783 ();
 FILLCELL_X2 FILLER_102_787 ();
 FILLCELL_X1 FILLER_102_789 ();
 FILLCELL_X2 FILLER_102_793 ();
 FILLCELL_X4 FILLER_102_811 ();
 FILLCELL_X1 FILLER_102_815 ();
 FILLCELL_X8 FILLER_102_832 ();
 FILLCELL_X2 FILLER_102_840 ();
 FILLCELL_X2 FILLER_102_860 ();
 FILLCELL_X2 FILLER_102_872 ();
 FILLCELL_X1 FILLER_102_890 ();
 FILLCELL_X2 FILLER_102_893 ();
 FILLCELL_X1 FILLER_102_895 ();
 FILLCELL_X2 FILLER_102_912 ();
 FILLCELL_X1 FILLER_102_914 ();
 FILLCELL_X1 FILLER_102_931 ();
 FILLCELL_X4 FILLER_102_944 ();
 FILLCELL_X2 FILLER_102_948 ();
 FILLCELL_X1 FILLER_102_950 ();
 FILLCELL_X8 FILLER_102_969 ();
 FILLCELL_X4 FILLER_102_977 ();
 FILLCELL_X1 FILLER_102_981 ();
 FILLCELL_X8 FILLER_103_1 ();
 FILLCELL_X4 FILLER_103_9 ();
 FILLCELL_X2 FILLER_103_16 ();
 FILLCELL_X1 FILLER_103_18 ();
 FILLCELL_X8 FILLER_103_22 ();
 FILLCELL_X2 FILLER_103_30 ();
 FILLCELL_X16 FILLER_103_35 ();
 FILLCELL_X4 FILLER_103_51 ();
 FILLCELL_X2 FILLER_103_55 ();
 FILLCELL_X1 FILLER_103_57 ();
 FILLCELL_X2 FILLER_103_61 ();
 FILLCELL_X4 FILLER_103_67 ();
 FILLCELL_X2 FILLER_103_71 ();
 FILLCELL_X8 FILLER_103_93 ();
 FILLCELL_X1 FILLER_103_101 ();
 FILLCELL_X1 FILLER_103_111 ();
 FILLCELL_X16 FILLER_103_121 ();
 FILLCELL_X4 FILLER_103_137 ();
 FILLCELL_X4 FILLER_103_148 ();
 FILLCELL_X2 FILLER_103_152 ();
 FILLCELL_X1 FILLER_103_154 ();
 FILLCELL_X8 FILLER_103_165 ();
 FILLCELL_X2 FILLER_103_173 ();
 FILLCELL_X1 FILLER_103_175 ();
 FILLCELL_X8 FILLER_103_190 ();
 FILLCELL_X4 FILLER_103_198 ();
 FILLCELL_X16 FILLER_103_216 ();
 FILLCELL_X4 FILLER_103_232 ();
 FILLCELL_X2 FILLER_103_236 ();
 FILLCELL_X8 FILLER_103_245 ();
 FILLCELL_X4 FILLER_103_253 ();
 FILLCELL_X1 FILLER_103_257 ();
 FILLCELL_X2 FILLER_103_265 ();
 FILLCELL_X1 FILLER_103_267 ();
 FILLCELL_X8 FILLER_103_278 ();
 FILLCELL_X2 FILLER_103_286 ();
 FILLCELL_X1 FILLER_103_288 ();
 FILLCELL_X16 FILLER_103_299 ();
 FILLCELL_X4 FILLER_103_315 ();
 FILLCELL_X2 FILLER_103_319 ();
 FILLCELL_X4 FILLER_103_328 ();
 FILLCELL_X1 FILLER_103_332 ();
 FILLCELL_X4 FILLER_103_405 ();
 FILLCELL_X2 FILLER_103_409 ();
 FILLCELL_X4 FILLER_103_425 ();
 FILLCELL_X2 FILLER_103_429 ();
 FILLCELL_X1 FILLER_103_431 ();
 FILLCELL_X4 FILLER_103_440 ();
 FILLCELL_X1 FILLER_103_444 ();
 FILLCELL_X4 FILLER_103_452 ();
 FILLCELL_X2 FILLER_103_456 ();
 FILLCELL_X1 FILLER_103_474 ();
 FILLCELL_X8 FILLER_103_489 ();
 FILLCELL_X2 FILLER_103_497 ();
 FILLCELL_X1 FILLER_103_499 ();
 FILLCELL_X2 FILLER_103_507 ();
 FILLCELL_X1 FILLER_103_509 ();
 FILLCELL_X2 FILLER_103_513 ();
 FILLCELL_X8 FILLER_103_524 ();
 FILLCELL_X4 FILLER_103_532 ();
 FILLCELL_X16 FILLER_103_553 ();
 FILLCELL_X2 FILLER_103_569 ();
 FILLCELL_X16 FILLER_103_578 ();
 FILLCELL_X4 FILLER_103_594 ();
 FILLCELL_X1 FILLER_103_598 ();
 FILLCELL_X16 FILLER_103_606 ();
 FILLCELL_X1 FILLER_103_622 ();
 FILLCELL_X4 FILLER_103_644 ();
 FILLCELL_X2 FILLER_103_648 ();
 FILLCELL_X1 FILLER_103_650 ();
 FILLCELL_X16 FILLER_103_672 ();
 FILLCELL_X2 FILLER_103_688 ();
 FILLCELL_X16 FILLER_103_697 ();
 FILLCELL_X2 FILLER_103_713 ();
 FILLCELL_X1 FILLER_103_715 ();
 FILLCELL_X16 FILLER_103_733 ();
 FILLCELL_X2 FILLER_103_749 ();
 FILLCELL_X1 FILLER_103_751 ();
 FILLCELL_X1 FILLER_103_758 ();
 FILLCELL_X2 FILLER_103_764 ();
 FILLCELL_X8 FILLER_103_801 ();
 FILLCELL_X1 FILLER_103_809 ();
 FILLCELL_X8 FILLER_103_812 ();
 FILLCELL_X4 FILLER_103_820 ();
 FILLCELL_X2 FILLER_103_824 ();
 FILLCELL_X1 FILLER_103_836 ();
 FILLCELL_X4 FILLER_103_839 ();
 FILLCELL_X8 FILLER_103_855 ();
 FILLCELL_X16 FILLER_103_881 ();
 FILLCELL_X2 FILLER_103_897 ();
 FILLCELL_X1 FILLER_103_899 ();
 FILLCELL_X32 FILLER_103_902 ();
 FILLCELL_X16 FILLER_103_934 ();
 FILLCELL_X8 FILLER_103_950 ();
 FILLCELL_X2 FILLER_103_958 ();
 FILLCELL_X4 FILLER_103_976 ();
 FILLCELL_X2 FILLER_103_980 ();
 FILLCELL_X1 FILLER_104_1 ();
 FILLCELL_X1 FILLER_104_19 ();
 FILLCELL_X4 FILLER_104_45 ();
 FILLCELL_X2 FILLER_104_49 ();
 FILLCELL_X1 FILLER_104_51 ();
 FILLCELL_X4 FILLER_104_58 ();
 FILLCELL_X2 FILLER_104_62 ();
 FILLCELL_X1 FILLER_104_64 ();
 FILLCELL_X8 FILLER_104_68 ();
 FILLCELL_X2 FILLER_104_76 ();
 FILLCELL_X1 FILLER_104_95 ();
 FILLCELL_X4 FILLER_104_137 ();
 FILLCELL_X8 FILLER_104_144 ();
 FILLCELL_X2 FILLER_104_152 ();
 FILLCELL_X4 FILLER_104_157 ();
 FILLCELL_X2 FILLER_104_161 ();
 FILLCELL_X2 FILLER_104_176 ();
 FILLCELL_X1 FILLER_104_178 ();
 FILLCELL_X1 FILLER_104_182 ();
 FILLCELL_X16 FILLER_104_186 ();
 FILLCELL_X2 FILLER_104_202 ();
 FILLCELL_X8 FILLER_104_214 ();
 FILLCELL_X4 FILLER_104_222 ();
 FILLCELL_X16 FILLER_104_229 ();
 FILLCELL_X8 FILLER_104_250 ();
 FILLCELL_X4 FILLER_104_258 ();
 FILLCELL_X1 FILLER_104_262 ();
 FILLCELL_X1 FILLER_104_273 ();
 FILLCELL_X2 FILLER_104_281 ();
 FILLCELL_X1 FILLER_104_283 ();
 FILLCELL_X2 FILLER_104_287 ();
 FILLCELL_X1 FILLER_104_289 ();
 FILLCELL_X16 FILLER_104_304 ();
 FILLCELL_X8 FILLER_104_327 ();
 FILLCELL_X1 FILLER_104_335 ();
 FILLCELL_X2 FILLER_104_339 ();
 FILLCELL_X1 FILLER_104_341 ();
 FILLCELL_X2 FILLER_104_349 ();
 FILLCELL_X2 FILLER_104_364 ();
 FILLCELL_X1 FILLER_104_366 ();
 FILLCELL_X1 FILLER_104_394 ();
 FILLCELL_X1 FILLER_104_398 ();
 FILLCELL_X1 FILLER_104_419 ();
 FILLCELL_X2 FILLER_104_432 ();
 FILLCELL_X1 FILLER_104_434 ();
 FILLCELL_X4 FILLER_104_442 ();
 FILLCELL_X8 FILLER_104_453 ();
 FILLCELL_X4 FILLER_104_461 ();
 FILLCELL_X1 FILLER_104_465 ();
 FILLCELL_X8 FILLER_104_473 ();
 FILLCELL_X16 FILLER_104_484 ();
 FILLCELL_X2 FILLER_104_507 ();
 FILLCELL_X1 FILLER_104_509 ();
 FILLCELL_X1 FILLER_104_517 ();
 FILLCELL_X8 FILLER_104_521 ();
 FILLCELL_X2 FILLER_104_529 ();
 FILLCELL_X1 FILLER_104_531 ();
 FILLCELL_X8 FILLER_104_546 ();
 FILLCELL_X4 FILLER_104_554 ();
 FILLCELL_X2 FILLER_104_558 ();
 FILLCELL_X1 FILLER_104_560 ();
 FILLCELL_X4 FILLER_104_585 ();
 FILLCELL_X16 FILLER_104_603 ();
 FILLCELL_X8 FILLER_104_619 ();
 FILLCELL_X4 FILLER_104_627 ();
 FILLCELL_X4 FILLER_104_653 ();
 FILLCELL_X2 FILLER_104_657 ();
 FILLCELL_X2 FILLER_104_666 ();
 FILLCELL_X1 FILLER_104_668 ();
 FILLCELL_X2 FILLER_104_676 ();
 FILLCELL_X8 FILLER_104_699 ();
 FILLCELL_X4 FILLER_104_707 ();
 FILLCELL_X2 FILLER_104_711 ();
 FILLCELL_X16 FILLER_104_720 ();
 FILLCELL_X8 FILLER_104_736 ();
 FILLCELL_X4 FILLER_104_744 ();
 FILLCELL_X2 FILLER_104_748 ();
 FILLCELL_X1 FILLER_104_750 ();
 FILLCELL_X8 FILLER_104_757 ();
 FILLCELL_X2 FILLER_104_765 ();
 FILLCELL_X1 FILLER_104_767 ();
 FILLCELL_X4 FILLER_104_785 ();
 FILLCELL_X1 FILLER_104_789 ();
 FILLCELL_X16 FILLER_104_793 ();
 FILLCELL_X2 FILLER_104_809 ();
 FILLCELL_X32 FILLER_104_829 ();
 FILLCELL_X8 FILLER_104_861 ();
 FILLCELL_X1 FILLER_104_869 ();
 FILLCELL_X4 FILLER_104_872 ();
 FILLCELL_X2 FILLER_104_876 ();
 FILLCELL_X1 FILLER_104_878 ();
 FILLCELL_X4 FILLER_104_889 ();
 FILLCELL_X2 FILLER_104_893 ();
 FILLCELL_X2 FILLER_104_911 ();
 FILLCELL_X16 FILLER_104_915 ();
 FILLCELL_X8 FILLER_104_931 ();
 FILLCELL_X4 FILLER_104_939 ();
 FILLCELL_X8 FILLER_104_953 ();
 FILLCELL_X2 FILLER_104_961 ();
 FILLCELL_X1 FILLER_104_973 ();
 FILLCELL_X4 FILLER_104_976 ();
 FILLCELL_X2 FILLER_104_980 ();
 FILLCELL_X8 FILLER_105_1 ();
 FILLCELL_X4 FILLER_105_12 ();
 FILLCELL_X1 FILLER_105_19 ();
 FILLCELL_X1 FILLER_105_23 ();
 FILLCELL_X8 FILLER_105_28 ();
 FILLCELL_X4 FILLER_105_36 ();
 FILLCELL_X1 FILLER_105_72 ();
 FILLCELL_X4 FILLER_105_93 ();
 FILLCELL_X2 FILLER_105_97 ();
 FILLCELL_X1 FILLER_105_99 ();
 FILLCELL_X16 FILLER_105_122 ();
 FILLCELL_X2 FILLER_105_138 ();
 FILLCELL_X1 FILLER_105_140 ();
 FILLCELL_X4 FILLER_105_144 ();
 FILLCELL_X1 FILLER_105_148 ();
 FILLCELL_X1 FILLER_105_163 ();
 FILLCELL_X2 FILLER_105_191 ();
 FILLCELL_X4 FILLER_105_224 ();
 FILLCELL_X2 FILLER_105_228 ();
 FILLCELL_X8 FILLER_105_247 ();
 FILLCELL_X2 FILLER_105_262 ();
 FILLCELL_X1 FILLER_105_271 ();
 FILLCELL_X1 FILLER_105_279 ();
 FILLCELL_X8 FILLER_105_287 ();
 FILLCELL_X1 FILLER_105_295 ();
 FILLCELL_X8 FILLER_105_315 ();
 FILLCELL_X1 FILLER_105_323 ();
 FILLCELL_X8 FILLER_105_338 ();
 FILLCELL_X2 FILLER_105_346 ();
 FILLCELL_X2 FILLER_105_360 ();
 FILLCELL_X1 FILLER_105_362 ();
 FILLCELL_X2 FILLER_105_366 ();
 FILLCELL_X1 FILLER_105_368 ();
 FILLCELL_X32 FILLER_105_376 ();
 FILLCELL_X2 FILLER_105_408 ();
 FILLCELL_X16 FILLER_105_417 ();
 FILLCELL_X4 FILLER_105_433 ();
 FILLCELL_X2 FILLER_105_437 ();
 FILLCELL_X8 FILLER_105_458 ();
 FILLCELL_X2 FILLER_105_466 ();
 FILLCELL_X16 FILLER_105_475 ();
 FILLCELL_X8 FILLER_105_491 ();
 FILLCELL_X4 FILLER_105_499 ();
 FILLCELL_X1 FILLER_105_503 ();
 FILLCELL_X4 FILLER_105_518 ();
 FILLCELL_X1 FILLER_105_522 ();
 FILLCELL_X4 FILLER_105_530 ();
 FILLCELL_X2 FILLER_105_534 ();
 FILLCELL_X16 FILLER_105_546 ();
 FILLCELL_X2 FILLER_105_562 ();
 FILLCELL_X1 FILLER_105_580 ();
 FILLCELL_X4 FILLER_105_588 ();
 FILLCELL_X2 FILLER_105_592 ();
 FILLCELL_X1 FILLER_105_594 ();
 FILLCELL_X8 FILLER_105_616 ();
 FILLCELL_X1 FILLER_105_624 ();
 FILLCELL_X4 FILLER_105_684 ();
 FILLCELL_X2 FILLER_105_688 ();
 FILLCELL_X1 FILLER_105_690 ();
 FILLCELL_X1 FILLER_105_704 ();
 FILLCELL_X32 FILLER_105_722 ();
 FILLCELL_X2 FILLER_105_754 ();
 FILLCELL_X4 FILLER_105_761 ();
 FILLCELL_X1 FILLER_105_791 ();
 FILLCELL_X16 FILLER_105_802 ();
 FILLCELL_X4 FILLER_105_834 ();
 FILLCELL_X2 FILLER_105_838 ();
 FILLCELL_X16 FILLER_105_843 ();
 FILLCELL_X8 FILLER_105_859 ();
 FILLCELL_X2 FILLER_105_867 ();
 FILLCELL_X1 FILLER_105_892 ();
 FILLCELL_X2 FILLER_105_905 ();
 FILLCELL_X1 FILLER_105_907 ();
 FILLCELL_X32 FILLER_105_924 ();
 FILLCELL_X1 FILLER_105_956 ();
 FILLCELL_X4 FILLER_105_959 ();
 FILLCELL_X8 FILLER_105_973 ();
 FILLCELL_X1 FILLER_105_981 ();
 FILLCELL_X4 FILLER_106_1 ();
 FILLCELL_X4 FILLER_106_8 ();
 FILLCELL_X2 FILLER_106_12 ();
 FILLCELL_X8 FILLER_106_31 ();
 FILLCELL_X4 FILLER_106_39 ();
 FILLCELL_X2 FILLER_106_43 ();
 FILLCELL_X1 FILLER_106_45 ();
 FILLCELL_X4 FILLER_106_70 ();
 FILLCELL_X1 FILLER_106_74 ();
 FILLCELL_X16 FILLER_106_118 ();
 FILLCELL_X4 FILLER_106_134 ();
 FILLCELL_X1 FILLER_106_138 ();
 FILLCELL_X16 FILLER_106_160 ();
 FILLCELL_X2 FILLER_106_176 ();
 FILLCELL_X8 FILLER_106_185 ();
 FILLCELL_X4 FILLER_106_193 ();
 FILLCELL_X1 FILLER_106_197 ();
 FILLCELL_X4 FILLER_106_208 ();
 FILLCELL_X4 FILLER_106_236 ();
 FILLCELL_X1 FILLER_106_240 ();
 FILLCELL_X4 FILLER_106_248 ();
 FILLCELL_X1 FILLER_106_252 ();
 FILLCELL_X8 FILLER_106_274 ();
 FILLCELL_X2 FILLER_106_282 ();
 FILLCELL_X1 FILLER_106_284 ();
 FILLCELL_X2 FILLER_106_292 ();
 FILLCELL_X1 FILLER_106_294 ();
 FILLCELL_X16 FILLER_106_310 ();
 FILLCELL_X4 FILLER_106_326 ();
 FILLCELL_X1 FILLER_106_330 ();
 FILLCELL_X1 FILLER_106_339 ();
 FILLCELL_X1 FILLER_106_343 ();
 FILLCELL_X4 FILLER_106_351 ();
 FILLCELL_X2 FILLER_106_355 ();
 FILLCELL_X1 FILLER_106_357 ();
 FILLCELL_X1 FILLER_106_368 ();
 FILLCELL_X8 FILLER_106_387 ();
 FILLCELL_X4 FILLER_106_395 ();
 FILLCELL_X2 FILLER_106_399 ();
 FILLCELL_X4 FILLER_106_415 ();
 FILLCELL_X1 FILLER_106_419 ();
 FILLCELL_X16 FILLER_106_427 ();
 FILLCELL_X4 FILLER_106_443 ();
 FILLCELL_X2 FILLER_106_447 ();
 FILLCELL_X8 FILLER_106_454 ();
 FILLCELL_X2 FILLER_106_462 ();
 FILLCELL_X1 FILLER_106_464 ();
 FILLCELL_X4 FILLER_106_471 ();
 FILLCELL_X2 FILLER_106_489 ();
 FILLCELL_X1 FILLER_106_491 ();
 FILLCELL_X2 FILLER_106_499 ();
 FILLCELL_X1 FILLER_106_501 ();
 FILLCELL_X1 FILLER_106_505 ();
 FILLCELL_X2 FILLER_106_509 ();
 FILLCELL_X2 FILLER_106_518 ();
 FILLCELL_X2 FILLER_106_533 ();
 FILLCELL_X4 FILLER_106_552 ();
 FILLCELL_X1 FILLER_106_556 ();
 FILLCELL_X8 FILLER_106_578 ();
 FILLCELL_X4 FILLER_106_586 ();
 FILLCELL_X2 FILLER_106_590 ();
 FILLCELL_X1 FILLER_106_592 ();
 FILLCELL_X4 FILLER_106_607 ();
 FILLCELL_X2 FILLER_106_611 ();
 FILLCELL_X1 FILLER_106_613 ();
 FILLCELL_X8 FILLER_106_619 ();
 FILLCELL_X4 FILLER_106_627 ();
 FILLCELL_X4 FILLER_106_632 ();
 FILLCELL_X2 FILLER_106_636 ();
 FILLCELL_X8 FILLER_106_657 ();
 FILLCELL_X8 FILLER_106_679 ();
 FILLCELL_X4 FILLER_106_687 ();
 FILLCELL_X1 FILLER_106_698 ();
 FILLCELL_X1 FILLER_106_705 ();
 FILLCELL_X2 FILLER_106_709 ();
 FILLCELL_X8 FILLER_106_714 ();
 FILLCELL_X16 FILLER_106_729 ();
 FILLCELL_X4 FILLER_106_745 ();
 FILLCELL_X8 FILLER_106_758 ();
 FILLCELL_X1 FILLER_106_791 ();
 FILLCELL_X2 FILLER_106_794 ();
 FILLCELL_X4 FILLER_106_812 ();
 FILLCELL_X2 FILLER_106_816 ();
 FILLCELL_X2 FILLER_106_831 ();
 FILLCELL_X4 FILLER_106_849 ();
 FILLCELL_X2 FILLER_106_853 ();
 FILLCELL_X1 FILLER_106_855 ();
 FILLCELL_X4 FILLER_106_866 ();
 FILLCELL_X2 FILLER_106_870 ();
 FILLCELL_X1 FILLER_106_872 ();
 FILLCELL_X16 FILLER_106_875 ();
 FILLCELL_X8 FILLER_106_891 ();
 FILLCELL_X2 FILLER_106_899 ();
 FILLCELL_X1 FILLER_106_919 ();
 FILLCELL_X8 FILLER_106_954 ();
 FILLCELL_X1 FILLER_106_962 ();
 FILLCELL_X8 FILLER_106_973 ();
 FILLCELL_X1 FILLER_106_981 ();
 FILLCELL_X8 FILLER_107_7 ();
 FILLCELL_X1 FILLER_107_15 ();
 FILLCELL_X1 FILLER_107_22 ();
 FILLCELL_X2 FILLER_107_27 ();
 FILLCELL_X16 FILLER_107_37 ();
 FILLCELL_X8 FILLER_107_53 ();
 FILLCELL_X4 FILLER_107_61 ();
 FILLCELL_X16 FILLER_107_68 ();
 FILLCELL_X8 FILLER_107_84 ();
 FILLCELL_X2 FILLER_107_92 ();
 FILLCELL_X1 FILLER_107_94 ();
 FILLCELL_X8 FILLER_107_127 ();
 FILLCELL_X1 FILLER_107_135 ();
 FILLCELL_X2 FILLER_107_157 ();
 FILLCELL_X1 FILLER_107_159 ();
 FILLCELL_X8 FILLER_107_167 ();
 FILLCELL_X4 FILLER_107_175 ();
 FILLCELL_X8 FILLER_107_189 ();
 FILLCELL_X2 FILLER_107_197 ();
 FILLCELL_X32 FILLER_107_202 ();
 FILLCELL_X1 FILLER_107_234 ();
 FILLCELL_X4 FILLER_107_242 ();
 FILLCELL_X1 FILLER_107_253 ();
 FILLCELL_X16 FILLER_107_268 ();
 FILLCELL_X8 FILLER_107_284 ();
 FILLCELL_X4 FILLER_107_292 ();
 FILLCELL_X2 FILLER_107_296 ();
 FILLCELL_X8 FILLER_107_317 ();
 FILLCELL_X4 FILLER_107_325 ();
 FILLCELL_X1 FILLER_107_329 ();
 FILLCELL_X8 FILLER_107_337 ();
 FILLCELL_X2 FILLER_107_345 ();
 FILLCELL_X1 FILLER_107_347 ();
 FILLCELL_X2 FILLER_107_368 ();
 FILLCELL_X2 FILLER_107_383 ();
 FILLCELL_X4 FILLER_107_390 ();
 FILLCELL_X2 FILLER_107_394 ();
 FILLCELL_X4 FILLER_107_410 ();
 FILLCELL_X1 FILLER_107_414 ();
 FILLCELL_X2 FILLER_107_436 ();
 FILLCELL_X8 FILLER_107_452 ();
 FILLCELL_X2 FILLER_107_460 ();
 FILLCELL_X8 FILLER_107_476 ();
 FILLCELL_X4 FILLER_107_484 ();
 FILLCELL_X2 FILLER_107_488 ();
 FILLCELL_X1 FILLER_107_490 ();
 FILLCELL_X4 FILLER_107_505 ();
 FILLCELL_X1 FILLER_107_523 ();
 FILLCELL_X16 FILLER_107_538 ();
 FILLCELL_X8 FILLER_107_554 ();
 FILLCELL_X4 FILLER_107_562 ();
 FILLCELL_X2 FILLER_107_566 ();
 FILLCELL_X1 FILLER_107_568 ();
 FILLCELL_X2 FILLER_107_583 ();
 FILLCELL_X32 FILLER_107_599 ();
 FILLCELL_X4 FILLER_107_631 ();
 FILLCELL_X4 FILLER_107_663 ();
 FILLCELL_X2 FILLER_107_667 ();
 FILLCELL_X1 FILLER_107_669 ();
 FILLCELL_X1 FILLER_107_688 ();
 FILLCELL_X1 FILLER_107_698 ();
 FILLCELL_X2 FILLER_107_702 ();
 FILLCELL_X1 FILLER_107_704 ();
 FILLCELL_X8 FILLER_107_711 ();
 FILLCELL_X1 FILLER_107_719 ();
 FILLCELL_X8 FILLER_107_737 ();
 FILLCELL_X1 FILLER_107_745 ();
 FILLCELL_X8 FILLER_107_780 ();
 FILLCELL_X4 FILLER_107_792 ();
 FILLCELL_X2 FILLER_107_796 ();
 FILLCELL_X8 FILLER_107_816 ();
 FILLCELL_X1 FILLER_107_824 ();
 FILLCELL_X1 FILLER_107_827 ();
 FILLCELL_X8 FILLER_107_846 ();
 FILLCELL_X32 FILLER_107_866 ();
 FILLCELL_X32 FILLER_107_898 ();
 FILLCELL_X2 FILLER_107_930 ();
 FILLCELL_X8 FILLER_107_934 ();
 FILLCELL_X4 FILLER_107_942 ();
 FILLCELL_X2 FILLER_107_946 ();
 FILLCELL_X1 FILLER_107_948 ();
 FILLCELL_X16 FILLER_107_959 ();
 FILLCELL_X4 FILLER_107_975 ();
 FILLCELL_X2 FILLER_107_979 ();
 FILLCELL_X1 FILLER_107_981 ();
 FILLCELL_X1 FILLER_108_1 ();
 FILLCELL_X1 FILLER_108_19 ();
 FILLCELL_X8 FILLER_108_37 ();
 FILLCELL_X4 FILLER_108_45 ();
 FILLCELL_X2 FILLER_108_49 ();
 FILLCELL_X16 FILLER_108_55 ();
 FILLCELL_X4 FILLER_108_71 ();
 FILLCELL_X2 FILLER_108_75 ();
 FILLCELL_X1 FILLER_108_77 ();
 FILLCELL_X1 FILLER_108_98 ();
 FILLCELL_X8 FILLER_108_119 ();
 FILLCELL_X8 FILLER_108_141 ();
 FILLCELL_X2 FILLER_108_149 ();
 FILLCELL_X1 FILLER_108_151 ();
 FILLCELL_X1 FILLER_108_180 ();
 FILLCELL_X16 FILLER_108_209 ();
 FILLCELL_X4 FILLER_108_225 ();
 FILLCELL_X16 FILLER_108_231 ();
 FILLCELL_X4 FILLER_108_247 ();
 FILLCELL_X2 FILLER_108_251 ();
 FILLCELL_X16 FILLER_108_257 ();
 FILLCELL_X2 FILLER_108_273 ();
 FILLCELL_X1 FILLER_108_275 ();
 FILLCELL_X2 FILLER_108_287 ();
 FILLCELL_X1 FILLER_108_289 ();
 FILLCELL_X4 FILLER_108_294 ();
 FILLCELL_X1 FILLER_108_298 ();
 FILLCELL_X2 FILLER_108_306 ();
 FILLCELL_X4 FILLER_108_311 ();
 FILLCELL_X2 FILLER_108_315 ();
 FILLCELL_X1 FILLER_108_317 ();
 FILLCELL_X8 FILLER_108_322 ();
 FILLCELL_X2 FILLER_108_330 ();
 FILLCELL_X1 FILLER_108_332 ();
 FILLCELL_X32 FILLER_108_341 ();
 FILLCELL_X16 FILLER_108_373 ();
 FILLCELL_X2 FILLER_108_389 ();
 FILLCELL_X4 FILLER_108_408 ();
 FILLCELL_X4 FILLER_108_433 ();
 FILLCELL_X2 FILLER_108_437 ();
 FILLCELL_X1 FILLER_108_439 ();
 FILLCELL_X2 FILLER_108_447 ();
 FILLCELL_X4 FILLER_108_470 ();
 FILLCELL_X2 FILLER_108_474 ();
 FILLCELL_X1 FILLER_108_476 ();
 FILLCELL_X16 FILLER_108_486 ();
 FILLCELL_X1 FILLER_108_502 ();
 FILLCELL_X16 FILLER_108_506 ();
 FILLCELL_X16 FILLER_108_536 ();
 FILLCELL_X8 FILLER_108_552 ();
 FILLCELL_X4 FILLER_108_560 ();
 FILLCELL_X1 FILLER_108_564 ();
 FILLCELL_X2 FILLER_108_572 ();
 FILLCELL_X1 FILLER_108_574 ();
 FILLCELL_X8 FILLER_108_582 ();
 FILLCELL_X4 FILLER_108_597 ();
 FILLCELL_X4 FILLER_108_605 ();
 FILLCELL_X2 FILLER_108_629 ();
 FILLCELL_X4 FILLER_108_645 ();
 FILLCELL_X1 FILLER_108_649 ();
 FILLCELL_X1 FILLER_108_679 ();
 FILLCELL_X32 FILLER_108_697 ();
 FILLCELL_X32 FILLER_108_729 ();
 FILLCELL_X8 FILLER_108_761 ();
 FILLCELL_X1 FILLER_108_769 ();
 FILLCELL_X2 FILLER_108_802 ();
 FILLCELL_X8 FILLER_108_823 ();
 FILLCELL_X1 FILLER_108_831 ();
 FILLCELL_X1 FILLER_108_861 ();
 FILLCELL_X1 FILLER_108_922 ();
 FILLCELL_X8 FILLER_108_939 ();
 FILLCELL_X1 FILLER_108_947 ();
 FILLCELL_X4 FILLER_108_958 ();
 FILLCELL_X8 FILLER_108_974 ();
 FILLCELL_X2 FILLER_109_1 ();
 FILLCELL_X2 FILLER_109_6 ();
 FILLCELL_X1 FILLER_109_8 ();
 FILLCELL_X2 FILLER_109_25 ();
 FILLCELL_X4 FILLER_109_30 ();
 FILLCELL_X2 FILLER_109_58 ();
 FILLCELL_X8 FILLER_109_67 ();
 FILLCELL_X2 FILLER_109_75 ();
 FILLCELL_X8 FILLER_109_126 ();
 FILLCELL_X2 FILLER_109_134 ();
 FILLCELL_X4 FILLER_109_168 ();
 FILLCELL_X16 FILLER_109_179 ();
 FILLCELL_X4 FILLER_109_195 ();
 FILLCELL_X2 FILLER_109_199 ();
 FILLCELL_X1 FILLER_109_201 ();
 FILLCELL_X2 FILLER_109_227 ();
 FILLCELL_X2 FILLER_109_253 ();
 FILLCELL_X4 FILLER_109_269 ();
 FILLCELL_X2 FILLER_109_273 ();
 FILLCELL_X8 FILLER_109_316 ();
 FILLCELL_X2 FILLER_109_324 ();
 FILLCELL_X1 FILLER_109_326 ();
 FILLCELL_X1 FILLER_109_338 ();
 FILLCELL_X8 FILLER_109_358 ();
 FILLCELL_X4 FILLER_109_375 ();
 FILLCELL_X2 FILLER_109_379 ();
 FILLCELL_X1 FILLER_109_381 ();
 FILLCELL_X1 FILLER_109_395 ();
 FILLCELL_X4 FILLER_109_401 ();
 FILLCELL_X4 FILLER_109_419 ();
 FILLCELL_X1 FILLER_109_423 ();
 FILLCELL_X16 FILLER_109_443 ();
 FILLCELL_X8 FILLER_109_459 ();
 FILLCELL_X4 FILLER_109_467 ();
 FILLCELL_X4 FILLER_109_482 ();
 FILLCELL_X4 FILLER_109_526 ();
 FILLCELL_X2 FILLER_109_530 ();
 FILLCELL_X1 FILLER_109_532 ();
 FILLCELL_X8 FILLER_109_542 ();
 FILLCELL_X1 FILLER_109_550 ();
 FILLCELL_X4 FILLER_109_568 ();
 FILLCELL_X2 FILLER_109_572 ();
 FILLCELL_X4 FILLER_109_585 ();
 FILLCELL_X2 FILLER_109_589 ();
 FILLCELL_X8 FILLER_109_605 ();
 FILLCELL_X2 FILLER_109_632 ();
 FILLCELL_X1 FILLER_109_634 ();
 FILLCELL_X4 FILLER_109_655 ();
 FILLCELL_X1 FILLER_109_659 ();
 FILLCELL_X32 FILLER_109_708 ();
 FILLCELL_X32 FILLER_109_740 ();
 FILLCELL_X2 FILLER_109_776 ();
 FILLCELL_X4 FILLER_109_780 ();
 FILLCELL_X2 FILLER_109_784 ();
 FILLCELL_X1 FILLER_109_786 ();
 FILLCELL_X16 FILLER_109_799 ();
 FILLCELL_X4 FILLER_109_815 ();
 FILLCELL_X8 FILLER_109_837 ();
 FILLCELL_X2 FILLER_109_845 ();
 FILLCELL_X1 FILLER_109_847 ();
 FILLCELL_X1 FILLER_109_850 ();
 FILLCELL_X16 FILLER_109_853 ();
 FILLCELL_X8 FILLER_109_869 ();
 FILLCELL_X2 FILLER_109_877 ();
 FILLCELL_X16 FILLER_109_881 ();
 FILLCELL_X4 FILLER_109_897 ();
 FILLCELL_X4 FILLER_109_933 ();
 FILLCELL_X4 FILLER_109_955 ();
 FILLCELL_X2 FILLER_109_959 ();
 FILLCELL_X4 FILLER_109_977 ();
 FILLCELL_X1 FILLER_109_981 ();
 FILLCELL_X1 FILLER_110_1 ();
 FILLCELL_X8 FILLER_110_5 ();
 FILLCELL_X4 FILLER_110_13 ();
 FILLCELL_X16 FILLER_110_34 ();
 FILLCELL_X1 FILLER_110_50 ();
 FILLCELL_X16 FILLER_110_74 ();
 FILLCELL_X2 FILLER_110_90 ();
 FILLCELL_X1 FILLER_110_92 ();
 FILLCELL_X1 FILLER_110_129 ();
 FILLCELL_X32 FILLER_110_144 ();
 FILLCELL_X4 FILLER_110_176 ();
 FILLCELL_X2 FILLER_110_180 ();
 FILLCELL_X2 FILLER_110_191 ();
 FILLCELL_X1 FILLER_110_193 ();
 FILLCELL_X16 FILLER_110_203 ();
 FILLCELL_X8 FILLER_110_219 ();
 FILLCELL_X2 FILLER_110_227 ();
 FILLCELL_X1 FILLER_110_229 ();
 FILLCELL_X4 FILLER_110_249 ();
 FILLCELL_X1 FILLER_110_253 ();
 FILLCELL_X1 FILLER_110_284 ();
 FILLCELL_X4 FILLER_110_321 ();
 FILLCELL_X1 FILLER_110_325 ();
 FILLCELL_X1 FILLER_110_334 ();
 FILLCELL_X8 FILLER_110_344 ();
 FILLCELL_X2 FILLER_110_352 ();
 FILLCELL_X4 FILLER_110_381 ();
 FILLCELL_X1 FILLER_110_385 ();
 FILLCELL_X2 FILLER_110_405 ();
 FILLCELL_X1 FILLER_110_407 ();
 FILLCELL_X16 FILLER_110_425 ();
 FILLCELL_X4 FILLER_110_441 ();
 FILLCELL_X2 FILLER_110_445 ();
 FILLCELL_X1 FILLER_110_447 ();
 FILLCELL_X8 FILLER_110_455 ();
 FILLCELL_X2 FILLER_110_463 ();
 FILLCELL_X1 FILLER_110_465 ();
 FILLCELL_X4 FILLER_110_483 ();
 FILLCELL_X1 FILLER_110_487 ();
 FILLCELL_X1 FILLER_110_499 ();
 FILLCELL_X4 FILLER_110_511 ();
 FILLCELL_X1 FILLER_110_526 ();
 FILLCELL_X8 FILLER_110_544 ();
 FILLCELL_X4 FILLER_110_552 ();
 FILLCELL_X4 FILLER_110_576 ();
 FILLCELL_X8 FILLER_110_597 ();
 FILLCELL_X1 FILLER_110_605 ();
 FILLCELL_X2 FILLER_110_612 ();
 FILLCELL_X1 FILLER_110_614 ();
 FILLCELL_X2 FILLER_110_620 ();
 FILLCELL_X2 FILLER_110_632 ();
 FILLCELL_X1 FILLER_110_634 ();
 FILLCELL_X4 FILLER_110_665 ();
 FILLCELL_X2 FILLER_110_669 ();
 FILLCELL_X1 FILLER_110_671 ();
 FILLCELL_X8 FILLER_110_689 ();
 FILLCELL_X16 FILLER_110_700 ();
 FILLCELL_X4 FILLER_110_716 ();
 FILLCELL_X2 FILLER_110_720 ();
 FILLCELL_X2 FILLER_110_726 ();
 FILLCELL_X1 FILLER_110_728 ();
 FILLCELL_X16 FILLER_110_733 ();
 FILLCELL_X8 FILLER_110_749 ();
 FILLCELL_X4 FILLER_110_757 ();
 FILLCELL_X2 FILLER_110_761 ();
 FILLCELL_X16 FILLER_110_766 ();
 FILLCELL_X8 FILLER_110_782 ();
 FILLCELL_X1 FILLER_110_790 ();
 FILLCELL_X4 FILLER_110_799 ();
 FILLCELL_X2 FILLER_110_803 ();
 FILLCELL_X1 FILLER_110_805 ();
 FILLCELL_X8 FILLER_110_815 ();
 FILLCELL_X2 FILLER_110_823 ();
 FILLCELL_X8 FILLER_110_841 ();
 FILLCELL_X32 FILLER_110_868 ();
 FILLCELL_X16 FILLER_110_900 ();
 FILLCELL_X2 FILLER_110_916 ();
 FILLCELL_X1 FILLER_110_918 ();
 FILLCELL_X8 FILLER_110_924 ();
 FILLCELL_X4 FILLER_110_932 ();
 FILLCELL_X4 FILLER_110_938 ();
 FILLCELL_X2 FILLER_110_960 ();
 FILLCELL_X1 FILLER_110_962 ();
 FILLCELL_X4 FILLER_110_975 ();
 FILLCELL_X2 FILLER_110_979 ();
 FILLCELL_X1 FILLER_110_981 ();
 FILLCELL_X1 FILLER_111_1 ();
 FILLCELL_X1 FILLER_111_19 ();
 FILLCELL_X1 FILLER_111_36 ();
 FILLCELL_X16 FILLER_111_44 ();
 FILLCELL_X4 FILLER_111_60 ();
 FILLCELL_X1 FILLER_111_64 ();
 FILLCELL_X2 FILLER_111_68 ();
 FILLCELL_X1 FILLER_111_70 ();
 FILLCELL_X16 FILLER_111_74 ();
 FILLCELL_X8 FILLER_111_90 ();
 FILLCELL_X4 FILLER_111_98 ();
 FILLCELL_X32 FILLER_111_110 ();
 FILLCELL_X16 FILLER_111_142 ();
 FILLCELL_X8 FILLER_111_158 ();
 FILLCELL_X1 FILLER_111_166 ();
 FILLCELL_X4 FILLER_111_184 ();
 FILLCELL_X2 FILLER_111_188 ();
 FILLCELL_X16 FILLER_111_207 ();
 FILLCELL_X4 FILLER_111_223 ();
 FILLCELL_X2 FILLER_111_227 ();
 FILLCELL_X2 FILLER_111_263 ();
 FILLCELL_X16 FILLER_111_272 ();
 FILLCELL_X2 FILLER_111_288 ();
 FILLCELL_X1 FILLER_111_290 ();
 FILLCELL_X4 FILLER_111_305 ();
 FILLCELL_X8 FILLER_111_316 ();
 FILLCELL_X1 FILLER_111_324 ();
 FILLCELL_X2 FILLER_111_329 ();
 FILLCELL_X4 FILLER_111_345 ();
 FILLCELL_X2 FILLER_111_349 ();
 FILLCELL_X2 FILLER_111_381 ();
 FILLCELL_X1 FILLER_111_383 ();
 FILLCELL_X1 FILLER_111_414 ();
 FILLCELL_X16 FILLER_111_422 ();
 FILLCELL_X4 FILLER_111_438 ();
 FILLCELL_X4 FILLER_111_476 ();
 FILLCELL_X2 FILLER_111_480 ();
 FILLCELL_X1 FILLER_111_482 ();
 FILLCELL_X16 FILLER_111_530 ();
 FILLCELL_X2 FILLER_111_546 ();
 FILLCELL_X1 FILLER_111_548 ();
 FILLCELL_X4 FILLER_111_606 ();
 FILLCELL_X1 FILLER_111_610 ();
 FILLCELL_X4 FILLER_111_628 ();
 FILLCELL_X2 FILLER_111_643 ();
 FILLCELL_X1 FILLER_111_645 ();
 FILLCELL_X4 FILLER_111_665 ();
 FILLCELL_X1 FILLER_111_692 ();
 FILLCELL_X4 FILLER_111_712 ();
 FILLCELL_X2 FILLER_111_719 ();
 FILLCELL_X8 FILLER_111_755 ();
 FILLCELL_X1 FILLER_111_763 ();
 FILLCELL_X4 FILLER_111_774 ();
 FILLCELL_X2 FILLER_111_778 ();
 FILLCELL_X8 FILLER_111_783 ();
 FILLCELL_X2 FILLER_111_821 ();
 FILLCELL_X2 FILLER_111_825 ();
 FILLCELL_X8 FILLER_111_843 ();
 FILLCELL_X2 FILLER_111_851 ();
 FILLCELL_X16 FILLER_111_855 ();
 FILLCELL_X1 FILLER_111_871 ();
 FILLCELL_X32 FILLER_111_892 ();
 FILLCELL_X16 FILLER_111_924 ();
 FILLCELL_X8 FILLER_111_940 ();
 FILLCELL_X2 FILLER_111_948 ();
 FILLCELL_X1 FILLER_111_950 ();
 FILLCELL_X4 FILLER_111_977 ();
 FILLCELL_X1 FILLER_111_981 ();
 FILLCELL_X2 FILLER_112_1 ();
 FILLCELL_X8 FILLER_112_6 ();
 FILLCELL_X1 FILLER_112_14 ();
 FILLCELL_X16 FILLER_112_49 ();
 FILLCELL_X8 FILLER_112_65 ();
 FILLCELL_X4 FILLER_112_73 ();
 FILLCELL_X1 FILLER_112_77 ();
 FILLCELL_X32 FILLER_112_95 ();
 FILLCELL_X16 FILLER_112_127 ();
 FILLCELL_X2 FILLER_112_143 ();
 FILLCELL_X1 FILLER_112_145 ();
 FILLCELL_X8 FILLER_112_169 ();
 FILLCELL_X1 FILLER_112_177 ();
 FILLCELL_X4 FILLER_112_181 ();
 FILLCELL_X1 FILLER_112_185 ();
 FILLCELL_X1 FILLER_112_203 ();
 FILLCELL_X32 FILLER_112_215 ();
 FILLCELL_X32 FILLER_112_247 ();
 FILLCELL_X8 FILLER_112_279 ();
 FILLCELL_X4 FILLER_112_287 ();
 FILLCELL_X4 FILLER_112_303 ();
 FILLCELL_X1 FILLER_112_307 ();
 FILLCELL_X1 FILLER_112_313 ();
 FILLCELL_X8 FILLER_112_328 ();
 FILLCELL_X2 FILLER_112_336 ();
 FILLCELL_X8 FILLER_112_357 ();
 FILLCELL_X4 FILLER_112_365 ();
 FILLCELL_X2 FILLER_112_369 ();
 FILLCELL_X1 FILLER_112_383 ();
 FILLCELL_X2 FILLER_112_414 ();
 FILLCELL_X8 FILLER_112_427 ();
 FILLCELL_X4 FILLER_112_435 ();
 FILLCELL_X2 FILLER_112_439 ();
 FILLCELL_X1 FILLER_112_441 ();
 FILLCELL_X1 FILLER_112_455 ();
 FILLCELL_X2 FILLER_112_505 ();
 FILLCELL_X1 FILLER_112_507 ();
 FILLCELL_X2 FILLER_112_519 ();
 FILLCELL_X8 FILLER_112_530 ();
 FILLCELL_X2 FILLER_112_538 ();
 FILLCELL_X1 FILLER_112_540 ();
 FILLCELL_X2 FILLER_112_615 ();
 FILLCELL_X2 FILLER_112_628 ();
 FILLCELL_X1 FILLER_112_630 ();
 FILLCELL_X4 FILLER_112_632 ();
 FILLCELL_X2 FILLER_112_636 ();
 FILLCELL_X16 FILLER_112_657 ();
 FILLCELL_X2 FILLER_112_690 ();
 FILLCELL_X1 FILLER_112_692 ();
 FILLCELL_X2 FILLER_112_700 ();
 FILLCELL_X1 FILLER_112_702 ();
 FILLCELL_X8 FILLER_112_715 ();
 FILLCELL_X2 FILLER_112_723 ();
 FILLCELL_X1 FILLER_112_725 ();
 FILLCELL_X2 FILLER_112_729 ();
 FILLCELL_X2 FILLER_112_734 ();
 FILLCELL_X1 FILLER_112_736 ();
 FILLCELL_X8 FILLER_112_743 ();
 FILLCELL_X2 FILLER_112_751 ();
 FILLCELL_X4 FILLER_112_756 ();
 FILLCELL_X8 FILLER_112_767 ();
 FILLCELL_X2 FILLER_112_777 ();
 FILLCELL_X1 FILLER_112_779 ();
 FILLCELL_X4 FILLER_112_783 ();
 FILLCELL_X2 FILLER_112_787 ();
 FILLCELL_X4 FILLER_112_796 ();
 FILLCELL_X1 FILLER_112_800 ();
 FILLCELL_X4 FILLER_112_811 ();
 FILLCELL_X8 FILLER_112_819 ();
 FILLCELL_X2 FILLER_112_827 ();
 FILLCELL_X1 FILLER_112_829 ();
 FILLCELL_X2 FILLER_112_849 ();
 FILLCELL_X1 FILLER_112_851 ();
 FILLCELL_X16 FILLER_112_873 ();
 FILLCELL_X2 FILLER_112_889 ();
 FILLCELL_X1 FILLER_112_891 ();
 FILLCELL_X1 FILLER_112_904 ();
 FILLCELL_X8 FILLER_112_915 ();
 FILLCELL_X1 FILLER_112_923 ();
 FILLCELL_X16 FILLER_112_938 ();
 FILLCELL_X16 FILLER_112_956 ();
 FILLCELL_X8 FILLER_112_972 ();
 FILLCELL_X2 FILLER_112_980 ();
 FILLCELL_X8 FILLER_113_1 ();
 FILLCELL_X4 FILLER_113_9 ();
 FILLCELL_X2 FILLER_113_13 ();
 FILLCELL_X1 FILLER_113_15 ();
 FILLCELL_X8 FILLER_113_19 ();
 FILLCELL_X16 FILLER_113_30 ();
 FILLCELL_X4 FILLER_113_46 ();
 FILLCELL_X2 FILLER_113_50 ();
 FILLCELL_X1 FILLER_113_52 ();
 FILLCELL_X4 FILLER_113_61 ();
 FILLCELL_X8 FILLER_113_68 ();
 FILLCELL_X32 FILLER_113_113 ();
 FILLCELL_X1 FILLER_113_145 ();
 FILLCELL_X8 FILLER_113_169 ();
 FILLCELL_X1 FILLER_113_177 ();
 FILLCELL_X2 FILLER_113_198 ();
 FILLCELL_X1 FILLER_113_200 ();
 FILLCELL_X4 FILLER_113_229 ();
 FILLCELL_X2 FILLER_113_240 ();
 FILLCELL_X1 FILLER_113_264 ();
 FILLCELL_X1 FILLER_113_276 ();
 FILLCELL_X2 FILLER_113_284 ();
 FILLCELL_X1 FILLER_113_286 ();
 FILLCELL_X4 FILLER_113_291 ();
 FILLCELL_X2 FILLER_113_295 ();
 FILLCELL_X4 FILLER_113_306 ();
 FILLCELL_X16 FILLER_113_340 ();
 FILLCELL_X8 FILLER_113_356 ();
 FILLCELL_X4 FILLER_113_364 ();
 FILLCELL_X2 FILLER_113_368 ();
 FILLCELL_X1 FILLER_113_407 ();
 FILLCELL_X8 FILLER_113_430 ();
 FILLCELL_X2 FILLER_113_438 ();
 FILLCELL_X4 FILLER_113_458 ();
 FILLCELL_X1 FILLER_113_462 ();
 FILLCELL_X8 FILLER_113_488 ();
 FILLCELL_X2 FILLER_113_527 ();
 FILLCELL_X1 FILLER_113_529 ();
 FILLCELL_X2 FILLER_113_567 ();
 FILLCELL_X4 FILLER_113_614 ();
 FILLCELL_X16 FILLER_113_661 ();
 FILLCELL_X8 FILLER_113_677 ();
 FILLCELL_X2 FILLER_113_685 ();
 FILLCELL_X1 FILLER_113_687 ();
 FILLCELL_X8 FILLER_113_705 ();
 FILLCELL_X4 FILLER_113_713 ();
 FILLCELL_X1 FILLER_113_717 ();
 FILLCELL_X1 FILLER_113_722 ();
 FILLCELL_X2 FILLER_113_726 ();
 FILLCELL_X1 FILLER_113_728 ();
 FILLCELL_X4 FILLER_113_758 ();
 FILLCELL_X1 FILLER_113_762 ();
 FILLCELL_X32 FILLER_113_773 ();
 FILLCELL_X4 FILLER_113_805 ();
 FILLCELL_X1 FILLER_113_809 ();
 FILLCELL_X2 FILLER_113_831 ();
 FILLCELL_X4 FILLER_113_853 ();
 FILLCELL_X32 FILLER_113_859 ();
 FILLCELL_X2 FILLER_113_891 ();
 FILLCELL_X4 FILLER_113_895 ();
 FILLCELL_X1 FILLER_113_899 ();
 FILLCELL_X8 FILLER_113_910 ();
 FILLCELL_X1 FILLER_113_944 ();
 FILLCELL_X16 FILLER_113_963 ();
 FILLCELL_X2 FILLER_113_979 ();
 FILLCELL_X1 FILLER_113_981 ();
 FILLCELL_X1 FILLER_114_1 ();
 FILLCELL_X2 FILLER_114_19 ();
 FILLCELL_X1 FILLER_114_28 ();
 FILLCELL_X4 FILLER_114_32 ();
 FILLCELL_X4 FILLER_114_39 ();
 FILLCELL_X2 FILLER_114_64 ();
 FILLCELL_X1 FILLER_114_66 ();
 FILLCELL_X8 FILLER_114_70 ();
 FILLCELL_X1 FILLER_114_78 ();
 FILLCELL_X16 FILLER_114_99 ();
 FILLCELL_X4 FILLER_114_115 ();
 FILLCELL_X2 FILLER_114_119 ();
 FILLCELL_X1 FILLER_114_121 ();
 FILLCELL_X2 FILLER_114_151 ();
 FILLCELL_X1 FILLER_114_162 ();
 FILLCELL_X2 FILLER_114_183 ();
 FILLCELL_X1 FILLER_114_185 ();
 FILLCELL_X8 FILLER_114_189 ();
 FILLCELL_X1 FILLER_114_197 ();
 FILLCELL_X8 FILLER_114_229 ();
 FILLCELL_X4 FILLER_114_259 ();
 FILLCELL_X1 FILLER_114_263 ();
 FILLCELL_X16 FILLER_114_306 ();
 FILLCELL_X1 FILLER_114_322 ();
 FILLCELL_X8 FILLER_114_349 ();
 FILLCELL_X4 FILLER_114_357 ();
 FILLCELL_X2 FILLER_114_361 ();
 FILLCELL_X2 FILLER_114_388 ();
 FILLCELL_X4 FILLER_114_418 ();
 FILLCELL_X4 FILLER_114_427 ();
 FILLCELL_X4 FILLER_114_450 ();
 FILLCELL_X2 FILLER_114_467 ();
 FILLCELL_X4 FILLER_114_486 ();
 FILLCELL_X4 FILLER_114_519 ();
 FILLCELL_X2 FILLER_114_523 ();
 FILLCELL_X1 FILLER_114_525 ();
 FILLCELL_X1 FILLER_114_551 ();
 FILLCELL_X2 FILLER_114_569 ();
 FILLCELL_X1 FILLER_114_571 ();
 FILLCELL_X1 FILLER_114_611 ();
 FILLCELL_X4 FILLER_114_632 ();
 FILLCELL_X1 FILLER_114_636 ();
 FILLCELL_X1 FILLER_114_643 ();
 FILLCELL_X1 FILLER_114_647 ();
 FILLCELL_X32 FILLER_114_651 ();
 FILLCELL_X32 FILLER_114_683 ();
 FILLCELL_X16 FILLER_114_749 ();
 FILLCELL_X4 FILLER_114_765 ();
 FILLCELL_X2 FILLER_114_769 ();
 FILLCELL_X8 FILLER_114_774 ();
 FILLCELL_X1 FILLER_114_782 ();
 FILLCELL_X4 FILLER_114_786 ();
 FILLCELL_X2 FILLER_114_790 ();
 FILLCELL_X1 FILLER_114_795 ();
 FILLCELL_X32 FILLER_114_799 ();
 FILLCELL_X4 FILLER_114_831 ();
 FILLCELL_X8 FILLER_114_853 ();
 FILLCELL_X1 FILLER_114_861 ();
 FILLCELL_X16 FILLER_114_878 ();
 FILLCELL_X8 FILLER_114_896 ();
 FILLCELL_X8 FILLER_114_914 ();
 FILLCELL_X4 FILLER_114_922 ();
 FILLCELL_X1 FILLER_114_926 ();
 FILLCELL_X1 FILLER_114_943 ();
 FILLCELL_X2 FILLER_114_946 ();
 FILLCELL_X1 FILLER_114_948 ();
 FILLCELL_X8 FILLER_114_951 ();
 FILLCELL_X2 FILLER_114_959 ();
 FILLCELL_X1 FILLER_114_961 ();
 FILLCELL_X4 FILLER_114_978 ();
 FILLCELL_X8 FILLER_115_1 ();
 FILLCELL_X1 FILLER_115_9 ();
 FILLCELL_X8 FILLER_115_13 ();
 FILLCELL_X16 FILLER_115_42 ();
 FILLCELL_X8 FILLER_115_58 ();
 FILLCELL_X8 FILLER_115_73 ();
 FILLCELL_X4 FILLER_115_81 ();
 FILLCELL_X1 FILLER_115_85 ();
 FILLCELL_X8 FILLER_115_95 ();
 FILLCELL_X4 FILLER_115_103 ();
 FILLCELL_X2 FILLER_115_107 ();
 FILLCELL_X1 FILLER_115_109 ();
 FILLCELL_X4 FILLER_115_130 ();
 FILLCELL_X1 FILLER_115_134 ();
 FILLCELL_X2 FILLER_115_141 ();
 FILLCELL_X1 FILLER_115_143 ();
 FILLCELL_X16 FILLER_115_147 ();
 FILLCELL_X8 FILLER_115_163 ();
 FILLCELL_X4 FILLER_115_171 ();
 FILLCELL_X2 FILLER_115_175 ();
 FILLCELL_X1 FILLER_115_177 ();
 FILLCELL_X32 FILLER_115_184 ();
 FILLCELL_X1 FILLER_115_216 ();
 FILLCELL_X4 FILLER_115_239 ();
 FILLCELL_X4 FILLER_115_245 ();
 FILLCELL_X2 FILLER_115_249 ();
 FILLCELL_X32 FILLER_115_260 ();
 FILLCELL_X4 FILLER_115_292 ();
 FILLCELL_X1 FILLER_115_296 ();
 FILLCELL_X16 FILLER_115_314 ();
 FILLCELL_X4 FILLER_115_330 ();
 FILLCELL_X16 FILLER_115_351 ();
 FILLCELL_X8 FILLER_115_367 ();
 FILLCELL_X2 FILLER_115_400 ();
 FILLCELL_X2 FILLER_115_425 ();
 FILLCELL_X8 FILLER_115_444 ();
 FILLCELL_X1 FILLER_115_474 ();
 FILLCELL_X4 FILLER_115_534 ();
 FILLCELL_X2 FILLER_115_538 ();
 FILLCELL_X1 FILLER_115_560 ();
 FILLCELL_X1 FILLER_115_588 ();
 FILLCELL_X8 FILLER_115_600 ();
 FILLCELL_X4 FILLER_115_645 ();
 FILLCELL_X1 FILLER_115_649 ();
 FILLCELL_X8 FILLER_115_654 ();
 FILLCELL_X2 FILLER_115_669 ();
 FILLCELL_X1 FILLER_115_671 ();
 FILLCELL_X8 FILLER_115_675 ();
 FILLCELL_X4 FILLER_115_687 ();
 FILLCELL_X2 FILLER_115_691 ();
 FILLCELL_X4 FILLER_115_696 ();
 FILLCELL_X16 FILLER_115_704 ();
 FILLCELL_X8 FILLER_115_720 ();
 FILLCELL_X4 FILLER_115_728 ();
 FILLCELL_X2 FILLER_115_732 ();
 FILLCELL_X16 FILLER_115_737 ();
 FILLCELL_X4 FILLER_115_753 ();
 FILLCELL_X2 FILLER_115_757 ();
 FILLCELL_X1 FILLER_115_775 ();
 FILLCELL_X16 FILLER_115_792 ();
 FILLCELL_X4 FILLER_115_808 ();
 FILLCELL_X1 FILLER_115_812 ();
 FILLCELL_X4 FILLER_115_871 ();
 FILLCELL_X1 FILLER_115_875 ();
 FILLCELL_X4 FILLER_115_894 ();
 FILLCELL_X8 FILLER_115_914 ();
 FILLCELL_X2 FILLER_115_922 ();
 FILLCELL_X1 FILLER_115_924 ();
 FILLCELL_X4 FILLER_115_927 ();
 FILLCELL_X2 FILLER_115_931 ();
 FILLCELL_X1 FILLER_115_933 ();
 FILLCELL_X8 FILLER_115_944 ();
 FILLCELL_X2 FILLER_115_952 ();
 FILLCELL_X1 FILLER_115_970 ();
 FILLCELL_X8 FILLER_115_973 ();
 FILLCELL_X1 FILLER_115_981 ();
 FILLCELL_X32 FILLER_116_1 ();
 FILLCELL_X16 FILLER_116_33 ();
 FILLCELL_X8 FILLER_116_49 ();
 FILLCELL_X4 FILLER_116_57 ();
 FILLCELL_X2 FILLER_116_61 ();
 FILLCELL_X4 FILLER_116_66 ();
 FILLCELL_X1 FILLER_116_73 ();
 FILLCELL_X8 FILLER_116_77 ();
 FILLCELL_X1 FILLER_116_85 ();
 FILLCELL_X16 FILLER_116_97 ();
 FILLCELL_X8 FILLER_116_113 ();
 FILLCELL_X4 FILLER_116_121 ();
 FILLCELL_X2 FILLER_116_131 ();
 FILLCELL_X16 FILLER_116_159 ();
 FILLCELL_X4 FILLER_116_175 ();
 FILLCELL_X1 FILLER_116_179 ();
 FILLCELL_X8 FILLER_116_197 ();
 FILLCELL_X4 FILLER_116_205 ();
 FILLCELL_X8 FILLER_116_216 ();
 FILLCELL_X2 FILLER_116_224 ();
 FILLCELL_X1 FILLER_116_226 ();
 FILLCELL_X16 FILLER_116_230 ();
 FILLCELL_X2 FILLER_116_246 ();
 FILLCELL_X16 FILLER_116_257 ();
 FILLCELL_X1 FILLER_116_273 ();
 FILLCELL_X32 FILLER_116_296 ();
 FILLCELL_X1 FILLER_116_328 ();
 FILLCELL_X4 FILLER_116_368 ();
 FILLCELL_X2 FILLER_116_372 ();
 FILLCELL_X1 FILLER_116_374 ();
 FILLCELL_X16 FILLER_116_380 ();
 FILLCELL_X8 FILLER_116_396 ();
 FILLCELL_X1 FILLER_116_404 ();
 FILLCELL_X8 FILLER_116_419 ();
 FILLCELL_X4 FILLER_116_427 ();
 FILLCELL_X2 FILLER_116_431 ();
 FILLCELL_X1 FILLER_116_433 ();
 FILLCELL_X8 FILLER_116_452 ();
 FILLCELL_X4 FILLER_116_460 ();
 FILLCELL_X1 FILLER_116_500 ();
 FILLCELL_X1 FILLER_116_557 ();
 FILLCELL_X4 FILLER_116_586 ();
 FILLCELL_X1 FILLER_116_590 ();
 FILLCELL_X8 FILLER_116_622 ();
 FILLCELL_X1 FILLER_116_630 ();
 FILLCELL_X4 FILLER_116_632 ();
 FILLCELL_X1 FILLER_116_636 ();
 FILLCELL_X2 FILLER_116_644 ();
 FILLCELL_X1 FILLER_116_646 ();
 FILLCELL_X8 FILLER_116_719 ();
 FILLCELL_X4 FILLER_116_727 ();
 FILLCELL_X1 FILLER_116_738 ();
 FILLCELL_X16 FILLER_116_756 ();
 FILLCELL_X1 FILLER_116_772 ();
 FILLCELL_X4 FILLER_116_775 ();
 FILLCELL_X2 FILLER_116_779 ();
 FILLCELL_X16 FILLER_116_797 ();
 FILLCELL_X4 FILLER_116_813 ();
 FILLCELL_X16 FILLER_116_820 ();
 FILLCELL_X8 FILLER_116_836 ();
 FILLCELL_X1 FILLER_116_844 ();
 FILLCELL_X1 FILLER_116_847 ();
 FILLCELL_X16 FILLER_116_868 ();
 FILLCELL_X4 FILLER_116_887 ();
 FILLCELL_X1 FILLER_116_896 ();
 FILLCELL_X4 FILLER_116_909 ();
 FILLCELL_X1 FILLER_116_913 ();
 FILLCELL_X16 FILLER_116_916 ();
 FILLCELL_X2 FILLER_116_932 ();
 FILLCELL_X2 FILLER_116_956 ();
 FILLCELL_X4 FILLER_116_960 ();
 FILLCELL_X2 FILLER_116_980 ();
 FILLCELL_X16 FILLER_117_1 ();
 FILLCELL_X8 FILLER_117_17 ();
 FILLCELL_X4 FILLER_117_25 ();
 FILLCELL_X2 FILLER_117_29 ();
 FILLCELL_X8 FILLER_117_34 ();
 FILLCELL_X4 FILLER_117_42 ();
 FILLCELL_X2 FILLER_117_46 ();
 FILLCELL_X2 FILLER_117_74 ();
 FILLCELL_X2 FILLER_117_130 ();
 FILLCELL_X16 FILLER_117_195 ();
 FILLCELL_X4 FILLER_117_218 ();
 FILLCELL_X2 FILLER_117_222 ();
 FILLCELL_X1 FILLER_117_224 ();
 FILLCELL_X4 FILLER_117_231 ();
 FILLCELL_X2 FILLER_117_235 ();
 FILLCELL_X1 FILLER_117_237 ();
 FILLCELL_X8 FILLER_117_258 ();
 FILLCELL_X4 FILLER_117_266 ();
 FILLCELL_X1 FILLER_117_270 ();
 FILLCELL_X16 FILLER_117_303 ();
 FILLCELL_X4 FILLER_117_319 ();
 FILLCELL_X1 FILLER_117_323 ();
 FILLCELL_X4 FILLER_117_343 ();
 FILLCELL_X2 FILLER_117_347 ();
 FILLCELL_X2 FILLER_117_354 ();
 FILLCELL_X8 FILLER_117_361 ();
 FILLCELL_X2 FILLER_117_400 ();
 FILLCELL_X1 FILLER_117_402 ();
 FILLCELL_X2 FILLER_117_434 ();
 FILLCELL_X1 FILLER_117_436 ();
 FILLCELL_X2 FILLER_117_457 ();
 FILLCELL_X2 FILLER_117_464 ();
 FILLCELL_X1 FILLER_117_466 ();
 FILLCELL_X2 FILLER_117_484 ();
 FILLCELL_X4 FILLER_117_512 ();
 FILLCELL_X2 FILLER_117_516 ();
 FILLCELL_X1 FILLER_117_518 ();
 FILLCELL_X8 FILLER_117_544 ();
 FILLCELL_X1 FILLER_117_552 ();
 FILLCELL_X16 FILLER_117_570 ();
 FILLCELL_X8 FILLER_117_586 ();
 FILLCELL_X1 FILLER_117_594 ();
 FILLCELL_X16 FILLER_117_604 ();
 FILLCELL_X4 FILLER_117_620 ();
 FILLCELL_X2 FILLER_117_624 ();
 FILLCELL_X32 FILLER_117_643 ();
 FILLCELL_X2 FILLER_117_675 ();
 FILLCELL_X1 FILLER_117_677 ();
 FILLCELL_X4 FILLER_117_705 ();
 FILLCELL_X1 FILLER_117_709 ();
 FILLCELL_X32 FILLER_117_730 ();
 FILLCELL_X8 FILLER_117_762 ();
 FILLCELL_X16 FILLER_117_780 ();
 FILLCELL_X1 FILLER_117_796 ();
 FILLCELL_X2 FILLER_117_799 ();
 FILLCELL_X16 FILLER_117_803 ();
 FILLCELL_X8 FILLER_117_819 ();
 FILLCELL_X4 FILLER_117_827 ();
 FILLCELL_X4 FILLER_117_833 ();
 FILLCELL_X2 FILLER_117_837 ();
 FILLCELL_X2 FILLER_117_867 ();
 FILLCELL_X8 FILLER_117_871 ();
 FILLCELL_X8 FILLER_117_889 ();
 FILLCELL_X4 FILLER_117_897 ();
 FILLCELL_X1 FILLER_117_911 ();
 FILLCELL_X4 FILLER_117_922 ();
 FILLCELL_X2 FILLER_117_928 ();
 FILLCELL_X32 FILLER_117_940 ();
 FILLCELL_X8 FILLER_117_972 ();
 FILLCELL_X2 FILLER_117_980 ();
 FILLCELL_X16 FILLER_118_1 ();
 FILLCELL_X4 FILLER_118_17 ();
 FILLCELL_X1 FILLER_118_21 ();
 FILLCELL_X16 FILLER_118_25 ();
 FILLCELL_X2 FILLER_118_41 ();
 FILLCELL_X1 FILLER_118_64 ();
 FILLCELL_X8 FILLER_118_68 ();
 FILLCELL_X2 FILLER_118_76 ();
 FILLCELL_X32 FILLER_118_89 ();
 FILLCELL_X1 FILLER_118_133 ();
 FILLCELL_X1 FILLER_118_140 ();
 FILLCELL_X4 FILLER_118_147 ();
 FILLCELL_X1 FILLER_118_151 ();
 FILLCELL_X4 FILLER_118_155 ();
 FILLCELL_X2 FILLER_118_159 ();
 FILLCELL_X1 FILLER_118_161 ();
 FILLCELL_X2 FILLER_118_168 ();
 FILLCELL_X16 FILLER_118_173 ();
 FILLCELL_X4 FILLER_118_189 ();
 FILLCELL_X1 FILLER_118_193 ();
 FILLCELL_X8 FILLER_118_200 ();
 FILLCELL_X1 FILLER_118_208 ();
 FILLCELL_X8 FILLER_118_212 ();
 FILLCELL_X1 FILLER_118_220 ();
 FILLCELL_X2 FILLER_118_244 ();
 FILLCELL_X2 FILLER_118_266 ();
 FILLCELL_X1 FILLER_118_268 ();
 FILLCELL_X2 FILLER_118_297 ();
 FILLCELL_X16 FILLER_118_316 ();
 FILLCELL_X8 FILLER_118_332 ();
 FILLCELL_X2 FILLER_118_340 ();
 FILLCELL_X1 FILLER_118_342 ();
 FILLCELL_X32 FILLER_118_350 ();
 FILLCELL_X4 FILLER_118_382 ();
 FILLCELL_X2 FILLER_118_386 ();
 FILLCELL_X1 FILLER_118_388 ();
 FILLCELL_X1 FILLER_118_406 ();
 FILLCELL_X1 FILLER_118_440 ();
 FILLCELL_X1 FILLER_118_452 ();
 FILLCELL_X2 FILLER_118_470 ();
 FILLCELL_X1 FILLER_118_472 ();
 FILLCELL_X16 FILLER_118_509 ();
 FILLCELL_X8 FILLER_118_525 ();
 FILLCELL_X1 FILLER_118_533 ();
 FILLCELL_X32 FILLER_118_539 ();
 FILLCELL_X32 FILLER_118_571 ();
 FILLCELL_X16 FILLER_118_603 ();
 FILLCELL_X8 FILLER_118_619 ();
 FILLCELL_X4 FILLER_118_627 ();
 FILLCELL_X2 FILLER_118_632 ();
 FILLCELL_X1 FILLER_118_634 ();
 FILLCELL_X8 FILLER_118_640 ();
 FILLCELL_X4 FILLER_118_648 ();
 FILLCELL_X1 FILLER_118_652 ();
 FILLCELL_X2 FILLER_118_657 ();
 FILLCELL_X2 FILLER_118_662 ();
 FILLCELL_X1 FILLER_118_664 ();
 FILLCELL_X16 FILLER_118_668 ();
 FILLCELL_X4 FILLER_118_684 ();
 FILLCELL_X4 FILLER_118_691 ();
 FILLCELL_X2 FILLER_118_695 ();
 FILLCELL_X8 FILLER_118_700 ();
 FILLCELL_X2 FILLER_118_708 ();
 FILLCELL_X4 FILLER_118_725 ();
 FILLCELL_X1 FILLER_118_729 ();
 FILLCELL_X8 FILLER_118_754 ();
 FILLCELL_X2 FILLER_118_762 ();
 FILLCELL_X2 FILLER_118_784 ();
 FILLCELL_X1 FILLER_118_786 ();
 FILLCELL_X16 FILLER_118_823 ();
 FILLCELL_X4 FILLER_118_839 ();
 FILLCELL_X2 FILLER_118_843 ();
 FILLCELL_X1 FILLER_118_845 ();
 FILLCELL_X8 FILLER_118_851 ();
 FILLCELL_X4 FILLER_118_859 ();
 FILLCELL_X2 FILLER_118_881 ();
 FILLCELL_X1 FILLER_118_883 ();
 FILLCELL_X2 FILLER_118_894 ();
 FILLCELL_X1 FILLER_118_898 ();
 FILLCELL_X2 FILLER_118_919 ();
 FILLCELL_X1 FILLER_118_939 ();
 FILLCELL_X1 FILLER_118_958 ();
 FILLCELL_X16 FILLER_118_961 ();
 FILLCELL_X4 FILLER_118_977 ();
 FILLCELL_X1 FILLER_118_981 ();
 FILLCELL_X32 FILLER_119_1 ();
 FILLCELL_X8 FILLER_119_33 ();
 FILLCELL_X4 FILLER_119_41 ();
 FILLCELL_X1 FILLER_119_45 ();
 FILLCELL_X8 FILLER_119_51 ();
 FILLCELL_X8 FILLER_119_62 ();
 FILLCELL_X4 FILLER_119_70 ();
 FILLCELL_X2 FILLER_119_74 ();
 FILLCELL_X1 FILLER_119_76 ();
 FILLCELL_X16 FILLER_119_96 ();
 FILLCELL_X2 FILLER_119_112 ();
 FILLCELL_X8 FILLER_119_148 ();
 FILLCELL_X1 FILLER_119_156 ();
 FILLCELL_X32 FILLER_119_212 ();
 FILLCELL_X1 FILLER_119_244 ();
 FILLCELL_X16 FILLER_119_253 ();
 FILLCELL_X2 FILLER_119_269 ();
 FILLCELL_X4 FILLER_119_288 ();
 FILLCELL_X1 FILLER_119_292 ();
 FILLCELL_X1 FILLER_119_310 ();
 FILLCELL_X8 FILLER_119_341 ();
 FILLCELL_X2 FILLER_119_349 ();
 FILLCELL_X1 FILLER_119_351 ();
 FILLCELL_X8 FILLER_119_377 ();
 FILLCELL_X2 FILLER_119_385 ();
 FILLCELL_X2 FILLER_119_404 ();
 FILLCELL_X4 FILLER_119_417 ();
 FILLCELL_X2 FILLER_119_421 ();
 FILLCELL_X16 FILLER_119_458 ();
 FILLCELL_X8 FILLER_119_474 ();
 FILLCELL_X4 FILLER_119_482 ();
 FILLCELL_X8 FILLER_119_503 ();
 FILLCELL_X4 FILLER_119_511 ();
 FILLCELL_X1 FILLER_119_518 ();
 FILLCELL_X2 FILLER_119_522 ();
 FILLCELL_X1 FILLER_119_524 ();
 FILLCELL_X4 FILLER_119_529 ();
 FILLCELL_X1 FILLER_119_533 ();
 FILLCELL_X4 FILLER_119_537 ();
 FILLCELL_X1 FILLER_119_555 ();
 FILLCELL_X4 FILLER_119_560 ();
 FILLCELL_X1 FILLER_119_567 ();
 FILLCELL_X8 FILLER_119_575 ();
 FILLCELL_X4 FILLER_119_583 ();
 FILLCELL_X1 FILLER_119_587 ();
 FILLCELL_X8 FILLER_119_591 ();
 FILLCELL_X1 FILLER_119_599 ();
 FILLCELL_X1 FILLER_119_606 ();
 FILLCELL_X8 FILLER_119_624 ();
 FILLCELL_X4 FILLER_119_632 ();
 FILLCELL_X2 FILLER_119_636 ();
 FILLCELL_X1 FILLER_119_644 ();
 FILLCELL_X4 FILLER_119_667 ();
 FILLCELL_X2 FILLER_119_671 ();
 FILLCELL_X1 FILLER_119_673 ();
 FILLCELL_X4 FILLER_119_678 ();
 FILLCELL_X2 FILLER_119_682 ();
 FILLCELL_X1 FILLER_119_684 ();
 FILLCELL_X2 FILLER_119_707 ();
 FILLCELL_X1 FILLER_119_709 ();
 FILLCELL_X32 FILLER_119_727 ();
 FILLCELL_X4 FILLER_119_759 ();
 FILLCELL_X1 FILLER_119_763 ();
 FILLCELL_X4 FILLER_119_780 ();
 FILLCELL_X1 FILLER_119_784 ();
 FILLCELL_X8 FILLER_119_797 ();
 FILLCELL_X2 FILLER_119_807 ();
 FILLCELL_X8 FILLER_119_825 ();
 FILLCELL_X4 FILLER_119_833 ();
 FILLCELL_X32 FILLER_119_847 ();
 FILLCELL_X8 FILLER_119_879 ();
 FILLCELL_X4 FILLER_119_887 ();
 FILLCELL_X1 FILLER_119_891 ();
 FILLCELL_X1 FILLER_119_894 ();
 FILLCELL_X8 FILLER_119_897 ();
 FILLCELL_X2 FILLER_119_905 ();
 FILLCELL_X1 FILLER_119_907 ();
 FILLCELL_X16 FILLER_119_910 ();
 FILLCELL_X8 FILLER_119_926 ();
 FILLCELL_X1 FILLER_119_934 ();
 FILLCELL_X1 FILLER_119_939 ();
 FILLCELL_X4 FILLER_119_970 ();
 FILLCELL_X2 FILLER_119_974 ();
 FILLCELL_X4 FILLER_119_978 ();
 FILLCELL_X32 FILLER_120_1 ();
 FILLCELL_X16 FILLER_120_33 ();
 FILLCELL_X8 FILLER_120_49 ();
 FILLCELL_X1 FILLER_120_57 ();
 FILLCELL_X8 FILLER_120_65 ();
 FILLCELL_X4 FILLER_120_73 ();
 FILLCELL_X32 FILLER_120_84 ();
 FILLCELL_X4 FILLER_120_116 ();
 FILLCELL_X2 FILLER_120_137 ();
 FILLCELL_X8 FILLER_120_156 ();
 FILLCELL_X1 FILLER_120_164 ();
 FILLCELL_X8 FILLER_120_182 ();
 FILLCELL_X4 FILLER_120_190 ();
 FILLCELL_X1 FILLER_120_194 ();
 FILLCELL_X4 FILLER_120_198 ();
 FILLCELL_X1 FILLER_120_202 ();
 FILLCELL_X16 FILLER_120_210 ();
 FILLCELL_X8 FILLER_120_226 ();
 FILLCELL_X2 FILLER_120_234 ();
 FILLCELL_X8 FILLER_120_258 ();
 FILLCELL_X2 FILLER_120_266 ();
 FILLCELL_X8 FILLER_120_271 ();
 FILLCELL_X2 FILLER_120_279 ();
 FILLCELL_X8 FILLER_120_284 ();
 FILLCELL_X4 FILLER_120_292 ();
 FILLCELL_X1 FILLER_120_296 ();
 FILLCELL_X8 FILLER_120_300 ();
 FILLCELL_X1 FILLER_120_308 ();
 FILLCELL_X32 FILLER_120_312 ();
 FILLCELL_X16 FILLER_120_344 ();
 FILLCELL_X4 FILLER_120_385 ();
 FILLCELL_X2 FILLER_120_389 ();
 FILLCELL_X8 FILLER_120_434 ();
 FILLCELL_X2 FILLER_120_442 ();
 FILLCELL_X1 FILLER_120_444 ();
 FILLCELL_X32 FILLER_120_467 ();
 FILLCELL_X16 FILLER_120_499 ();
 FILLCELL_X1 FILLER_120_515 ();
 FILLCELL_X1 FILLER_120_533 ();
 FILLCELL_X1 FILLER_120_571 ();
 FILLCELL_X4 FILLER_120_596 ();
 FILLCELL_X1 FILLER_120_600 ();
 FILLCELL_X1 FILLER_120_608 ();
 FILLCELL_X4 FILLER_120_616 ();
 FILLCELL_X2 FILLER_120_620 ();
 FILLCELL_X1 FILLER_120_622 ();
 FILLCELL_X2 FILLER_120_628 ();
 FILLCELL_X1 FILLER_120_630 ();
 FILLCELL_X4 FILLER_120_632 ();
 FILLCELL_X1 FILLER_120_636 ();
 FILLCELL_X2 FILLER_120_659 ();
 FILLCELL_X1 FILLER_120_661 ();
 FILLCELL_X8 FILLER_120_669 ();
 FILLCELL_X4 FILLER_120_677 ();
 FILLCELL_X2 FILLER_120_681 ();
 FILLCELL_X32 FILLER_120_700 ();
 FILLCELL_X2 FILLER_120_732 ();
 FILLCELL_X1 FILLER_120_734 ();
 FILLCELL_X8 FILLER_120_756 ();
 FILLCELL_X4 FILLER_120_764 ();
 FILLCELL_X2 FILLER_120_768 ();
 FILLCELL_X1 FILLER_120_770 ();
 FILLCELL_X16 FILLER_120_773 ();
 FILLCELL_X2 FILLER_120_789 ();
 FILLCELL_X1 FILLER_120_791 ();
 FILLCELL_X16 FILLER_120_794 ();
 FILLCELL_X8 FILLER_120_810 ();
 FILLCELL_X4 FILLER_120_818 ();
 FILLCELL_X2 FILLER_120_822 ();
 FILLCELL_X4 FILLER_120_834 ();
 FILLCELL_X1 FILLER_120_838 ();
 FILLCELL_X8 FILLER_120_854 ();
 FILLCELL_X2 FILLER_120_862 ();
 FILLCELL_X8 FILLER_120_880 ();
 FILLCELL_X1 FILLER_120_888 ();
 FILLCELL_X1 FILLER_120_899 ();
 FILLCELL_X8 FILLER_120_914 ();
 FILLCELL_X1 FILLER_120_922 ();
 FILLCELL_X4 FILLER_120_925 ();
 FILLCELL_X1 FILLER_120_929 ();
 FILLCELL_X2 FILLER_120_940 ();
 FILLCELL_X1 FILLER_120_942 ();
 FILLCELL_X4 FILLER_120_975 ();
 FILLCELL_X2 FILLER_120_979 ();
 FILLCELL_X1 FILLER_120_981 ();
 FILLCELL_X32 FILLER_121_1 ();
 FILLCELL_X8 FILLER_121_33 ();
 FILLCELL_X4 FILLER_121_41 ();
 FILLCELL_X1 FILLER_121_45 ();
 FILLCELL_X2 FILLER_121_80 ();
 FILLCELL_X8 FILLER_121_87 ();
 FILLCELL_X4 FILLER_121_95 ();
 FILLCELL_X1 FILLER_121_99 ();
 FILLCELL_X32 FILLER_121_102 ();
 FILLCELL_X32 FILLER_121_134 ();
 FILLCELL_X32 FILLER_121_166 ();
 FILLCELL_X4 FILLER_121_215 ();
 FILLCELL_X2 FILLER_121_219 ();
 FILLCELL_X1 FILLER_121_221 ();
 FILLCELL_X4 FILLER_121_231 ();
 FILLCELL_X2 FILLER_121_235 ();
 FILLCELL_X8 FILLER_121_256 ();
 FILLCELL_X4 FILLER_121_264 ();
 FILLCELL_X16 FILLER_121_271 ();
 FILLCELL_X8 FILLER_121_287 ();
 FILLCELL_X4 FILLER_121_299 ();
 FILLCELL_X1 FILLER_121_303 ();
 FILLCELL_X32 FILLER_121_312 ();
 FILLCELL_X32 FILLER_121_344 ();
 FILLCELL_X4 FILLER_121_376 ();
 FILLCELL_X1 FILLER_121_414 ();
 FILLCELL_X8 FILLER_121_424 ();
 FILLCELL_X2 FILLER_121_432 ();
 FILLCELL_X4 FILLER_121_456 ();
 FILLCELL_X1 FILLER_121_460 ();
 FILLCELL_X8 FILLER_121_464 ();
 FILLCELL_X4 FILLER_121_472 ();
 FILLCELL_X1 FILLER_121_476 ();
 FILLCELL_X4 FILLER_121_480 ();
 FILLCELL_X1 FILLER_121_484 ();
 FILLCELL_X4 FILLER_121_489 ();
 FILLCELL_X8 FILLER_121_496 ();
 FILLCELL_X4 FILLER_121_504 ();
 FILLCELL_X4 FILLER_121_515 ();
 FILLCELL_X8 FILLER_121_522 ();
 FILLCELL_X4 FILLER_121_530 ();
 FILLCELL_X2 FILLER_121_534 ();
 FILLCELL_X8 FILLER_121_540 ();
 FILLCELL_X8 FILLER_121_551 ();
 FILLCELL_X8 FILLER_121_562 ();
 FILLCELL_X1 FILLER_121_591 ();
 FILLCELL_X2 FILLER_121_595 ();
 FILLCELL_X16 FILLER_121_614 ();
 FILLCELL_X8 FILLER_121_630 ();
 FILLCELL_X2 FILLER_121_638 ();
 FILLCELL_X1 FILLER_121_640 ();
 FILLCELL_X2 FILLER_121_658 ();
 FILLCELL_X2 FILLER_121_677 ();
 FILLCELL_X1 FILLER_121_679 ();
 FILLCELL_X8 FILLER_121_691 ();
 FILLCELL_X1 FILLER_121_699 ();
 FILLCELL_X2 FILLER_121_705 ();
 FILLCELL_X2 FILLER_121_732 ();
 FILLCELL_X4 FILLER_121_738 ();
 FILLCELL_X16 FILLER_121_748 ();
 FILLCELL_X8 FILLER_121_764 ();
 FILLCELL_X4 FILLER_121_772 ();
 FILLCELL_X2 FILLER_121_776 ();
 FILLCELL_X4 FILLER_121_794 ();
 FILLCELL_X2 FILLER_121_798 ();
 FILLCELL_X1 FILLER_121_800 ();
 FILLCELL_X4 FILLER_121_815 ();
 FILLCELL_X1 FILLER_121_831 ();
 FILLCELL_X8 FILLER_121_834 ();
 FILLCELL_X2 FILLER_121_842 ();
 FILLCELL_X1 FILLER_121_844 ();
 FILLCELL_X16 FILLER_121_855 ();
 FILLCELL_X4 FILLER_121_871 ();
 FILLCELL_X1 FILLER_121_875 ();
 FILLCELL_X2 FILLER_121_880 ();
 FILLCELL_X1 FILLER_121_882 ();
 FILLCELL_X16 FILLER_121_885 ();
 FILLCELL_X8 FILLER_121_901 ();
 FILLCELL_X1 FILLER_121_909 ();
 FILLCELL_X8 FILLER_121_920 ();
 FILLCELL_X4 FILLER_121_928 ();
 FILLCELL_X2 FILLER_121_932 ();
 FILLCELL_X8 FILLER_121_938 ();
 FILLCELL_X4 FILLER_121_946 ();
 FILLCELL_X2 FILLER_121_950 ();
 FILLCELL_X1 FILLER_121_952 ();
 FILLCELL_X16 FILLER_121_955 ();
 FILLCELL_X8 FILLER_121_971 ();
 FILLCELL_X2 FILLER_121_979 ();
 FILLCELL_X1 FILLER_121_981 ();
 FILLCELL_X32 FILLER_122_1 ();
 FILLCELL_X32 FILLER_122_33 ();
 FILLCELL_X16 FILLER_122_65 ();
 FILLCELL_X4 FILLER_122_81 ();
 FILLCELL_X2 FILLER_122_85 ();
 FILLCELL_X32 FILLER_122_118 ();
 FILLCELL_X4 FILLER_122_150 ();
 FILLCELL_X16 FILLER_122_160 ();
 FILLCELL_X2 FILLER_122_176 ();
 FILLCELL_X1 FILLER_122_178 ();
 FILLCELL_X8 FILLER_122_187 ();
 FILLCELL_X2 FILLER_122_195 ();
 FILLCELL_X4 FILLER_122_200 ();
 FILLCELL_X2 FILLER_122_204 ();
 FILLCELL_X4 FILLER_122_209 ();
 FILLCELL_X2 FILLER_122_213 ();
 FILLCELL_X1 FILLER_122_215 ();
 FILLCELL_X16 FILLER_122_239 ();
 FILLCELL_X2 FILLER_122_259 ();
 FILLCELL_X1 FILLER_122_261 ();
 FILLCELL_X4 FILLER_122_265 ();
 FILLCELL_X2 FILLER_122_269 ();
 FILLCELL_X1 FILLER_122_271 ();
 FILLCELL_X8 FILLER_122_276 ();
 FILLCELL_X4 FILLER_122_284 ();
 FILLCELL_X2 FILLER_122_291 ();
 FILLCELL_X1 FILLER_122_293 ();
 FILLCELL_X8 FILLER_122_301 ();
 FILLCELL_X8 FILLER_122_313 ();
 FILLCELL_X2 FILLER_122_321 ();
 FILLCELL_X2 FILLER_122_326 ();
 FILLCELL_X1 FILLER_122_336 ();
 FILLCELL_X2 FILLER_122_340 ();
 FILLCELL_X16 FILLER_122_345 ();
 FILLCELL_X4 FILLER_122_361 ();
 FILLCELL_X1 FILLER_122_365 ();
 FILLCELL_X16 FILLER_122_373 ();
 FILLCELL_X8 FILLER_122_389 ();
 FILLCELL_X4 FILLER_122_397 ();
 FILLCELL_X1 FILLER_122_401 ();
 FILLCELL_X4 FILLER_122_405 ();
 FILLCELL_X2 FILLER_122_409 ();
 FILLCELL_X4 FILLER_122_428 ();
 FILLCELL_X2 FILLER_122_432 ();
 FILLCELL_X2 FILLER_122_451 ();
 FILLCELL_X16 FILLER_122_456 ();
 FILLCELL_X2 FILLER_122_472 ();
 FILLCELL_X1 FILLER_122_481 ();
 FILLCELL_X1 FILLER_122_499 ();
 FILLCELL_X2 FILLER_122_517 ();
 FILLCELL_X8 FILLER_122_523 ();
 FILLCELL_X2 FILLER_122_531 ();
 FILLCELL_X1 FILLER_122_533 ();
 FILLCELL_X1 FILLER_122_539 ();
 FILLCELL_X2 FILLER_122_543 ();
 FILLCELL_X1 FILLER_122_545 ();
 FILLCELL_X2 FILLER_122_550 ();
 FILLCELL_X1 FILLER_122_552 ();
 FILLCELL_X8 FILLER_122_556 ();
 FILLCELL_X2 FILLER_122_564 ();
 FILLCELL_X2 FILLER_122_571 ();
 FILLCELL_X32 FILLER_122_587 ();
 FILLCELL_X8 FILLER_122_619 ();
 FILLCELL_X4 FILLER_122_627 ();
 FILLCELL_X1 FILLER_122_632 ();
 FILLCELL_X8 FILLER_122_650 ();
 FILLCELL_X4 FILLER_122_658 ();
 FILLCELL_X2 FILLER_122_662 ();
 FILLCELL_X1 FILLER_122_664 ();
 FILLCELL_X4 FILLER_122_670 ();
 FILLCELL_X2 FILLER_122_674 ();
 FILLCELL_X4 FILLER_122_716 ();
 FILLCELL_X2 FILLER_122_720 ();
 FILLCELL_X1 FILLER_122_722 ();
 FILLCELL_X4 FILLER_122_726 ();
 FILLCELL_X2 FILLER_122_730 ();
 FILLCELL_X1 FILLER_122_732 ();
 FILLCELL_X2 FILLER_122_750 ();
 FILLCELL_X16 FILLER_122_755 ();
 FILLCELL_X8 FILLER_122_798 ();
 FILLCELL_X4 FILLER_122_806 ();
 FILLCELL_X2 FILLER_122_810 ();
 FILLCELL_X2 FILLER_122_828 ();
 FILLCELL_X1 FILLER_122_830 ();
 FILLCELL_X4 FILLER_122_841 ();
 FILLCELL_X1 FILLER_122_845 ();
 FILLCELL_X4 FILLER_122_886 ();
 FILLCELL_X2 FILLER_122_906 ();
 FILLCELL_X8 FILLER_122_910 ();
 FILLCELL_X4 FILLER_122_918 ();
 FILLCELL_X4 FILLER_122_932 ();
 FILLCELL_X32 FILLER_122_946 ();
 FILLCELL_X4 FILLER_122_978 ();
 FILLCELL_X32 FILLER_123_1 ();
 FILLCELL_X32 FILLER_123_33 ();
 FILLCELL_X16 FILLER_123_65 ();
 FILLCELL_X4 FILLER_123_81 ();
 FILLCELL_X1 FILLER_123_85 ();
 FILLCELL_X2 FILLER_123_90 ();
 FILLCELL_X1 FILLER_123_92 ();
 FILLCELL_X8 FILLER_123_96 ();
 FILLCELL_X2 FILLER_123_104 ();
 FILLCELL_X1 FILLER_123_106 ();
 FILLCELL_X2 FILLER_123_110 ();
 FILLCELL_X1 FILLER_123_112 ();
 FILLCELL_X8 FILLER_123_120 ();
 FILLCELL_X2 FILLER_123_128 ();
 FILLCELL_X1 FILLER_123_130 ();
 FILLCELL_X2 FILLER_123_137 ();
 FILLCELL_X1 FILLER_123_139 ();
 FILLCELL_X8 FILLER_123_144 ();
 FILLCELL_X4 FILLER_123_152 ();
 FILLCELL_X2 FILLER_123_156 ();
 FILLCELL_X1 FILLER_123_161 ();
 FILLCELL_X8 FILLER_123_165 ();
 FILLCELL_X4 FILLER_123_173 ();
 FILLCELL_X1 FILLER_123_177 ();
 FILLCELL_X4 FILLER_123_181 ();
 FILLCELL_X1 FILLER_123_205 ();
 FILLCELL_X8 FILLER_123_210 ();
 FILLCELL_X4 FILLER_123_218 ();
 FILLCELL_X2 FILLER_123_222 ();
 FILLCELL_X16 FILLER_123_227 ();
 FILLCELL_X4 FILLER_123_263 ();
 FILLCELL_X1 FILLER_123_267 ();
 FILLCELL_X1 FILLER_123_288 ();
 FILLCELL_X2 FILLER_123_323 ();
 FILLCELL_X8 FILLER_123_349 ();
 FILLCELL_X4 FILLER_123_357 ();
 FILLCELL_X16 FILLER_123_378 ();
 FILLCELL_X4 FILLER_123_394 ();
 FILLCELL_X2 FILLER_123_398 ();
 FILLCELL_X1 FILLER_123_400 ();
 FILLCELL_X4 FILLER_123_407 ();
 FILLCELL_X2 FILLER_123_411 ();
 FILLCELL_X4 FILLER_123_421 ();
 FILLCELL_X2 FILLER_123_425 ();
 FILLCELL_X1 FILLER_123_427 ();
 FILLCELL_X16 FILLER_123_445 ();
 FILLCELL_X1 FILLER_123_465 ();
 FILLCELL_X1 FILLER_123_469 ();
 FILLCELL_X8 FILLER_123_487 ();
 FILLCELL_X1 FILLER_123_495 ();
 FILLCELL_X4 FILLER_123_499 ();
 FILLCELL_X2 FILLER_123_535 ();
 FILLCELL_X1 FILLER_123_542 ();
 FILLCELL_X32 FILLER_123_563 ();
 FILLCELL_X4 FILLER_123_595 ();
 FILLCELL_X2 FILLER_123_599 ();
 FILLCELL_X2 FILLER_123_608 ();
 FILLCELL_X1 FILLER_123_610 ();
 FILLCELL_X2 FILLER_123_614 ();
 FILLCELL_X2 FILLER_123_627 ();
 FILLCELL_X2 FILLER_123_632 ();
 FILLCELL_X8 FILLER_123_637 ();
 FILLCELL_X4 FILLER_123_645 ();
 FILLCELL_X1 FILLER_123_656 ();
 FILLCELL_X1 FILLER_123_667 ();
 FILLCELL_X8 FILLER_123_671 ();
 FILLCELL_X4 FILLER_123_679 ();
 FILLCELL_X1 FILLER_123_683 ();
 FILLCELL_X4 FILLER_123_692 ();
 FILLCELL_X2 FILLER_123_696 ();
 FILLCELL_X4 FILLER_123_702 ();
 FILLCELL_X16 FILLER_123_709 ();
 FILLCELL_X4 FILLER_123_725 ();
 FILLCELL_X2 FILLER_123_729 ();
 FILLCELL_X2 FILLER_123_735 ();
 FILLCELL_X16 FILLER_123_769 ();
 FILLCELL_X4 FILLER_123_795 ();
 FILLCELL_X16 FILLER_123_829 ();
 FILLCELL_X1 FILLER_123_845 ();
 FILLCELL_X2 FILLER_123_850 ();
 FILLCELL_X16 FILLER_123_854 ();
 FILLCELL_X2 FILLER_123_870 ();
 FILLCELL_X1 FILLER_123_872 ();
 FILLCELL_X8 FILLER_123_883 ();
 FILLCELL_X4 FILLER_123_891 ();
 FILLCELL_X2 FILLER_123_895 ();
 FILLCELL_X2 FILLER_123_899 ();
 FILLCELL_X1 FILLER_123_917 ();
 FILLCELL_X32 FILLER_123_950 ();
 FILLCELL_X32 FILLER_124_1 ();
 FILLCELL_X32 FILLER_124_33 ();
 FILLCELL_X8 FILLER_124_65 ();
 FILLCELL_X4 FILLER_124_73 ();
 FILLCELL_X2 FILLER_124_77 ();
 FILLCELL_X2 FILLER_124_96 ();
 FILLCELL_X2 FILLER_124_127 ();
 FILLCELL_X1 FILLER_124_129 ();
 FILLCELL_X1 FILLER_124_133 ();
 FILLCELL_X2 FILLER_124_141 ();
 FILLCELL_X1 FILLER_124_143 ();
 FILLCELL_X1 FILLER_124_165 ();
 FILLCELL_X8 FILLER_124_169 ();
 FILLCELL_X8 FILLER_124_184 ();
 FILLCELL_X4 FILLER_124_192 ();
 FILLCELL_X4 FILLER_124_200 ();
 FILLCELL_X8 FILLER_124_207 ();
 FILLCELL_X4 FILLER_124_215 ();
 FILLCELL_X16 FILLER_124_226 ();
 FILLCELL_X4 FILLER_124_242 ();
 FILLCELL_X2 FILLER_124_246 ();
 FILLCELL_X2 FILLER_124_251 ();
 FILLCELL_X1 FILLER_124_253 ();
 FILLCELL_X32 FILLER_124_257 ();
 FILLCELL_X4 FILLER_124_289 ();
 FILLCELL_X1 FILLER_124_293 ();
 FILLCELL_X2 FILLER_124_298 ();
 FILLCELL_X2 FILLER_124_303 ();
 FILLCELL_X1 FILLER_124_305 ();
 FILLCELL_X4 FILLER_124_309 ();
 FILLCELL_X4 FILLER_124_321 ();
 FILLCELL_X8 FILLER_124_334 ();
 FILLCELL_X32 FILLER_124_346 ();
 FILLCELL_X16 FILLER_124_378 ();
 FILLCELL_X2 FILLER_124_394 ();
 FILLCELL_X1 FILLER_124_396 ();
 FILLCELL_X2 FILLER_124_400 ();
 FILLCELL_X1 FILLER_124_402 ();
 FILLCELL_X32 FILLER_124_406 ();
 FILLCELL_X16 FILLER_124_438 ();
 FILLCELL_X4 FILLER_124_471 ();
 FILLCELL_X2 FILLER_124_475 ();
 FILLCELL_X1 FILLER_124_477 ();
 FILLCELL_X16 FILLER_124_481 ();
 FILLCELL_X2 FILLER_124_497 ();
 FILLCELL_X8 FILLER_124_502 ();
 FILLCELL_X4 FILLER_124_510 ();
 FILLCELL_X2 FILLER_124_514 ();
 FILLCELL_X2 FILLER_124_519 ();
 FILLCELL_X16 FILLER_124_524 ();
 FILLCELL_X4 FILLER_124_540 ();
 FILLCELL_X8 FILLER_124_547 ();
 FILLCELL_X1 FILLER_124_555 ();
 FILLCELL_X8 FILLER_124_563 ();
 FILLCELL_X2 FILLER_124_571 ();
 FILLCELL_X4 FILLER_124_577 ();
 FILLCELL_X1 FILLER_124_581 ();
 FILLCELL_X8 FILLER_124_586 ();
 FILLCELL_X2 FILLER_124_594 ();
 FILLCELL_X1 FILLER_124_596 ();
 FILLCELL_X8 FILLER_124_635 ();
 FILLCELL_X2 FILLER_124_643 ();
 FILLCELL_X1 FILLER_124_645 ();
 FILLCELL_X8 FILLER_124_669 ();
 FILLCELL_X4 FILLER_124_682 ();
 FILLCELL_X2 FILLER_124_686 ();
 FILLCELL_X1 FILLER_124_688 ();
 FILLCELL_X16 FILLER_124_711 ();
 FILLCELL_X2 FILLER_124_727 ();
 FILLCELL_X1 FILLER_124_729 ();
 FILLCELL_X32 FILLER_124_747 ();
 FILLCELL_X2 FILLER_124_779 ();
 FILLCELL_X8 FILLER_124_783 ();
 FILLCELL_X4 FILLER_124_791 ();
 FILLCELL_X2 FILLER_124_795 ();
 FILLCELL_X16 FILLER_124_801 ();
 FILLCELL_X4 FILLER_124_817 ();
 FILLCELL_X2 FILLER_124_821 ();
 FILLCELL_X2 FILLER_124_825 ();
 FILLCELL_X8 FILLER_124_829 ();
 FILLCELL_X4 FILLER_124_837 ();
 FILLCELL_X8 FILLER_124_857 ();
 FILLCELL_X1 FILLER_124_865 ();
 FILLCELL_X2 FILLER_124_896 ();
 FILLCELL_X16 FILLER_124_908 ();
 FILLCELL_X8 FILLER_124_924 ();
 FILLCELL_X4 FILLER_124_932 ();
 FILLCELL_X32 FILLER_124_938 ();
 FILLCELL_X8 FILLER_124_970 ();
 FILLCELL_X4 FILLER_124_978 ();
 FILLCELL_X32 FILLER_125_1 ();
 FILLCELL_X32 FILLER_125_33 ();
 FILLCELL_X16 FILLER_125_65 ();
 FILLCELL_X8 FILLER_125_81 ();
 FILLCELL_X4 FILLER_125_89 ();
 FILLCELL_X2 FILLER_125_93 ();
 FILLCELL_X8 FILLER_125_112 ();
 FILLCELL_X2 FILLER_125_120 ();
 FILLCELL_X1 FILLER_125_122 ();
 FILLCELL_X4 FILLER_125_140 ();
 FILLCELL_X1 FILLER_125_144 ();
 FILLCELL_X1 FILLER_125_152 ();
 FILLCELL_X1 FILLER_125_170 ();
 FILLCELL_X1 FILLER_125_188 ();
 FILLCELL_X1 FILLER_125_206 ();
 FILLCELL_X2 FILLER_125_231 ();
 FILLCELL_X1 FILLER_125_233 ();
 FILLCELL_X8 FILLER_125_251 ();
 FILLCELL_X16 FILLER_125_266 ();
 FILLCELL_X2 FILLER_125_282 ();
 FILLCELL_X1 FILLER_125_284 ();
 FILLCELL_X4 FILLER_125_330 ();
 FILLCELL_X2 FILLER_125_334 ();
 FILLCELL_X1 FILLER_125_336 ();
 FILLCELL_X16 FILLER_125_354 ();
 FILLCELL_X8 FILLER_125_370 ();
 FILLCELL_X4 FILLER_125_378 ();
 FILLCELL_X1 FILLER_125_382 ();
 FILLCELL_X8 FILLER_125_390 ();
 FILLCELL_X4 FILLER_125_398 ();
 FILLCELL_X16 FILLER_125_406 ();
 FILLCELL_X8 FILLER_125_422 ();
 FILLCELL_X2 FILLER_125_430 ();
 FILLCELL_X4 FILLER_125_435 ();
 FILLCELL_X2 FILLER_125_439 ();
 FILLCELL_X1 FILLER_125_441 ();
 FILLCELL_X8 FILLER_125_445 ();
 FILLCELL_X16 FILLER_125_460 ();
 FILLCELL_X8 FILLER_125_476 ();
 FILLCELL_X4 FILLER_125_484 ();
 FILLCELL_X1 FILLER_125_488 ();
 FILLCELL_X4 FILLER_125_493 ();
 FILLCELL_X1 FILLER_125_497 ();
 FILLCELL_X4 FILLER_125_502 ();
 FILLCELL_X2 FILLER_125_506 ();
 FILLCELL_X4 FILLER_125_511 ();
 FILLCELL_X1 FILLER_125_515 ();
 FILLCELL_X4 FILLER_125_520 ();
 FILLCELL_X4 FILLER_125_527 ();
 FILLCELL_X2 FILLER_125_531 ();
 FILLCELL_X1 FILLER_125_533 ();
 FILLCELL_X1 FILLER_125_539 ();
 FILLCELL_X2 FILLER_125_562 ();
 FILLCELL_X1 FILLER_125_564 ();
 FILLCELL_X4 FILLER_125_599 ();
 FILLCELL_X1 FILLER_125_612 ();
 FILLCELL_X8 FILLER_125_616 ();
 FILLCELL_X1 FILLER_125_632 ();
 FILLCELL_X16 FILLER_125_636 ();
 FILLCELL_X32 FILLER_125_671 ();
 FILLCELL_X8 FILLER_125_703 ();
 FILLCELL_X1 FILLER_125_711 ();
 FILLCELL_X8 FILLER_125_719 ();
 FILLCELL_X16 FILLER_125_731 ();
 FILLCELL_X4 FILLER_125_747 ();
 FILLCELL_X1 FILLER_125_751 ();
 FILLCELL_X8 FILLER_125_773 ();
 FILLCELL_X2 FILLER_125_781 ();
 FILLCELL_X1 FILLER_125_783 ();
 FILLCELL_X8 FILLER_125_800 ();
 FILLCELL_X2 FILLER_125_812 ();
 FILLCELL_X1 FILLER_125_814 ();
 FILLCELL_X1 FILLER_125_817 ();
 FILLCELL_X4 FILLER_125_834 ();
 FILLCELL_X16 FILLER_125_840 ();
 FILLCELL_X8 FILLER_125_856 ();
 FILLCELL_X2 FILLER_125_864 ();
 FILLCELL_X1 FILLER_125_866 ();
 FILLCELL_X8 FILLER_125_869 ();
 FILLCELL_X2 FILLER_125_877 ();
 FILLCELL_X4 FILLER_125_895 ();
 FILLCELL_X1 FILLER_125_899 ();
 FILLCELL_X2 FILLER_125_916 ();
 FILLCELL_X1 FILLER_125_928 ();
 FILLCELL_X2 FILLER_125_931 ();
 FILLCELL_X32 FILLER_125_937 ();
 FILLCELL_X8 FILLER_125_969 ();
 FILLCELL_X4 FILLER_125_977 ();
 FILLCELL_X1 FILLER_125_981 ();
 FILLCELL_X32 FILLER_126_1 ();
 FILLCELL_X32 FILLER_126_33 ();
 FILLCELL_X32 FILLER_126_65 ();
 FILLCELL_X32 FILLER_126_97 ();
 FILLCELL_X16 FILLER_126_129 ();
 FILLCELL_X2 FILLER_126_145 ();
 FILLCELL_X1 FILLER_126_147 ();
 FILLCELL_X4 FILLER_126_156 ();
 FILLCELL_X2 FILLER_126_160 ();
 FILLCELL_X32 FILLER_126_165 ();
 FILLCELL_X16 FILLER_126_197 ();
 FILLCELL_X2 FILLER_126_213 ();
 FILLCELL_X4 FILLER_126_232 ();
 FILLCELL_X2 FILLER_126_236 ();
 FILLCELL_X2 FILLER_126_245 ();
 FILLCELL_X4 FILLER_126_251 ();
 FILLCELL_X2 FILLER_126_255 ();
 FILLCELL_X1 FILLER_126_257 ();
 FILLCELL_X4 FILLER_126_275 ();
 FILLCELL_X2 FILLER_126_279 ();
 FILLCELL_X2 FILLER_126_285 ();
 FILLCELL_X4 FILLER_126_297 ();
 FILLCELL_X2 FILLER_126_301 ();
 FILLCELL_X1 FILLER_126_303 ();
 FILLCELL_X4 FILLER_126_312 ();
 FILLCELL_X8 FILLER_126_321 ();
 FILLCELL_X2 FILLER_126_329 ();
 FILLCELL_X1 FILLER_126_331 ();
 FILLCELL_X1 FILLER_126_342 ();
 FILLCELL_X4 FILLER_126_360 ();
 FILLCELL_X2 FILLER_126_381 ();
 FILLCELL_X1 FILLER_126_383 ();
 FILLCELL_X8 FILLER_126_408 ();
 FILLCELL_X1 FILLER_126_416 ();
 FILLCELL_X8 FILLER_126_438 ();
 FILLCELL_X2 FILLER_126_446 ();
 FILLCELL_X4 FILLER_126_468 ();
 FILLCELL_X2 FILLER_126_472 ();
 FILLCELL_X2 FILLER_126_491 ();
 FILLCELL_X2 FILLER_126_510 ();
 FILLCELL_X1 FILLER_126_512 ();
 FILLCELL_X2 FILLER_126_530 ();
 FILLCELL_X1 FILLER_126_532 ();
 FILLCELL_X2 FILLER_126_537 ();
 FILLCELL_X1 FILLER_126_539 ();
 FILLCELL_X1 FILLER_126_544 ();
 FILLCELL_X16 FILLER_126_548 ();
 FILLCELL_X1 FILLER_126_564 ();
 FILLCELL_X1 FILLER_126_568 ();
 FILLCELL_X16 FILLER_126_587 ();
 FILLCELL_X4 FILLER_126_603 ();
 FILLCELL_X1 FILLER_126_607 ();
 FILLCELL_X16 FILLER_126_612 ();
 FILLCELL_X2 FILLER_126_628 ();
 FILLCELL_X1 FILLER_126_630 ();
 FILLCELL_X16 FILLER_126_632 ();
 FILLCELL_X4 FILLER_126_648 ();
 FILLCELL_X2 FILLER_126_652 ();
 FILLCELL_X4 FILLER_126_658 ();
 FILLCELL_X8 FILLER_126_682 ();
 FILLCELL_X4 FILLER_126_694 ();
 FILLCELL_X2 FILLER_126_701 ();
 FILLCELL_X1 FILLER_126_707 ();
 FILLCELL_X4 FILLER_126_745 ();
 FILLCELL_X1 FILLER_126_749 ();
 FILLCELL_X4 FILLER_126_777 ();
 FILLCELL_X2 FILLER_126_781 ();
 FILLCELL_X1 FILLER_126_783 ();
 FILLCELL_X4 FILLER_126_794 ();
 FILLCELL_X1 FILLER_126_798 ();
 FILLCELL_X8 FILLER_126_825 ();
 FILLCELL_X2 FILLER_126_833 ();
 FILLCELL_X1 FILLER_126_835 ();
 FILLCELL_X2 FILLER_126_878 ();
 FILLCELL_X2 FILLER_126_892 ();
 FILLCELL_X32 FILLER_126_918 ();
 FILLCELL_X32 FILLER_126_950 ();
 FILLCELL_X32 FILLER_127_1 ();
 FILLCELL_X32 FILLER_127_33 ();
 FILLCELL_X32 FILLER_127_65 ();
 FILLCELL_X16 FILLER_127_97 ();
 FILLCELL_X8 FILLER_127_137 ();
 FILLCELL_X4 FILLER_127_145 ();
 FILLCELL_X1 FILLER_127_149 ();
 FILLCELL_X16 FILLER_127_157 ();
 FILLCELL_X4 FILLER_127_173 ();
 FILLCELL_X2 FILLER_127_177 ();
 FILLCELL_X8 FILLER_127_186 ();
 FILLCELL_X2 FILLER_127_194 ();
 FILLCELL_X16 FILLER_127_199 ();
 FILLCELL_X16 FILLER_127_249 ();
 FILLCELL_X2 FILLER_127_265 ();
 FILLCELL_X1 FILLER_127_267 ();
 FILLCELL_X1 FILLER_127_275 ();
 FILLCELL_X2 FILLER_127_314 ();
 FILLCELL_X8 FILLER_127_319 ();
 FILLCELL_X2 FILLER_127_327 ();
 FILLCELL_X1 FILLER_127_329 ();
 FILLCELL_X16 FILLER_127_335 ();
 FILLCELL_X8 FILLER_127_351 ();
 FILLCELL_X4 FILLER_127_359 ();
 FILLCELL_X1 FILLER_127_363 ();
 FILLCELL_X8 FILLER_127_392 ();
 FILLCELL_X2 FILLER_127_400 ();
 FILLCELL_X1 FILLER_127_402 ();
 FILLCELL_X8 FILLER_127_410 ();
 FILLCELL_X4 FILLER_127_418 ();
 FILLCELL_X2 FILLER_127_422 ();
 FILLCELL_X1 FILLER_127_424 ();
 FILLCELL_X8 FILLER_127_446 ();
 FILLCELL_X4 FILLER_127_454 ();
 FILLCELL_X8 FILLER_127_462 ();
 FILLCELL_X4 FILLER_127_470 ();
 FILLCELL_X1 FILLER_127_474 ();
 FILLCELL_X2 FILLER_127_489 ();
 FILLCELL_X16 FILLER_127_494 ();
 FILLCELL_X1 FILLER_127_510 ();
 FILLCELL_X4 FILLER_127_514 ();
 FILLCELL_X8 FILLER_127_522 ();
 FILLCELL_X4 FILLER_127_530 ();
 FILLCELL_X2 FILLER_127_534 ();
 FILLCELL_X4 FILLER_127_553 ();
 FILLCELL_X1 FILLER_127_557 ();
 FILLCELL_X4 FILLER_127_561 ();
 FILLCELL_X1 FILLER_127_565 ();
 FILLCELL_X2 FILLER_127_574 ();
 FILLCELL_X8 FILLER_127_593 ();
 FILLCELL_X4 FILLER_127_601 ();
 FILLCELL_X1 FILLER_127_605 ();
 FILLCELL_X2 FILLER_127_623 ();
 FILLCELL_X16 FILLER_127_629 ();
 FILLCELL_X1 FILLER_127_662 ();
 FILLCELL_X8 FILLER_127_670 ();
 FILLCELL_X4 FILLER_127_678 ();
 FILLCELL_X1 FILLER_127_682 ();
 FILLCELL_X16 FILLER_127_720 ();
 FILLCELL_X8 FILLER_127_736 ();
 FILLCELL_X4 FILLER_127_744 ();
 FILLCELL_X2 FILLER_127_748 ();
 FILLCELL_X1 FILLER_127_750 ();
 FILLCELL_X2 FILLER_127_755 ();
 FILLCELL_X16 FILLER_127_760 ();
 FILLCELL_X8 FILLER_127_776 ();
 FILLCELL_X2 FILLER_127_784 ();
 FILLCELL_X4 FILLER_127_796 ();
 FILLCELL_X2 FILLER_127_800 ();
 FILLCELL_X1 FILLER_127_802 ();
 FILLCELL_X8 FILLER_127_819 ();
 FILLCELL_X4 FILLER_127_827 ();
 FILLCELL_X2 FILLER_127_831 ();
 FILLCELL_X1 FILLER_127_867 ();
 FILLCELL_X2 FILLER_127_870 ();
 FILLCELL_X1 FILLER_127_872 ();
 FILLCELL_X8 FILLER_127_889 ();
 FILLCELL_X1 FILLER_127_899 ();
 FILLCELL_X32 FILLER_127_910 ();
 FILLCELL_X32 FILLER_127_942 ();
 FILLCELL_X8 FILLER_127_974 ();
 FILLCELL_X32 FILLER_128_1 ();
 FILLCELL_X32 FILLER_128_33 ();
 FILLCELL_X32 FILLER_128_65 ();
 FILLCELL_X32 FILLER_128_97 ();
 FILLCELL_X1 FILLER_128_133 ();
 FILLCELL_X1 FILLER_128_145 ();
 FILLCELL_X8 FILLER_128_166 ();
 FILLCELL_X2 FILLER_128_174 ();
 FILLCELL_X2 FILLER_128_200 ();
 FILLCELL_X1 FILLER_128_202 ();
 FILLCELL_X2 FILLER_128_224 ();
 FILLCELL_X8 FILLER_128_229 ();
 FILLCELL_X1 FILLER_128_237 ();
 FILLCELL_X4 FILLER_128_241 ();
 FILLCELL_X2 FILLER_128_245 ();
 FILLCELL_X1 FILLER_128_247 ();
 FILLCELL_X4 FILLER_128_256 ();
 FILLCELL_X2 FILLER_128_260 ();
 FILLCELL_X1 FILLER_128_262 ();
 FILLCELL_X2 FILLER_128_280 ();
 FILLCELL_X1 FILLER_128_282 ();
 FILLCELL_X4 FILLER_128_286 ();
 FILLCELL_X1 FILLER_128_290 ();
 FILLCELL_X16 FILLER_128_308 ();
 FILLCELL_X8 FILLER_128_332 ();
 FILLCELL_X1 FILLER_128_340 ();
 FILLCELL_X32 FILLER_128_351 ();
 FILLCELL_X4 FILLER_128_383 ();
 FILLCELL_X8 FILLER_128_410 ();
 FILLCELL_X2 FILLER_128_418 ();
 FILLCELL_X4 FILLER_128_426 ();
 FILLCELL_X2 FILLER_128_430 ();
 FILLCELL_X1 FILLER_128_432 ();
 FILLCELL_X4 FILLER_128_436 ();
 FILLCELL_X1 FILLER_128_440 ();
 FILLCELL_X2 FILLER_128_444 ();
 FILLCELL_X1 FILLER_128_446 ();
 FILLCELL_X2 FILLER_128_450 ();
 FILLCELL_X4 FILLER_128_472 ();
 FILLCELL_X4 FILLER_128_479 ();
 FILLCELL_X2 FILLER_128_483 ();
 FILLCELL_X1 FILLER_128_489 ();
 FILLCELL_X8 FILLER_128_493 ();
 FILLCELL_X4 FILLER_128_501 ();
 FILLCELL_X2 FILLER_128_505 ();
 FILLCELL_X1 FILLER_128_507 ();
 FILLCELL_X1 FILLER_128_511 ();
 FILLCELL_X1 FILLER_128_532 ();
 FILLCELL_X8 FILLER_128_536 ();
 FILLCELL_X2 FILLER_128_544 ();
 FILLCELL_X1 FILLER_128_546 ();
 FILLCELL_X4 FILLER_128_550 ();
 FILLCELL_X1 FILLER_128_554 ();
 FILLCELL_X4 FILLER_128_560 ();
 FILLCELL_X1 FILLER_128_564 ();
 FILLCELL_X1 FILLER_128_570 ();
 FILLCELL_X1 FILLER_128_576 ();
 FILLCELL_X16 FILLER_128_580 ();
 FILLCELL_X2 FILLER_128_596 ();
 FILLCELL_X1 FILLER_128_598 ();
 FILLCELL_X4 FILLER_128_632 ();
 FILLCELL_X2 FILLER_128_636 ();
 FILLCELL_X4 FILLER_128_642 ();
 FILLCELL_X1 FILLER_128_646 ();
 FILLCELL_X4 FILLER_128_650 ();
 FILLCELL_X2 FILLER_128_654 ();
 FILLCELL_X1 FILLER_128_681 ();
 FILLCELL_X32 FILLER_128_692 ();
 FILLCELL_X2 FILLER_128_724 ();
 FILLCELL_X1 FILLER_128_726 ();
 FILLCELL_X4 FILLER_128_731 ();
 FILLCELL_X8 FILLER_128_738 ();
 FILLCELL_X2 FILLER_128_746 ();
 FILLCELL_X16 FILLER_128_765 ();
 FILLCELL_X8 FILLER_128_781 ();
 FILLCELL_X4 FILLER_128_789 ();
 FILLCELL_X1 FILLER_128_793 ();
 FILLCELL_X32 FILLER_128_804 ();
 FILLCELL_X8 FILLER_128_836 ();
 FILLCELL_X4 FILLER_128_844 ();
 FILLCELL_X2 FILLER_128_848 ();
 FILLCELL_X1 FILLER_128_852 ();
 FILLCELL_X1 FILLER_128_855 ();
 FILLCELL_X32 FILLER_128_866 ();
 FILLCELL_X32 FILLER_128_898 ();
 FILLCELL_X32 FILLER_128_930 ();
 FILLCELL_X16 FILLER_128_962 ();
 FILLCELL_X4 FILLER_128_978 ();
 FILLCELL_X32 FILLER_129_1 ();
 FILLCELL_X32 FILLER_129_33 ();
 FILLCELL_X32 FILLER_129_65 ();
 FILLCELL_X16 FILLER_129_97 ();
 FILLCELL_X4 FILLER_129_113 ();
 FILLCELL_X1 FILLER_129_117 ();
 FILLCELL_X16 FILLER_129_135 ();
 FILLCELL_X8 FILLER_129_157 ();
 FILLCELL_X2 FILLER_129_165 ();
 FILLCELL_X16 FILLER_129_198 ();
 FILLCELL_X1 FILLER_129_214 ();
 FILLCELL_X8 FILLER_129_225 ();
 FILLCELL_X4 FILLER_129_233 ();
 FILLCELL_X1 FILLER_129_237 ();
 FILLCELL_X16 FILLER_129_242 ();
 FILLCELL_X8 FILLER_129_258 ();
 FILLCELL_X2 FILLER_129_266 ();
 FILLCELL_X16 FILLER_129_271 ();
 FILLCELL_X4 FILLER_129_287 ();
 FILLCELL_X1 FILLER_129_291 ();
 FILLCELL_X4 FILLER_129_295 ();
 FILLCELL_X1 FILLER_129_299 ();
 FILLCELL_X4 FILLER_129_320 ();
 FILLCELL_X2 FILLER_129_341 ();
 FILLCELL_X1 FILLER_129_343 ();
 FILLCELL_X8 FILLER_129_356 ();
 FILLCELL_X4 FILLER_129_364 ();
 FILLCELL_X2 FILLER_129_368 ();
 FILLCELL_X32 FILLER_129_394 ();
 FILLCELL_X2 FILLER_129_426 ();
 FILLCELL_X1 FILLER_129_428 ();
 FILLCELL_X8 FILLER_129_432 ();
 FILLCELL_X4 FILLER_129_440 ();
 FILLCELL_X2 FILLER_129_444 ();
 FILLCELL_X1 FILLER_129_446 ();
 FILLCELL_X8 FILLER_129_451 ();
 FILLCELL_X1 FILLER_129_459 ();
 FILLCELL_X16 FILLER_129_463 ();
 FILLCELL_X2 FILLER_129_479 ();
 FILLCELL_X32 FILLER_129_498 ();
 FILLCELL_X2 FILLER_129_530 ();
 FILLCELL_X8 FILLER_129_539 ();
 FILLCELL_X4 FILLER_129_547 ();
 FILLCELL_X2 FILLER_129_551 ();
 FILLCELL_X8 FILLER_129_585 ();
 FILLCELL_X1 FILLER_129_593 ();
 FILLCELL_X8 FILLER_129_614 ();
 FILLCELL_X4 FILLER_129_622 ();
 FILLCELL_X2 FILLER_129_626 ();
 FILLCELL_X2 FILLER_129_631 ();
 FILLCELL_X1 FILLER_129_633 ();
 FILLCELL_X16 FILLER_129_651 ();
 FILLCELL_X4 FILLER_129_667 ();
 FILLCELL_X2 FILLER_129_671 ();
 FILLCELL_X1 FILLER_129_673 ();
 FILLCELL_X8 FILLER_129_679 ();
 FILLCELL_X4 FILLER_129_687 ();
 FILLCELL_X2 FILLER_129_695 ();
 FILLCELL_X1 FILLER_129_697 ();
 FILLCELL_X4 FILLER_129_703 ();
 FILLCELL_X4 FILLER_129_722 ();
 FILLCELL_X1 FILLER_129_726 ();
 FILLCELL_X2 FILLER_129_744 ();
 FILLCELL_X8 FILLER_129_750 ();
 FILLCELL_X2 FILLER_129_758 ();
 FILLCELL_X4 FILLER_129_763 ();
 FILLCELL_X2 FILLER_129_767 ();
 FILLCELL_X1 FILLER_129_769 ();
 FILLCELL_X32 FILLER_129_794 ();
 FILLCELL_X32 FILLER_129_826 ();
 FILLCELL_X32 FILLER_129_858 ();
 FILLCELL_X32 FILLER_129_890 ();
 FILLCELL_X32 FILLER_129_922 ();
 FILLCELL_X16 FILLER_129_954 ();
 FILLCELL_X8 FILLER_129_970 ();
 FILLCELL_X4 FILLER_129_978 ();
 FILLCELL_X32 FILLER_130_1 ();
 FILLCELL_X32 FILLER_130_33 ();
 FILLCELL_X32 FILLER_130_65 ();
 FILLCELL_X32 FILLER_130_97 ();
 FILLCELL_X4 FILLER_130_129 ();
 FILLCELL_X2 FILLER_130_133 ();
 FILLCELL_X1 FILLER_130_135 ();
 FILLCELL_X2 FILLER_130_160 ();
 FILLCELL_X4 FILLER_130_169 ();
 FILLCELL_X2 FILLER_130_173 ();
 FILLCELL_X2 FILLER_130_192 ();
 FILLCELL_X4 FILLER_130_205 ();
 FILLCELL_X4 FILLER_130_230 ();
 FILLCELL_X2 FILLER_130_234 ();
 FILLCELL_X2 FILLER_130_265 ();
 FILLCELL_X4 FILLER_130_271 ();
 FILLCELL_X2 FILLER_130_275 ();
 FILLCELL_X1 FILLER_130_277 ();
 FILLCELL_X4 FILLER_130_285 ();
 FILLCELL_X2 FILLER_130_289 ();
 FILLCELL_X1 FILLER_130_291 ();
 FILLCELL_X16 FILLER_130_296 ();
 FILLCELL_X4 FILLER_130_312 ();
 FILLCELL_X1 FILLER_130_316 ();
 FILLCELL_X4 FILLER_130_321 ();
 FILLCELL_X2 FILLER_130_325 ();
 FILLCELL_X1 FILLER_130_327 ();
 FILLCELL_X4 FILLER_130_332 ();
 FILLCELL_X2 FILLER_130_336 ();
 FILLCELL_X2 FILLER_130_344 ();
 FILLCELL_X4 FILLER_130_363 ();
 FILLCELL_X2 FILLER_130_367 ();
 FILLCELL_X1 FILLER_130_369 ();
 FILLCELL_X1 FILLER_130_394 ();
 FILLCELL_X1 FILLER_130_399 ();
 FILLCELL_X1 FILLER_130_417 ();
 FILLCELL_X1 FILLER_130_422 ();
 FILLCELL_X2 FILLER_130_427 ();
 FILLCELL_X1 FILLER_130_458 ();
 FILLCELL_X1 FILLER_130_463 ();
 FILLCELL_X4 FILLER_130_467 ();
 FILLCELL_X2 FILLER_130_471 ();
 FILLCELL_X1 FILLER_130_473 ();
 FILLCELL_X8 FILLER_130_478 ();
 FILLCELL_X4 FILLER_130_486 ();
 FILLCELL_X1 FILLER_130_490 ();
 FILLCELL_X2 FILLER_130_495 ();
 FILLCELL_X1 FILLER_130_497 ();
 FILLCELL_X4 FILLER_130_501 ();
 FILLCELL_X2 FILLER_130_505 ();
 FILLCELL_X1 FILLER_130_507 ();
 FILLCELL_X2 FILLER_130_532 ();
 FILLCELL_X1 FILLER_130_543 ();
 FILLCELL_X2 FILLER_130_548 ();
 FILLCELL_X1 FILLER_130_550 ();
 FILLCELL_X2 FILLER_130_554 ();
 FILLCELL_X1 FILLER_130_556 ();
 FILLCELL_X2 FILLER_130_561 ();
 FILLCELL_X4 FILLER_130_566 ();
 FILLCELL_X2 FILLER_130_570 ();
 FILLCELL_X16 FILLER_130_579 ();
 FILLCELL_X1 FILLER_130_595 ();
 FILLCELL_X8 FILLER_130_617 ();
 FILLCELL_X2 FILLER_130_629 ();
 FILLCELL_X2 FILLER_130_635 ();
 FILLCELL_X4 FILLER_130_641 ();
 FILLCELL_X1 FILLER_130_645 ();
 FILLCELL_X1 FILLER_130_654 ();
 FILLCELL_X4 FILLER_130_659 ();
 FILLCELL_X2 FILLER_130_663 ();
 FILLCELL_X2 FILLER_130_668 ();
 FILLCELL_X1 FILLER_130_670 ();
 FILLCELL_X4 FILLER_130_675 ();
 FILLCELL_X4 FILLER_130_682 ();
 FILLCELL_X1 FILLER_130_686 ();
 FILLCELL_X8 FILLER_130_727 ();
 FILLCELL_X4 FILLER_130_735 ();
 FILLCELL_X32 FILLER_130_793 ();
 FILLCELL_X32 FILLER_130_825 ();
 FILLCELL_X32 FILLER_130_857 ();
 FILLCELL_X32 FILLER_130_889 ();
 FILLCELL_X32 FILLER_130_921 ();
 FILLCELL_X16 FILLER_130_953 ();
 FILLCELL_X8 FILLER_130_969 ();
 FILLCELL_X4 FILLER_130_977 ();
 FILLCELL_X1 FILLER_130_981 ();
 FILLCELL_X32 FILLER_131_1 ();
 FILLCELL_X32 FILLER_131_33 ();
 FILLCELL_X32 FILLER_131_65 ();
 FILLCELL_X4 FILLER_131_97 ();
 FILLCELL_X2 FILLER_131_101 ();
 FILLCELL_X16 FILLER_131_106 ();
 FILLCELL_X8 FILLER_131_122 ();
 FILLCELL_X2 FILLER_131_130 ();
 FILLCELL_X1 FILLER_131_132 ();
 FILLCELL_X1 FILLER_131_157 ();
 FILLCELL_X8 FILLER_131_175 ();
 FILLCELL_X8 FILLER_131_203 ();
 FILLCELL_X4 FILLER_131_211 ();
 FILLCELL_X1 FILLER_131_235 ();
 FILLCELL_X1 FILLER_131_341 ();
 FILLCELL_X16 FILLER_131_345 ();
 FILLCELL_X8 FILLER_131_361 ();
 FILLCELL_X2 FILLER_131_369 ();
 FILLCELL_X1 FILLER_131_371 ();
 FILLCELL_X2 FILLER_131_375 ();
 FILLCELL_X1 FILLER_131_377 ();
 FILLCELL_X8 FILLER_131_398 ();
 FILLCELL_X4 FILLER_131_440 ();
 FILLCELL_X2 FILLER_131_444 ();
 FILLCELL_X2 FILLER_131_517 ();
 FILLCELL_X1 FILLER_131_714 ();
 FILLCELL_X1 FILLER_131_742 ();
 FILLCELL_X1 FILLER_131_749 ();
 FILLCELL_X2 FILLER_131_793 ();
 FILLCELL_X2 FILLER_131_798 ();
 FILLCELL_X1 FILLER_131_800 ();
 FILLCELL_X32 FILLER_131_807 ();
 FILLCELL_X32 FILLER_131_839 ();
 FILLCELL_X32 FILLER_131_871 ();
 FILLCELL_X32 FILLER_131_903 ();
 FILLCELL_X32 FILLER_131_935 ();
 FILLCELL_X8 FILLER_131_967 ();
 FILLCELL_X4 FILLER_131_975 ();
 FILLCELL_X2 FILLER_131_979 ();
 FILLCELL_X1 FILLER_131_981 ();
 FILLCELL_X32 FILLER_132_1 ();
 FILLCELL_X16 FILLER_132_33 ();
 FILLCELL_X8 FILLER_132_49 ();
 FILLCELL_X4 FILLER_132_57 ();
 FILLCELL_X1 FILLER_132_61 ();
 FILLCELL_X8 FILLER_132_65 ();
 FILLCELL_X2 FILLER_132_73 ();
 FILLCELL_X1 FILLER_132_75 ();
 FILLCELL_X8 FILLER_132_79 ();
 FILLCELL_X4 FILLER_132_87 ();
 FILLCELL_X8 FILLER_132_94 ();
 FILLCELL_X4 FILLER_132_102 ();
 FILLCELL_X2 FILLER_132_106 ();
 FILLCELL_X4 FILLER_132_111 ();
 FILLCELL_X1 FILLER_132_115 ();
 FILLCELL_X8 FILLER_132_119 ();
 FILLCELL_X2 FILLER_132_130 ();
 FILLCELL_X1 FILLER_132_132 ();
 FILLCELL_X8 FILLER_132_139 ();
 FILLCELL_X1 FILLER_132_147 ();
 FILLCELL_X1 FILLER_132_151 ();
 FILLCELL_X1 FILLER_132_155 ();
 FILLCELL_X2 FILLER_132_159 ();
 FILLCELL_X2 FILLER_132_164 ();
 FILLCELL_X2 FILLER_132_169 ();
 FILLCELL_X8 FILLER_132_174 ();
 FILLCELL_X2 FILLER_132_182 ();
 FILLCELL_X1 FILLER_132_184 ();
 FILLCELL_X1 FILLER_132_200 ();
 FILLCELL_X4 FILLER_132_207 ();
 FILLCELL_X1 FILLER_132_211 ();
 FILLCELL_X1 FILLER_132_221 ();
 FILLCELL_X4 FILLER_132_231 ();
 FILLCELL_X1 FILLER_132_235 ();
 FILLCELL_X2 FILLER_132_245 ();
 FILLCELL_X1 FILLER_132_250 ();
 FILLCELL_X1 FILLER_132_260 ();
 FILLCELL_X1 FILLER_132_264 ();
 FILLCELL_X1 FILLER_132_268 ();
 FILLCELL_X1 FILLER_132_272 ();
 FILLCELL_X1 FILLER_132_276 ();
 FILLCELL_X4 FILLER_132_286 ();
 FILLCELL_X1 FILLER_132_311 ();
 FILLCELL_X2 FILLER_132_315 ();
 FILLCELL_X2 FILLER_132_320 ();
 FILLCELL_X1 FILLER_132_325 ();
 FILLCELL_X1 FILLER_132_329 ();
 FILLCELL_X1 FILLER_132_333 ();
 FILLCELL_X1 FILLER_132_337 ();
 FILLCELL_X4 FILLER_132_344 ();
 FILLCELL_X2 FILLER_132_348 ();
 FILLCELL_X1 FILLER_132_350 ();
 FILLCELL_X16 FILLER_132_354 ();
 FILLCELL_X4 FILLER_132_370 ();
 FILLCELL_X2 FILLER_132_374 ();
 FILLCELL_X1 FILLER_132_376 ();
 FILLCELL_X2 FILLER_132_386 ();
 FILLCELL_X1 FILLER_132_388 ();
 FILLCELL_X4 FILLER_132_398 ();
 FILLCELL_X8 FILLER_132_405 ();
 FILLCELL_X4 FILLER_132_413 ();
 FILLCELL_X2 FILLER_132_417 ();
 FILLCELL_X2 FILLER_132_422 ();
 FILLCELL_X4 FILLER_132_427 ();
 FILLCELL_X2 FILLER_132_431 ();
 FILLCELL_X1 FILLER_132_433 ();
 FILLCELL_X4 FILLER_132_437 ();
 FILLCELL_X2 FILLER_132_450 ();
 FILLCELL_X2 FILLER_132_455 ();
 FILLCELL_X4 FILLER_132_460 ();
 FILLCELL_X1 FILLER_132_464 ();
 FILLCELL_X2 FILLER_132_468 ();
 FILLCELL_X1 FILLER_132_470 ();
 FILLCELL_X2 FILLER_132_483 ();
 FILLCELL_X1 FILLER_132_485 ();
 FILLCELL_X2 FILLER_132_489 ();
 FILLCELL_X1 FILLER_132_491 ();
 FILLCELL_X1 FILLER_132_506 ();
 FILLCELL_X2 FILLER_132_513 ();
 FILLCELL_X2 FILLER_132_534 ();
 FILLCELL_X1 FILLER_132_539 ();
 FILLCELL_X2 FILLER_132_629 ();
 FILLCELL_X1 FILLER_132_762 ();
 FILLCELL_X2 FILLER_132_793 ();
 FILLCELL_X4 FILLER_132_798 ();
 FILLCELL_X1 FILLER_132_802 ();
 FILLCELL_X32 FILLER_132_806 ();
 FILLCELL_X32 FILLER_132_838 ();
 FILLCELL_X32 FILLER_132_870 ();
 FILLCELL_X32 FILLER_132_902 ();
 FILLCELL_X32 FILLER_132_934 ();
 FILLCELL_X16 FILLER_132_966 ();
endmodule
