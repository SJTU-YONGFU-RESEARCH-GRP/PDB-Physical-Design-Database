module clock_gating (clk_in,
    clk_out,
    enable,
    test_enable);
 input clk_in;
 output clk_out;
 input enable;
 input test_enable;

 wire _0_;
 wire \gen_latch.latch_out ;
 wire net1;
 wire net2;
 wire net3;
 wire clk_in_regs;
 wire clknet_0_clk_in;
 wire clknet_1_0__leaf_clk_in;
 wire clknet_0_clk_in_regs;
 wire clknet_1_0__leaf_clk_in_regs;

 gf180mcu_fd_sc_mcu9t5v0__or2_2 _1_ (.A1(net2),
    .A2(net1),
    .Z(_0_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _2_ (.A1(\gen_latch.latch_out ),
    .A2(clknet_1_0__leaf_clk_in),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__latsnq_1 \gen_latch.latch_out$_DLATCH_N_  (.D(_0_),
    .E(clknet_1_0__leaf_clk_in_regs),
    .Q(\gen_latch.latch_out ));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_53 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_54 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_55 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_56 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_57 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_58 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_59 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_60 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_61 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_62 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_63 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_64 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_65 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_67 ();
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input1 (.I(enable),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(test_enable),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output3 (.I(net3),
    .Z(clk_out));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_regs_0_core_clock (.I(clk_in),
    .Z(clk_in_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_0_clk_in (.I(clk_in),
    .Z(clknet_0_clk_in));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_0__f_clk_in (.I(clknet_0_clk_in),
    .Z(clknet_1_0__leaf_clk_in));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_0_clk_in_regs (.I(clk_in_regs),
    .Z(clknet_0_clk_in_regs));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_0__f_clk_in_regs (.I(clknet_0_clk_in_regs),
    .Z(clknet_1_0__leaf_clk_in_regs));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_178 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_31 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_25_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_252 ();
endmodule
