
* cell configurable_mult
* pin b[5]
* pin a[6]
* pin b[7]
* pin b[4]
* pin a[4]
* pin b[3]
* pin a[3]
* pin b[1]
* pin a[7]
* pin b[0]
* pin NWELL
* pin PWELL
* pin product[1]
* pin product[2]
* pin product[0]
* pin b[2]
* pin a[0]
* pin product[3]
* pin a[2]
* pin a[1]
* pin a[5]
* pin product[4]
* pin b[6]
* pin product[5]
* pin product[6]
* pin product[15]
* pin product[14]
* pin product[12]
* pin product[13]
* pin sign_mode
* pin product[8]
* pin product[11]
* pin product[10]
* pin product[7]
* pin product[9]
.SUBCKT configurable_mult 1 2 3 4 5 6 7 8 9 10 11 12 23 36 37 51 65 87 122 123
+ 160 171 204 290 449 569 596 597 598 599 604 606 607 608 609
* net 1 b[5]
* net 2 a[6]
* net 3 b[7]
* net 4 b[4]
* net 5 a[4]
* net 6 b[3]
* net 7 a[3]
* net 8 b[1]
* net 9 a[7]
* net 10 b[0]
* net 11 NWELL
* net 12 PWELL
* net 23 product[1]
* net 36 product[2]
* net 37 product[0]
* net 51 b[2]
* net 65 a[0]
* net 87 product[3]
* net 122 a[2]
* net 123 a[1]
* net 160 a[5]
* net 171 product[4]
* net 204 b[6]
* net 290 product[5]
* net 449 product[6]
* net 569 product[15]
* net 596 product[14]
* net 597 product[12]
* net 598 product[13]
* net 599 sign_mode
* net 604 product[8]
* net 606 product[11]
* net 607 product[10]
* net 608 product[7]
* net 609 product[9]
* cell instance $5 r0 *1 155.23,152.6
X$5 12 1 18 11 BUF_X16
* cell instance $12 m0 *1 154.66,158.2
X$12 2 11 25 12 BUF_X4
* cell instance $14 r0 *1 155.04,155.4
X$14 12 57 11 3 BUF_X8
* cell instance $21 m0 *1 159.98,155.4
X$21 12 29 11 4 BUF_X8
* cell instance $26 r0 *1 164.54,152.6
X$26 12 15 11 5 BUF_X8
* cell instance $33 m0 *1 169.48,155.4
X$33 12 19 11 6 BUF_X8
* cell instance $39 r0 *1 169.1,152.6
X$39 12 7 14 11 BUF_X16
* cell instance $44 m0 *1 181.83,149.8
X$44 12 8 13 11 BUF_X16
* cell instance $51 r0 *1 186.39,1.4
X$51 12 9 17 11 BUF_X32
* cell instance $57 r0 *1 190.38,155.4
X$57 12 22 11 10 BUF_X8
* cell instance $59 m0 *1 189.24,152.6
X$59 12 24 11 10 BUF_X8
* cell instance $64 r0 *1 158.65,191.8
X$64 508 415 509 555 545 582 12 11 OAI221_X2
* cell instance $68 m0 *1 158.46,194.6
X$68 520 582 561 12 11 581 OR3_X4
* cell instance $70 m0 *1 160.74,194.6
X$70 510 583 12 11 556 NAND2_X2
* cell instance $72 r0 *1 162.07,191.8
X$72 543 544 555 11 545 12 OAI21_X1
* cell instance $74 r0 *1 162.83,191.8
X$74 562 557 511 12 561 11 AOI21_X2
* cell instance $78 m0 *1 163.02,194.6
X$78 579 571 11 12 585 AND2_X1
* cell instance $79 m0 *1 163.78,194.6
X$79 557 521 585 12 562 11 AOI21_X2
* cell instance $80 r0 *1 165.3,191.8
X$80 483 12 11 571 BUF_X1
* cell instance $81 r0 *1 164.54,191.8
X$81 459 521 483 12 11 544 NOR3_X1
* cell instance $85 m0 *1 165.87,194.6
X$85 589 439 484 11 12 587 OAI21_X2
* cell instance $87 r0 *1 167.01,191.8
X$87 525 572 564 11 12 523 OAI21_X2
* cell instance $90 r0 *1 172.33,191.8
X$90 526 513 439 11 12 568 AND3_X1
* cell instance $91 r0 *1 173.28,191.8
X$91 485 513 393 12 593 11 AOI21_X1
* cell instance $92 r0 *1 174.04,191.8
X$92 526 393 513 11 564 12 OAI21_X1
* cell instance $96 m0 *1 167.58,194.6
X$96 586 564 572 11 12 589 OAI21_X2
* cell instance $97 m0 *1 168.91,194.6
X$97 484 485 12 11 586 NOR2_X1
* cell instance $99 m0 *1 169.67,194.6
X$99 592 591 11 12 590 XNOR2_X1
* cell instance $100 m0 *1 170.81,194.6
X$100 568 565 484 439 573 557 11 12 AOI221_X2
* cell instance $103 m0 *1 173.47,194.6
X$103 593 12 11 573 INV_X1
* cell instance $104 m0 *1 173.85,194.6
X$104 485 513 566 12 592 11 AOI21_X2
* cell instance $108 r0 *1 176.7,191.8
X$108 514 513 12 11 558 XOR2_X1
* cell instance $111 m0 *1 177.27,194.6
X$111 558 594 510 11 12 574 MUX2_X2
* cell instance $113 r0 *1 181.64,191.8
X$113 529 527 528 11 12 566 OAI21_X4
* cell instance $114 r0 *1 181.26,191.8
X$114 526 12 11 527 INV_X1
* cell instance $115 r0 *1 184.11,191.8
X$115 393 12 11 529 INV_X1
* cell instance $117 r0 *1 184.68,191.8
X$117 567 443 528 12 11 NOR2_X4
* cell instance $118 r0 *1 186.39,191.8
X$118 519 443 12 11 565 OR2_X2
* cell instance $120 r0 *1 187.53,191.8
X$120 443 12 11 552 INV_X1
* cell instance $121 r0 *1 187.91,191.8
X$121 515 552 529 12 11 595 NAND3_X2
* cell instance $122 r0 *1 189.24,191.8
X$122 530 551 443 491 531 554 11 12 AOI221_X2
* cell instance $126 m0 *1 182.21,194.6
X$126 527 528 12 11 575 XNOR2_X2
* cell instance $129 m0 *1 187.53,194.6
X$129 12 572 595 530 551 11 AOI21_X4
* cell instance $133 r0 *1 193.23,191.8
X$133 492 491 11 12 530 AND2_X2
* cell instance $134 r0 *1 195.7,191.8
X$134 531 492 551 12 563 11 AOI21_X1
* cell instance $137 m0 *1 193.61,194.6
X$137 555 12 11 510 INV_X4
* cell instance $140 m0 *1 195.51,194.6
X$140 491 563 11 12 578 XNOR2_X1
* cell instance $142 r0 *1 197.03,191.8
X$142 517 532 539 11 12 551 OAI21_X4
* cell instance $144 r0 *1 199.5,191.8
X$144 532 469 517 11 560 12 OAI21_X1
* cell instance $147 m0 *1 197.6,194.6
X$147 492 560 12 11 577 XOR2_X1
* cell instance $151 m0 *1 200.07,194.6
X$151 577 559 510 11 12 601 MUX2_X2
* cell instance $153 r0 *1 200.64,191.8
X$153 547 474 11 12 534 XNOR2_X1
* cell instance $157 r0 *1 202.92,191.8
X$157 494 546 12 11 559 XOR2_X1
* cell instance $159 r0 *1 205.01,191.8
X$159 536 12 11 539 BUF_X2
* cell instance $231 r0 *1 197.98,359.8
X$231 605 12 11 608 BUF_X1
* cell instance $235 r0 *1 200.83,359.8
X$235 603 12 11 609 BUF_X1
* cell instance $425 r0 *1 6.65,194.6
X$425 600 12 11 598 BUF_X1
* cell instance $426 r0 *1 7.22,194.6
X$426 576 12 11 569 BUF_X2
* cell instance $427 r0 *1 7.98,194.6
X$427 581 12 11 596 BUF_X1
* cell instance $459 m0 *1 3.23,197.4
X$459 570 12 11 597 BUF_X2
* cell instance $495 r0 *1 159.79,194.6
X$495 556 510 584 11 12 600 OAI21_X4
* cell instance $500 r0 *1 165.87,194.6
X$500 571 12 11 588 BUF_X1
* cell instance $501 r0 *1 164.16,194.6
X$501 588 587 11 584 12 XOR2_X2
* cell instance $505 r0 *1 170.05,194.6
X$505 439 12 11 591 BUF_X1
* cell instance $507 r0 *1 170.62,194.6
X$507 590 548 510 11 12 570 MUX2_X2
* cell instance $511 r0 *1 182.97,194.6
X$511 12 602 489 555 575 11 AOI21_X4
* cell instance $516 r0 *1 199.88,194.6
X$516 578 534 510 11 12 603 MUX2_X2
* cell instance $2812 r0 *1 180.88,155.4
X$2812 12 16 28 102 26 27 11 FA_X1
* cell instance $2813 m0 *1 181.83,158.2
X$2813 19 33 11 12 26 AND2_X2
* cell instance $2820 m0 *1 185.63,158.2
X$2820 13 22 11 20 12 XOR2_X2
* cell instance $2821 r0 *1 186.2,155.4
X$2821 24 13 17 11 12 21 AND3_X1
* cell instance $11551 r0 *1 152.38,180.6
X$11551 319 12 11 374 INV_X1
* cell instance $11555 r0 *1 160.55,180.6
X$11555 12 358 389 404 343 344 11 FA_X1
* cell instance $11564 m0 *1 151.05,183.4
X$11564 278 383 11 12 386 XNOR2_X1
* cell instance $11565 m0 *1 152.19,183.4
X$11565 342 374 383 11 12 611 HA_X1
* cell instance $11570 m0 *1 156.94,183.4
X$11570 206 110 429 11 12 436 HA_X1
* cell instance $11573 r0 *1 165.68,180.6
X$11573 12 281 417 375 359 346 11 FA_X1
* cell instance $11576 r0 *1 168.91,180.6
X$11576 163 12 11 376 INV_X1
* cell instance $11581 m0 *1 168.91,183.4
X$11581 239 376 418 11 12 419 HA_X1
* cell instance $11585 r0 *1 172.71,180.6
X$11585 360 12 11 476 INV_X1
* cell instance $11589 m0 *1 173.47,183.4
X$11589 362 363 390 11 12 391 HA_X1
* cell instance $11590 m0 *1 175.37,183.4
X$11590 365 12 11 406 INV_X1
* cell instance $11594 r0 *1 178.03,180.6
X$11594 325 12 11 408 INV_X1
* cell instance $11597 m0 *1 178.41,183.4
X$11597 408 384 464 11 12 441 HA_X1
* cell instance $11599 r0 *1 180.5,180.6
X$11599 367 12 11 377 INV_X1
* cell instance $11603 m0 *1 181.07,183.4
X$11603 382 12 11 392 INV_X1
* cell instance $11605 r0 *1 182.21,180.6
X$11605 276 12 11 384 INV_X1
* cell instance $11609 r0 *1 185.82,180.6
X$11609 12 369 382 411 370 372 11 FA_X1
* cell instance $11610 r0 *1 188.86,180.6
X$11610 12 333 372 413 371 348 11 FA_X1
* cell instance $11613 r0 *1 194.18,180.6
X$11613 350 349 409 11 12 410 HA_X1
* cell instance $11614 r0 *1 196.08,180.6
X$11614 12 297 351 361 398 249 11 FA_X1
* cell instance $11615 r0 *1 199.12,180.6
X$11615 361 12 11 378 INV_X2
* cell instance $11618 r0 *1 202.92,180.6
X$11618 12 266 379 380 356 354 11 FA_X1
* cell instance $11620 r0 *1 207.48,180.6
X$11620 251 355 400 11 12 424 HA_X1
* cell instance $11651 m0 *1 192.09,183.4
X$11651 12 351 396 412 413 414 11 FA_X1
* cell instance $11652 m0 *1 195.13,183.4
X$11652 410 12 11 414 INV_X1
* cell instance $11655 m0 *1 196.08,183.4
X$11655 409 12 11 398 INV_X1
* cell instance $11659 m0 *1 199.12,183.4
X$11659 12 266 407 405 378 354 11 FA_X1
* cell instance $11662 m0 *1 209.76,183.4
X$11662 400 381 399 11 12 403 HA_X1
* cell instance $13143 r0 *1 152.38,191.8
X$13143 12 538 537 523 507 11 AOI21_X4
* cell instance $13144 r0 *1 154.85,191.8
X$13144 555 540 538 11 12 580 OAI21_X4
* cell instance $13154 m0 *1 154.28,194.6
X$13154 580 478 555 11 12 576 OAI21_X4
* cell instance $13155 m0 *1 156.75,194.6
X$13155 579 11 555 12 BUF_X4
* cell instance $13221 r0 *1 156.94,186.2
X$13221 451 450 436 12 497 11 AOI21_X1
* cell instance $13223 r0 *1 163.78,186.2
X$13223 437 433 483 11 12 459 HA_X1
* cell instance $13235 m0 *1 156.75,189
X$13235 497 458 479 11 12 498 OAI21_X4
* cell instance $13236 m0 *1 159.22,189
X$13236 450 415 12 11 458 NAND2_X1
* cell instance $13237 m0 *1 159.79,189
X$13237 450 12 11 480 INV_X1
* cell instance $13239 m0 *1 163.21,189
X$13239 481 12 11 521 INV_X1
* cell instance $13241 m0 *1 164.35,189
X$13241 459 12 11 482 INV_X1
* cell instance $13243 r0 *1 170.24,186.2
X$13243 454 11 439 12 BUF_X4
* cell instance $13244 r0 *1 168.34,186.2
X$13244 453 438 454 11 12 484 HA_X1
* cell instance $13245 r0 *1 171.57,186.2
X$13245 420 455 11 12 548 XNOR2_X1
* cell instance $13249 m0 *1 172.33,189
X$13249 406 476 501 11 12 485 HA_X1
* cell instance $13251 r0 *1 174.8,186.2
X$13251 419 420 391 12 486 11 AOI21_X1
* cell instance $13253 r0 *1 175.56,186.2
X$13253 420 421 12 11 460 NAND2_X1
* cell instance $13255 r0 *1 176.32,186.2
X$13255 391 421 477 12 455 11 AOI21_X1
* cell instance $13258 r0 *1 178.03,186.2
X$13258 441 464 12 11 442 NOR2_X1
* cell instance $13262 m0 *1 175.56,189
X$13262 461 460 440 11 524 12 OAI21_X1
* cell instance $13264 m0 *1 176.51,189
X$13264 461 463 12 11 477 NAND2_X1
* cell instance $13266 m0 *1 177.27,189
X$13266 442 460 486 11 462 12 OAI21_X1
* cell instance $13268 m0 *1 178.22,189
X$13268 486 504 463 12 11 487 NAND3_X1
* cell instance $13269 m0 *1 178.98,189
X$13269 464 466 488 11 12 465 OAI21_X2
* cell instance $13270 r0 *1 179.17,186.2
X$13270 441 12 11 463 INV_X1
* cell instance $13276 m0 *1 180.31,189
X$13276 466 12 11 504 INV_X1
* cell instance $13278 m0 *1 181.45,189
X$13278 464 466 467 11 12 461 OAI21_X4
* cell instance $13279 m0 *1 183.92,189
X$13279 464 467 466 12 11 490 OR3_X2
* cell instance $13282 r0 *1 188.29,186.2
X$13282 457 394 445 11 12 466 HA_X1
* cell instance $13283 r0 *1 190.76,186.2
X$13283 395 456 506 11 12 443 HA_X1
* cell instance $13287 r0 *1 195.89,186.2
X$13287 407 397 505 11 12 531 HA_X1
* cell instance $13291 r0 *1 200.26,186.2
X$13291 405 424 444 11 12 475 HA_X1
* cell instance $13292 r0 *1 202.16,186.2
X$13292 445 12 11 474 BUF_X1
* cell instance $13293 r0 *1 202.73,186.2
X$13293 445 422 431 12 11 473 NAND3_X1
* cell instance $13294 r0 *1 203.49,186.2
X$13294 422 12 11 470 BUF_X2
* cell instance $13295 r0 *1 204.25,186.2
X$13295 445 12 11 446 BUF_X2
* cell instance $13296 r0 *1 205.01,186.2
X$13296 452 447 12 11 471 NOR2_X1
* cell instance $13297 r0 *1 205.58,186.2
X$13297 447 12 11 448 INV_X1
* cell instance $13324 r0 *1 354.16,186.2
X$13324 426 12 11 449 BUF_X2
* cell instance $13333 m0 *1 201.78,189
X$13333 468 448 473 469 472 467 12 11 OAI221_X2
* cell instance $13334 m0 *1 203.87,189
X$13334 452 446 12 11 472 NAND2_X1
* cell instance $13335 m0 *1 204.44,189
X$13335 495 452 470 11 12 496 OAI21_X4
* cell instance $13336 m0 *1 206.91,189
X$13336 12 488 496 471 518 11 AOI21_X4
* cell instance $13441 r0 *1 151.05,183.4
X$13441 316 386 11 12 537 XNOR2_X1
* cell instance $13443 r0 *1 153.71,183.4
X$13443 387 320 428 11 12 388 HA_X1
* cell instance $13457 m0 *1 155.23,186.2
X$13457 428 199 450 11 12 451 HA_X1
* cell instance $13458 m0 *1 157.13,186.2
X$13458 429 12 11 415 BUF_X1
* cell instance $13460 r0 *1 159.98,183.4
X$13460 357 12 11 432 INV_X1
* cell instance $13464 r0 *1 161.31,183.4
X$13464 389 12 11 416 INV_X1
* cell instance $13467 r0 *1 163.4,183.4
X$13467 404 12 11 433 INV_X1
* cell instance $13470 r0 *1 168.34,183.4
X$13470 375 12 11 438 INV_X2
* cell instance $13476 m0 *1 161.31,186.2
X$13476 432 416 481 11 12 512 HA_X1
* cell instance $13480 m0 *1 165.3,186.2
X$13480 417 12 11 437 INV_X1
* cell instance $13484 m0 *1 168.15,186.2
X$13484 385 12 11 453 INV_X1
* cell instance $13488 m0 *1 169.86,186.2
X$13488 418 12 11 420 BUF_X1
* cell instance $13491 r0 *1 174.04,183.4
X$13491 390 12 11 421 BUF_X1
* cell instance $13498 m0 *1 175.37,186.2
X$13498 419 420 435 12 440 11 AOI21_X1
* cell instance $13499 m0 *1 176.13,186.2
X$13499 434 12 11 435 INV_X1
* cell instance $13501 m0 *1 176.7,186.2
X$13501 391 421 441 12 434 11 AOI21_X1
* cell instance $13503 r0 *1 180.5,183.4
X$13503 392 377 526 11 12 393 HA_X1
* cell instance $13512 m0 *1 188.48,186.2
X$13512 248 12 11 457 INV_X2
* cell instance $13515 m0 *1 190.19,186.2
X$13515 411 12 11 456 INV_X2
* cell instance $13517 r0 *1 191.71,183.4
X$13517 396 12 11 395 INV_X1
* cell instance $13518 r0 *1 191.14,183.4
X$13518 332 12 11 394 INV_X2
* cell instance $13522 r0 *1 196.08,183.4
X$13522 412 12 11 397 INV_X2
* cell instance $13527 r0 *1 202.16,183.4
X$13527 379 352 422 11 12 452 HA_X1
* cell instance $13537 m0 *1 202.16,186.2
X$13537 445 422 12 11 468 NAND2_X1
* cell instance $13538 m0 *1 202.73,186.2
X$13538 431 12 11 423 BUF_X1
* cell instance $13542 m0 *1 205.39,186.2
X$13542 424 380 431 11 12 447 HA_X1
* cell instance $13545 r0 *1 209,183.4
X$13545 12 469 403 399 402 11 AOI21_X4
* cell instance $13546 r0 *1 212.23,183.4
X$13546 400 12 11 430 INV_X1
* cell instance $13549 m0 *1 211.85,186.2
X$13549 12 427 536 426 430 425 11 FA_X1
* cell instance $13550 r0 *1 213.18,183.4
X$13550 381 12 11 427 INV_X1
* cell instance $13552 r0 *1 213.56,183.4
X$13552 401 12 11 425 INV_X2
* cell instance $13553 r0 *1 214.13,183.4
X$13553 401 12 11 402 BUF_X1
* cell instance $13669 r0 *1 154.85,189
X$13669 498 388 12 11 478 XNOR2_X2
* cell instance $13678 m0 *1 153.52,191.8
X$13678 537 523 507 12 11 540 AND3_X4
* cell instance $13681 r0 *1 158.84,189
X$13681 436 480 12 11 509 NAND2_X1
* cell instance $13682 r0 *1 157.89,189
X$13682 555 480 436 12 11 508 OR3_X1
* cell instance $13684 r0 *1 160.93,189
X$13684 482 481 12 11 543 NOR2_X1
* cell instance $13685 r0 *1 161.5,189
X$13685 482 481 555 12 11 511 NAND3_X1
* cell instance $13686 r0 *1 162.26,189
X$13686 12 522 521 499 482 11 AOI21_X4
* cell instance $13687 r0 *1 164.73,189
X$13687 483 500 484 11 12 499 OAI21_X4
* cell instance $13688 r0 *1 167.2,189
X$13688 439 11 500 12 BUF_X4
* cell instance $13691 r0 *1 172.33,189
X$13691 501 12 11 513 BUF_X2
* cell instance $13695 r0 *1 177.84,189
X$13695 462 487 503 11 12 479 OAI21_X4
* cell instance $13696 r0 *1 180.31,189
X$13696 488 11 503 12 BUF_X4
* cell instance $13700 m0 *1 158.46,191.8
X$13700 508 524 542 11 520 12 OAI21_X1
* cell instance $13701 m0 *1 159.22,191.8
X$13701 524 480 415 510 12 11 542 NAND4_X1
* cell instance $13704 m0 *1 160.74,191.8
X$13704 479 415 12 11 583 XNOR2_X2
* cell instance $13707 m0 *1 163.21,191.8
X$13707 522 512 12 507 11 OR2_X4
* cell instance $13710 m0 *1 165.49,191.8
X$13710 459 484 485 512 11 525 12 NOR4_X2
* cell instance $13715 m0 *1 176.89,191.8
X$13715 549 421 12 11 594 XOR2_X1
* cell instance $13718 m0 *1 179.17,191.8
X$13718 463 465 12 11 549 NAND2_X1
* cell instance $13720 r0 *1 182.21,189
X$13720 12 489 555 461 490 11 AOI21_X4
* cell instance $13724 r0 *1 190.95,189
X$13724 506 11 491 12 BUF_X4
* cell instance $13727 m0 *1 182.78,191.8
X$13727 529 527 554 11 12 514 OAI21_X2
* cell instance $13729 m0 *1 185.63,191.8
X$13729 519 12 11 567 BUF_X2
* cell instance $13735 m0 *1 192.28,191.8
X$13735 531 491 12 515 11 NAND2_X4
* cell instance $13736 r0 *1 193.61,189
X$13736 491 492 12 11 516 NAND2_X1
* cell instance $13741 m0 *1 194.18,191.8
X$13741 516 517 553 469 515 519 12 11 OAI221_X2
* cell instance $13743 r0 *1 196.08,189
X$13743 505 12 11 492 BUF_X2
* cell instance $13744 r0 *1 197.03,189
X$13744 502 555 493 12 11 550 MUX2_X1
* cell instance $13746 m0 *1 196.27,191.8
X$13746 493 491 492 12 11 553 NAND3_X2
* cell instance $13748 m0 *1 197.79,191.8
X$13748 550 539 12 11 605 XNOR2_X2
* cell instance $13749 r0 *1 198.93,189
X$13749 475 12 11 517 INV_X1
* cell instance $13752 m0 *1 199.69,191.8
X$13752 533 12 11 532 INV_X2
* cell instance $13753 r0 *1 199.88,189
X$13753 444 12 11 493 BUF_X2
* cell instance $13758 m0 *1 200.26,191.8
X$13758 444 12 11 533 BUF_X1
* cell instance $13761 m0 *1 201.78,191.8
X$13761 423 12 11 502 BUF_X1
* cell instance $13762 m0 *1 202.35,191.8
X$13762 535 469 448 11 546 12 OAI21_X1
* cell instance $13763 m0 *1 203.11,191.8
X$13763 452 494 541 12 547 11 AOI21_X2
* cell instance $13764 r0 *1 204.63,189
X$13764 446 11 495 12 BUF_X4
* cell instance $13765 r0 *1 203.3,189
X$13765 470 11 494 12 BUF_X4
* cell instance $13766 r0 *1 205.96,189
X$13766 423 12 11 535 INV_X1
* cell instance $13796 m0 *1 204.63,191.8
X$13796 535 536 12 11 518 OR2_X2
* cell instance $13797 m0 *1 205.58,191.8
X$13797 448 518 12 11 541 NAND2_X2
* cell instance $13874 m0 *1 1.33,200.2
X$13874 599 12 11 579 CLKBUF_X3
* cell instance $14175 r0 *1 183.16,359.8
X$14175 602 12 11 607 BUF_X1
* cell instance $14344 r0 *1 178.22,359.8
X$14344 574 12 11 606 BUF_X2
* cell instance $18032 m0 *1 201.4,359.8
X$18032 601 12 11 604 BUF_X2
* cell instance $19050 r0 *1 148.2,169.4
X$19050 204 12 11 190 BUF_X2
* cell instance $19053 r0 *1 154.28,169.4
X$19053 25 57 11 12 205 AND2_X1
* cell instance $19056 r0 *1 156.75,169.4
X$19056 25 190 11 12 187 AND2_X1
* cell instance $19057 r0 *1 157.51,169.4
X$19057 72 33 12 11 207 NOR2_X1
* cell instance $19061 m0 *1 152.57,172.2
X$19061 190 43 11 12 224 AND2_X1
* cell instance $19063 m0 *1 153.52,172.2
X$19063 205 224 201 11 12 387 HA_X1
* cell instance $19066 m0 *1 157.13,172.2
X$19066 207 187 225 11 12 255 HA_X1
* cell instance $19067 r0 *1 158.65,169.4
X$19067 12 161 208 209 176 74 11 FA_X1
* cell instance $19070 r0 *1 162.45,169.4
X$19070 12 176 210 211 162 74 11 FA_X1
* cell instance $19072 r0 *1 166.25,169.4
X$19072 188 189 227 11 12 228 HA_X1
* cell instance $19075 r0 *1 171.38,169.4
X$19075 72 14 12 11 230 NOR2_X1
* cell instance $19076 r0 *1 171.95,169.4
X$19076 229 230 263 11 12 257 HA_X1
* cell instance $19078 r0 *1 176.89,169.4
X$19078 114 12 11 259 INV_X1
* cell instance $19081 r0 *1 178.98,169.4
X$19081 57 63 12 11 213 NAND2_X1
* cell instance $19082 r0 *1 179.55,169.4
X$19082 190 14 12 11 214 NAND2_X1
* cell instance $19084 r0 *1 180.31,169.4
X$19084 28 12 11 215 INV_X1
* cell instance $19086 r0 *1 181.45,169.4
X$19086 12 237 236 216 101 185 11 FA_X1
* cell instance $19088 r0 *1 187.53,169.4
X$19088 57 50 12 11 192 NAND2_X1
* cell instance $19091 r0 *1 191.33,169.4
X$19091 12 168 235 232 167 231 11 FA_X1
* cell instance $19094 r0 *1 200.64,169.4
X$19094 35 18 12 226 11 NAND2_X4
* cell instance $19095 r0 *1 202.35,169.4
X$19095 12 193 218 223 226 219 11 FA_X1
* cell instance $19096 r0 *1 205.39,169.4
X$19096 12 223 220 221 143 181 11 FA_X1
* cell instance $19097 r0 *1 208.43,169.4
X$19097 194 12 11 222 INV_X1
* cell instance $19130 m0 *1 161.5,172.2
X$19130 12 225 260 240 210 228 11 FA_X1
* cell instance $19135 m0 *1 167.39,172.2
X$19135 12 227 241 212 257 73 11 FA_X1
* cell instance $19139 m0 *1 175.37,172.2
X$19139 12 259 347 325 233 236 11 FA_X1
* cell instance $19140 m0 *1 178.41,172.2
X$19140 12 215 233 237 213 214 11 FA_X1
* cell instance $19144 m0 *1 186.2,172.2
X$19144 12 235 247 217 258 192 11 FA_X1
* cell instance $19148 m0 *1 192.85,172.2
X$19148 12 119 254 273 232 79 11 FA_X1
* cell instance $19152 m0 *1 202.54,172.2
X$19152 218 12 11 250 INV_X1
* cell instance $19154 m0 *1 209,172.2
X$19154 221 12 11 252 INV_X2
* cell instance $19268 r0 *1 146.87,175
X$19268 293 277 11 12 329 XNOR2_X1
* cell instance $19270 r0 *1 148.77,175
X$19270 12 270 293 295 294 208 11 FA_X1
* cell instance $19272 r0 *1 152.57,175
X$19272 295 12 11 279 INV_X1
* cell instance $19274 r0 *1 155.99,175
X$19274 298 12 11 321 INV_X1
* cell instance $19277 r0 *1 160.17,175
X$19277 12 301 337 322 262 242 11 FA_X1
* cell instance $19280 r0 *1 164.16,175
X$19280 12 242 323 307 302 262 11 FA_X1
* cell instance $19283 r0 *1 168.15,175
X$19283 12 261 281 282 303 307 11 FA_X1
* cell instance $19290 m0 *1 151.62,177.8
X$19290 12 279 317 296 318 337 11 FA_X1
* cell instance $19295 m0 *1 159.03,177.8
X$19295 280 12 11 338 INV_X1
* cell instance $19302 m0 *1 171.38,177.8
X$19302 283 12 11 324 INV_X1
* cell instance $19306 m0 *1 173.85,177.8
X$19306 12 308 341 366 309 310 11 FA_X1
* cell instance $19307 r0 *1 174.8,175
X$19307 305 12 11 309 INV_X1
* cell instance $19311 r0 *1 176.13,175
X$19311 183 12 11 310 INV_X1
* cell instance $19315 r0 *1 178.98,175
X$19315 12 275 340 284 314 28 11 FA_X1
* cell instance $19321 m0 *1 183.73,177.8
X$19321 186 12 11 335 INV_X1
* cell instance $19322 m0 *1 184.11,177.8
X$19322 118 12 11 334 INV_X1
* cell instance $19325 r0 *1 186.96,175
X$19325 312 264 326 11 12 314 HA_X1
* cell instance $19330 r0 *1 191.52,175
X$19330 12 313 315 285 306 231 11 FA_X1
* cell instance $19332 r0 *1 196.27,175
X$19332 12 306 286 299 287 300 11 FA_X1
* cell instance $19333 r0 *1 199.31,175
X$19333 12 297 288 353 273 299 11 FA_X1
* cell instance $19337 m0 *1 194.18,177.8
X$19337 12 311 332 304 288 286 11 FA_X1
* cell instance $19342 r0 *1 202.92,175
X$19342 265 12 11 292 INV_X1
* cell instance $19347 r0 *1 215.65,175
X$19347 289 12 11 291 BUF_X2
* cell instance $19377 m0 *1 203.3,177.8
X$19377 12 220 327 328 106 292 11 FA_X1
* cell instance $19414 m0 *1 353.97,177.8
X$19414 291 12 11 290 BUF_X1
* cell instance $19475 r0 *1 150.1,177.8
X$19475 329 330 11 12 316 XNOR2_X1
* cell instance $19476 r0 *1 151.24,177.8
X$19476 317 331 11 12 330 XNOR2_X1
* cell instance $19487 r0 *1 152.76,177.8
X$19487 318 12 11 319 BUF_X1
* cell instance $19489 r0 *1 155.04,177.8
X$19489 12 296 331 357 336 321 11 FA_X1
* cell instance $19491 m0 *1 153.33,180.6
X$19491 337 12 11 342 INV_X1
* cell instance $19493 r0 *1 158.65,177.8
X$19493 12 318 336 343 338 337 11 FA_X1
* cell instance $19499 m0 *1 162.07,180.6
X$19499 260 12 11 358 INV_X1
* cell instance $19500 m0 *1 162.45,180.6
X$19500 12 323 344 359 322 345 11 FA_X1
* cell instance $19501 r0 *1 163.02,177.8
X$19501 322 12 11 318 BUF_X2
* cell instance $19504 r0 *1 163.97,177.8
X$19504 240 12 11 345 INV_X1
* cell instance $19509 r0 *1 169.86,177.8
X$19509 12 341 385 360 282 324 11 FA_X1
* cell instance $19515 m0 *1 167.2,180.6
X$19515 241 12 11 346 INV_X1
* cell instance $19520 m0 *1 173.28,180.6
X$19520 164 12 11 362 INV_X1
* cell instance $19524 m0 *1 174.99,180.6
X$19524 347 12 11 363 INV_X1
* cell instance $19528 m0 *1 176.7,180.6
X$19528 12 368 365 367 364 366 11 FA_X1
* cell instance $19529 r0 *1 178.03,177.8
X$19529 340 12 11 364 INV_X1
* cell instance $19534 r0 *1 182.02,177.8
X$19534 284 12 11 339 INV_X1
* cell instance $19538 r0 *1 182.78,177.8
X$19538 12 334 368 370 335 339 11 FA_X1
* cell instance $19541 r0 *1 188.29,177.8
X$19541 326 12 11 373 INV_X1
* cell instance $19546 m0 *1 187.15,180.6
X$19546 12 234 369 371 315 373 11 FA_X1
* cell instance $19547 r0 *1 189.24,177.8
X$19547 166 12 11 333 INV_X2
* cell instance $19557 m0 *1 194.56,180.6
X$19557 285 12 11 350 INV_X2
* cell instance $19561 m0 *1 197.22,180.6
X$19561 287 12 11 349 INV_X1
* cell instance $19567 m0 *1 201.4,180.6
X$19567 304 12 11 352 INV_X2
* cell instance $19570 m0 *1 202.54,180.6
X$19570 353 12 11 356 INV_X1
* cell instance $19573 r0 *1 203.11,177.8
X$19573 327 12 11 354 INV_X1
* cell instance $19577 r0 *1 206.15,177.8
X$19577 328 12 11 355 INV_X1
* cell instance $19711 m0 *1 148.39,175
X$19711 208 270 277 11 12 610 HA_X1
* cell instance $19712 m0 *1 150.29,175
X$19712 238 224 270 11 12 278 HA_X1
* cell instance $19713 m0 *1 152.19,175
X$19713 253 224 272 11 12 294 HA_X1
* cell instance $19714 r0 *1 153.71,172.2
X$19714 72 43 12 11 238 NOR2_X1
* cell instance $19716 r0 *1 154.28,172.2
X$19716 72 25 12 11 253 NOR2_X1
* cell instance $19720 r0 *1 165.49,172.2
X$19720 211 12 11 302 INV_X1
* cell instance $19724 m0 *1 154.09,175
X$19724 43 57 11 12 320 AND2_X1
* cell instance $19727 m0 *1 155.99,175
X$19727 12 208 298 280 255 272 11 FA_X1
* cell instance $19730 m0 *1 161.31,175
X$19730 209 12 11 301 INV_X2
* cell instance $19735 m0 *1 170.05,175
X$19735 212 12 11 303 INV_X1
* cell instance $19736 r0 *1 170.62,172.2
X$19736 191 12 11 262 INV_X2
* cell instance $19737 r0 *1 170.05,172.2
X$19737 140 12 11 242 INV_X2
* cell instance $19739 r0 *1 171.95,172.2
X$19739 12 191 243 244 140 45 11 FA_X1
* cell instance $19743 r0 *1 178.98,172.2
X$19743 72 63 12 11 245 NOR2_X1
* cell instance $19744 r0 *1 179.55,172.2
X$19744 214 12 11 246 INV_X1
* cell instance $19747 m0 *1 170.43,175
X$19747 243 12 11 261 INV_X1
* cell instance $19750 m0 *1 171.95,175
X$19750 12 274 283 305 263 138 11 FA_X1
* cell instance $19751 m0 *1 174.99,175
X$19751 244 12 11 308 INV_X1
* cell instance $19756 m0 *1 179.74,175
X$19756 246 245 275 11 12 274 HA_X1
* cell instance $19758 r0 *1 183.54,172.2
X$19758 12 247 276 248 216 256 11 FA_X1
* cell instance $19764 r0 *1 186.96,172.2
X$19764 190 63 12 11 258 NAND2_X1
* cell instance $19767 m0 *1 187.15,175
X$19767 258 12 11 312 INV_X1
* cell instance $19769 m0 *1 187.72,175
X$19769 72 50 12 11 264 NOR2_X1
* cell instance $19771 r0 *1 188.86,172.2
X$19771 12 182 256 311 217 254 11 FA_X1
* cell instance $19777 r0 *1 208.62,172.2
X$19777 12 222 251 269 252 174 11 FA_X1
* cell instance $19806 m0 *1 192.47,175
X$19806 35 72 12 11 313 OR2_X1
* cell instance $19810 m0 *1 197.22,175
X$19810 57 35 12 11 300 NAND2_X1
* cell instance $19811 m0 *1 197.79,175
X$19811 190 50 12 11 306 NAND2_X1
* cell instance $19816 m0 *1 201.4,175
X$19816 35 190 11 12 271 AND2_X1
* cell instance $19818 m0 *1 202.35,175
X$19818 250 271 265 11 12 266 HA_X1
* cell instance $19823 m0 *1 212.99,175
X$19823 195 269 268 11 12 381 HA_X1
* cell instance $19824 m0 *1 214.89,175
X$19824 268 267 289 11 12 401 HA_X1
* cell instance $19971 m0 *1 180.88,155.4
X$19971 15 29 11 12 27 AND2_X2
* cell instance $19973 m0 *1 182.02,155.4
X$19973 14 18 11 16 12 AND2_X4
* cell instance $19978 m0 *1 186.58,155.4
X$19978 12 17 30 11 BUF_X16
* cell instance $20094 m0 *1 168.53,161
X$20094 12 44 92 45 52 31 11 FA_X1
* cell instance $20096 r0 *1 169.67,158.2
X$20096 25 29 12 11 52 NAND2_X1
* cell instance $20097 r0 *1 170.24,158.2
X$20097 18 33 12 11 31 NAND2_X1
* cell instance $20103 m0 *1 174.04,161
X$20103 12 55 138 46 32 56 11 FA_X1
* cell instance $20105 r0 *1 174.23,158.2
X$20105 19 25 11 12 32 AND2_X1
* cell instance $20106 r0 *1 175.75,158.2
X$20106 29 33 11 12 55 AND2_X2
* cell instance $20107 r0 *1 176.7,158.2
X$20107 15 18 11 12 56 AND2_X2
* cell instance $20113 m0 *1 179.36,161
X$20113 46 12 11 98 INV_X1
* cell instance $20116 r0 *1 184.87,158.2
X$20116 13 43 11 12 34 AND2_X1
* cell instance $20117 r0 *1 185.82,158.2
X$20117 30 20 11 117 12 AND2_X4
* cell instance $20151 m0 *1 188.48,161
X$20151 30 22 12 47 11 NAND2_X4
* cell instance $20152 m0 *1 190.19,161
X$20152 57 47 12 11 48 XNOR2_X2
* cell instance $20153 m0 *1 192.09,161
X$20153 58 48 42 11 12 70 HA_X1
* cell instance $20154 m0 *1 193.99,161
X$20154 25 22 12 11 71 NAND2_X1
* cell instance $20157 m0 *1 196.84,161
X$20157 33 22 12 11 69 NAND2_X1
* cell instance $20158 m0 *1 197.41,161
X$20158 33 13 12 11 60 NAND2_X1
* cell instance $20160 m0 *1 198.36,161
X$20160 15 22 12 11 41 NAND2_X1
* cell instance $20161 m0 *1 198.93,161
X$20161 15 49 12 11 61 NAND2_X1
* cell instance $20164 m0 *1 201.21,161
X$20164 15 13 12 11 68 NAND2_X1
* cell instance $20168 m0 *1 204.25,161
X$20168 14 49 12 11 62 NAND2_X1
* cell instance $20171 m0 *1 211.09,161
X$20171 49 50 12 11 81 NAND2_X1
* cell instance $20175 m0 *1 216.6,161
X$20175 49 35 12 11 85 NAND2_X1
* cell instance $20176 m0 *1 217.17,161
X$20176 13 50 12 11 64 NAND2_X1
* cell instance $20178 m0 *1 218.12,161
X$20178 35 13 11 12 54 AND2_X1
* cell instance $20180 m0 *1 219.26,161
X$20180 24 50 11 12 40 AND2_X1
* cell instance $20181 m0 *1 220.02,161
X$20181 54 40 53 11 12 89 HA_X1
* cell instance $20184 m0 *1 228.19,161
X$20184 53 12 11 39 BUF_X2
* cell instance $20186 m0 *1 229.33,161
X$20186 24 35 11 12 38 AND2_X2
* cell instance $20188 m0 *1 230.66,161
X$20188 12 49 11 51 BUF_X8
* cell instance $20213 r0 *1 355.87,158.2
X$20213 39 12 11 23 BUF_X1
* cell instance $20221 m0 *1 360.81,161
X$20221 38 12 11 37 BUF_X1
* cell instance $20293 r0 *1 155.42,163.8
X$20293 33 57 11 12 109 AND2_X1
* cell instance $20303 m0 *1 155.23,166.6
X$20303 12 187 147 135 109 150 11 FA_X1
* cell instance $20304 m0 *1 158.27,166.6
X$20304 135 136 148 11 12 177 HA_X1
* cell instance $20305 r0 *1 159.79,163.8
X$20305 12 148 110 239 127 126 11 FA_X1
* cell instance $20312 m0 *1 161.5,166.6
X$20312 30 29 11 176 12 AND2_X4
* cell instance $20313 m0 *1 163.21,166.6
X$20313 176 162 149 11 12 150 HA_X1
* cell instance $20314 r0 *1 164.16,163.8
X$20314 149 128 151 11 12 127 HA_X1
* cell instance $20318 r0 *1 170.62,163.8
X$20318 131 12 11 112 INV_X1
* cell instance $20323 m0 *1 166.06,166.6
X$20323 151 12 11 178 INV_X1
* cell instance $20325 m0 *1 169.48,166.6
X$20325 17 11 43 12 BUF_X4
* cell instance $20327 m0 *1 171,166.6
X$20327 12 165 137 157 154 156 11 FA_X1
* cell instance $20329 r0 *1 172.14,163.8
X$20329 57 14 12 11 154 NAND2_X1
* cell instance $20332 r0 *1 173.85,163.8
X$20332 12 113 131 114 139 45 11 FA_X1
* cell instance $20335 m0 *1 174.04,166.6
X$20335 138 12 11 156 INV_X1
* cell instance $20336 m0 *1 174.42,166.6
X$20336 157 12 11 139 INV_X1
* cell instance $20340 m0 *1 178.79,166.6
X$20340 115 12 11 191 BUF_X2
* cell instance $20343 r0 *1 179.55,163.8
X$20343 117 133 115 11 12 116 HA_X1
* cell instance $20345 m0 *1 181.07,166.6
X$20345 116 21 12 11 140 OR2_X1
* cell instance $20348 r0 *1 183.54,163.8
X$20348 76 117 134 11 12 159 HA_X1
* cell instance $20351 r0 *1 185.63,163.8
X$20351 12 104 118 166 102 134 11 FA_X1
* cell instance $20356 m0 *1 184.49,166.6
X$20356 159 21 12 11 158 OR2_X2
* cell instance $20359 m0 *1 187.34,166.6
X$20359 155 12 11 184 INV_X2
* cell instance $20360 m0 *1 187.91,166.6
X$20360 102 12 11 155 BUF_X2
* cell instance $20363 r0 *1 191.33,163.8
X$20363 12 59 153 119 47 132 11 FA_X1
* cell instance $20367 m0 *1 192.66,166.6
X$20367 29 14 12 11 168 NAND2_X1
* cell instance $20370 m0 *1 199.5,166.6
X$20370 12 120 287 142 152 141 11 FA_X1
* cell instance $20372 r0 *1 200.83,163.8
X$20372 19 14 12 11 152 NAND2_X1
* cell instance $20374 r0 *1 201.78,163.8
X$20374 29 63 12 11 120 NAND2_X1
* cell instance $20381 m0 *1 206.91,166.6
X$20381 50 19 11 12 180 AND2_X1
* cell instance $20384 r0 *1 210.33,163.8
X$20384 19 35 12 11 121 NAND2_X1
* cell instance $20387 r0 *1 212.23,163.8
X$20387 12 84 146 129 130 121 11 FA_X1
* cell instance $20392 m0 *1 212.8,166.6
X$20392 146 12 11 170 INV_X1
* cell instance $20394 r0 *1 215.84,163.8
X$20394 129 12 11 124 INV_X1
* cell instance $20400 r0 *1 220.59,163.8
X$20400 124 86 125 11 12 173 HA_X1
* cell instance $20404 r0 *1 222.87,163.8
X$20404 125 12 11 88 BUF_X2
* cell instance $20406 r0 *1 229.52,163.8
X$20406 12 50 11 123 BUF_X8
* cell instance $20407 r0 *1 224.77,163.8
X$20407 12 122 63 11 BUF_X16
* cell instance $20535 r0 *1 166.06,161
X$20535 57 15 12 11 91 NAND2_X1
* cell instance $20546 m0 *1 157.51,163.8
X$20546 57 12 11 72 INV_X4
* cell instance $20550 m0 *1 162.07,163.8
X$20550 90 12 11 126 INV_X1
* cell instance $20553 m0 *1 163.02,163.8
X$20553 12 92 90 94 111 91 11 FA_X1
* cell instance $20554 m0 *1 166.06,163.8
X$20554 94 12 11 128 INV_X1
* cell instance $20557 r0 *1 168.53,161
X$20557 92 12 11 73 INV_X1
* cell instance $20560 m0 *1 169.86,163.8
X$20560 44 12 11 74 INV_X2
* cell instance $20562 r0 *1 170.05,161
X$20562 30 19 12 44 11 NAND2_X4
* cell instance $20569 m0 *1 176.32,163.8
X$20569 97 12 11 113 INV_X1
* cell instance $20571 r0 *1 181.26,161
X$20571 99 12 11 100 INV_X1
* cell instance $20572 r0 *1 178.22,161
X$20572 12 75 97 101 98 100 11 FA_X1
* cell instance $20575 m0 *1 180.12,163.8
X$20575 75 12 11 133 INV_X1
* cell instance $20577 r0 *1 182.21,161
X$20577 43 49 12 11 75 NAND2_X1
* cell instance $20582 r0 *1 184.68,161
X$20582 34 76 77 11 12 99 HA_X1
* cell instance $20583 r0 *1 183.92,161
X$20583 49 25 11 12 76 AND2_X1
* cell instance $20590 m0 *1 186.2,163.8
X$20590 77 12 11 103 INV_X1
* cell instance $20595 m0 *1 191.71,163.8
X$20595 72 47 78 11 104 12 OAI21_X1
* cell instance $20596 r0 *1 192.66,161
X$20596 59 12 11 58 INV_X1
* cell instance $20597 r0 *1 192.28,161
X$20597 70 12 11 78 INV_X1
* cell instance $20599 r0 *1 193.23,161
X$20599 25 13 12 11 59 NAND2_X1
* cell instance $20602 m0 *1 192.47,163.8
X$20602 33 49 12 11 132 NAND2_X1
* cell instance $20604 r0 *1 195.89,161
X$20604 42 12 11 202 INV_X1
* cell instance $20607 r0 *1 197.03,161
X$20607 12 60 79 107 71 61 11 FA_X1
* cell instance $20613 m0 *1 200.45,163.8
X$20613 12 142 297 106 108 107 11 FA_X1
* cell instance $20615 r0 *1 201.97,161
X$20615 12 62 108 181 69 68 11 FA_X1
* cell instance $20617 r0 *1 206.72,161
X$20617 49 63 12 11 105 NAND2_X1
* cell instance $20618 r0 *1 207.29,161
X$20618 14 13 12 11 80 NAND2_X1
* cell instance $20620 r0 *1 208.62,161
X$20620 14 24 12 11 82 NAND2_X1
* cell instance $20623 r0 *1 212.99,161
X$20623 63 13 12 11 83 NAND2_X1
* cell instance $20628 m0 *1 205.77,163.8
X$20628 12 41 143 144 105 80 11 FA_X1
* cell instance $20631 m0 *1 210.52,163.8
X$20631 12 83 145 130 81 82 11 FA_X1
* cell instance $20633 r0 *1 214.89,161
X$20633 63 24 12 11 67 NAND2_X1
* cell instance $20635 r0 *1 215.46,161
X$20635 12 64 84 95 67 85 11 FA_X1
* cell instance $20637 r0 *1 219.07,161
X$20637 95 12 11 96 INV_X1
* cell instance $20642 r0 *1 220.78,161
X$20642 89 96 93 11 12 86 HA_X1
* cell instance $20646 r0 *1 224.01,161
X$20646 93 12 11 66 BUF_X2
* cell instance $20670 r0 *1 353.21,161
X$20670 12 65 35 11 BUF_X16
* cell instance $20698 m0 *1 358.34,163.8
X$20698 88 12 11 87 BUF_X1
* cell instance $20701 r0 *1 359.1,161
X$20701 66 12 11 36 BUF_X1
* cell instance $20788 r0 *1 139.46,166.6
X$20788 12 33 11 160 BUF_X8
* cell instance $20807 m0 *1 155.23,169.4
X$20807 12 201 199 206 147 177 11 FA_X1
* cell instance $20810 r0 *1 158.27,166.6
X$20810 18 30 11 161 12 AND2_X4
* cell instance $20811 r0 *1 163.02,166.6
X$20811 18 25 11 12 162 AND2_X1
* cell instance $20816 m0 *1 159.41,169.4
X$20816 161 12 11 136 BUF_X1
* cell instance $20820 m0 *1 165.3,169.4
X$20820 190 33 12 11 111 NAND2_X1
* cell instance $20822 m0 *1 166.06,169.4
X$20822 111 12 11 188 INV_X1
* cell instance $20823 m0 *1 166.44,169.4
X$20823 72 15 12 11 189 NOR2_X1
* cell instance $20826 r0 *1 168.72,166.6
X$20826 12 112 163 164 178 137 11 FA_X1
* cell instance $20833 m0 *1 172.14,169.4
X$20833 190 15 12 11 165 NAND2_X1
* cell instance $20834 m0 *1 172.71,169.4
X$20834 165 12 11 229 INV_X1
* cell instance $20836 r0 *1 177.65,166.6
X$20836 12 46 183 186 115 158 11 FA_X1
* cell instance $20844 r0 *1 185.63,166.6
X$20844 12 103 185 182 184 153 11 FA_X1
* cell instance $20847 r0 *1 191.14,166.6
X$20847 12 132 234 203 167 168 11 FA_X1
* cell instance $20851 r0 *1 201.21,166.6
X$20851 18 50 12 11 141 NAND2_X1
* cell instance $20855 r0 *1 205.77,166.6
X$20855 35 29 11 12 179 AND2_X1
* cell instance $20859 m0 *1 191.9,169.4
X$20859 15 19 12 11 167 NAND2_X1
* cell instance $20861 m0 *1 192.85,169.4
X$20861 18 63 12 11 231 NAND2_X2
* cell instance $20864 m0 *1 194.94,169.4
X$20864 12 203 348 249 202 79 11 FA_X1
* cell instance $20874 m0 *1 203.3,169.4
X$20874 19 63 12 219 11 NAND2_X4
* cell instance $20875 m0 *1 205.01,169.4
X$20875 29 50 12 11 193 NAND2_X2
* cell instance $20877 r0 *1 208.81,166.6
X$20877 175 12 11 169 INV_X1
* cell instance $20878 r0 *1 206.91,166.6
X$20878 180 179 175 11 12 174 HA_X1
* cell instance $20906 r0 *1 357.58,166.6
X$20906 172 12 11 171 BUF_X1
* cell instance $20912 m0 *1 208.05,169.4
X$20912 12 145 194 200 169 144 11 FA_X1
* cell instance $20914 m0 *1 211.85,169.4
X$20914 200 12 11 198 INV_X1
* cell instance $20917 m0 *1 213.37,169.4
X$20917 170 198 196 11 12 195 HA_X1
* cell instance $20918 m0 *1 215.27,169.4
X$20918 196 173 197 11 12 267 HA_X1
* cell instance $20919 m0 *1 217.17,169.4
X$20919 197 12 11 172 BUF_X2
.ENDS configurable_mult

* cell BUF_X32
* pin PWELL,VSS
* pin A
* pin Z
* pin NWELL,VDD
.SUBCKT BUF_X32 1 2 4 5
* net 1 PWELL,VSS
* net 2 A
* net 4 Z
* net 5 NWELL,VDD
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 3 2 5 5 PMOS_VTL L=0.05U W=10.08U AS=0.729225P AD=0.707175P PS=13.025U
+ PD=12.325U
* device instance $17 r0 *1 3.215,0.995 PMOS_VTL
M$17 4 3 5 5 PMOS_VTL L=0.05U W=20.16U AS=1.4175P AD=1.43955P PS=24.66U
+ PD=25.36U
* device instance $49 r0 *1 0.17,0.2975 NMOS_VTL
M$49 3 2 1 1 NMOS_VTL L=0.05U W=6.64U AS=0.4803625P AD=0.4658375P PS=9.37U
+ PD=8.885U
* device instance $65 r0 *1 3.215,0.2975 NMOS_VTL
M$65 4 3 1 1 NMOS_VTL L=0.05U W=13.28U AS=0.93375P AD=0.948275P PS=17.78U
+ PD=18.265U
.ENDS BUF_X32

* cell BUF_X8
* pin PWELL,VSS
* pin Z
* pin NWELL,VDD
* pin A
.SUBCKT BUF_X8 1 3 4 5
* net 1 PWELL,VSS
* net 3 Z
* net 4 NWELL,VDD
* net 5 A
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 2 5 4 4 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 3 2 4 4 PMOS_VTL L=0.05U W=5.04U AS=0.3528P AD=0.37485P PS=6.16U PD=6.86U
* device instance $13 r0 *1 0.17,0.2975 NMOS_VTL
M$13 2 5 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $17 r0 *1 0.93,0.2975 NMOS_VTL
M$17 3 2 1 1 NMOS_VTL L=0.05U W=3.32U AS=0.2324P AD=0.246925P PS=4.44U PD=4.925U
.ENDS BUF_X8

* cell AND2_X4
* pin A2
* pin A1
* pin NWELL,VDD
* pin ZN
* pin PWELL,VSS
.SUBCKT AND2_X4 1 2 4 5 6
* net 1 A2
* net 2 A1
* net 4 NWELL,VDD
* net 5 ZN
* net 6 PWELL,VSS
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 3 1 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 4 2 3 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 5 3 4 4 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $9 r0 *1 0.17,0.2975 NMOS_VTL
M$9 8 1 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $10 r0 *1 0.36,0.2975 NMOS_VTL
M$10 3 2 8 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.55,0.2975 NMOS_VTL
M$11 7 2 3 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 0.74,0.2975 NMOS_VTL
M$12 6 1 7 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.93,0.2975 NMOS_VTL
M$13 5 3 6 6 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS AND2_X4

* cell BUF_X16
* pin PWELL,VSS
* pin A
* pin Z
* pin NWELL,VDD
.SUBCKT BUF_X16 1 2 4 5
* net 1 PWELL,VSS
* net 2 A
* net 4 Z
* net 5 NWELL,VDD
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 3 2 5 5 PMOS_VTL L=0.05U W=5.04U AS=0.37485P AD=0.3528P PS=6.86U PD=6.16U
* device instance $9 r0 *1 1.705,0.995 PMOS_VTL
M$9 4 3 5 5 PMOS_VTL L=0.05U W=10.08U AS=0.7056P AD=0.72765P PS=12.32U PD=13.02U
* device instance $25 r0 *1 0.185,0.2975 NMOS_VTL
M$25 3 2 1 1 NMOS_VTL L=0.05U W=3.32U AS=0.246925P AD=0.2324P PS=4.925U PD=4.44U
* device instance $33 r0 *1 1.705,0.2975 NMOS_VTL
M$33 4 3 1 1 NMOS_VTL L=0.05U W=6.64U AS=0.4648P AD=0.479325P PS=8.88U PD=9.365U
.ENDS BUF_X16

* cell NOR4_X2
* pin A3
* pin A2
* pin A1
* pin A4
* pin NWELL,VDD
* pin ZN
* pin PWELL,VSS
.SUBCKT NOR4_X2 1 2 3 4 5 6 7
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 A4
* net 5 NWELL,VDD
* net 6 ZN
* net 7 PWELL,VSS
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 12 4 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 11 1 12 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 10 2 11 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 6 3 10 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 9 3 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.16,0.995 PMOS_VTL
M$6 13 2 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.35,0.995 PMOS_VTL
M$7 8 1 13 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.54,0.995 PMOS_VTL
M$8 5 4 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 0.21,0.2975 NMOS_VTL
M$9 6 4 7 7 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.072625P PS=1.595U
+ PD=1.595U
* device instance $10 r0 *1 0.4,0.2975 NMOS_VTL
M$10 7 1 6 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $11 r0 *1 0.59,0.2975 NMOS_VTL
M$11 6 2 7 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $12 r0 *1 0.78,0.2975 NMOS_VTL
M$12 7 3 6 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
.ENDS NOR4_X2

* cell OR2_X4
* pin A2
* pin A1
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT OR2_X4 1 2 3 5 6
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 5 ZN
* net 6 NWELL,VDD
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 8 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 4 2 8 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 7 2 4 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 6 1 7 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 5 4 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $9 r0 *1 0.17,0.2975 NMOS_VTL
M$9 4 1 3 3 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $10 r0 *1 0.36,0.2975 NMOS_VTL
M$10 3 2 4 3 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $13 r0 *1 0.93,0.2975 NMOS_VTL
M$13 5 4 3 3 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS OR2_X4

* cell NAND4_X1
* pin A4
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND4_X1 1 2 3 4 5 6 7
* net 1 A4
* net 2 A3
* net 3 A2
* net 4 A1
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 6 2 7 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 7 3 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 6 4 7 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 10 1 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.36,0.2975 NMOS_VTL
M$6 9 2 10 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.55,0.2975 NMOS_VTL
M$7 8 3 9 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.74,0.2975 NMOS_VTL
M$8 7 4 8 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND4_X1

* cell AND2_X1
* pin A1
* pin A2
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND2_X1 1 2 4 5 6
* net 1 A1
* net 2 A2
* net 4 NWELL,VDD
* net 5 PWELL,VSS
* net 6 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 3 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 3 2 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.195 NMOS_VTL
M$4 7 1 3 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $5 r0 *1 0.36,0.195 NMOS_VTL
M$5 5 2 7 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 3 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AND2_X1

* cell XOR2_X2
* pin B
* pin A
* pin NWELL,VDD
* pin Z
* pin PWELL,VSS
.SUBCKT XOR2_X2 1 2 4 5 7
* net 1 B
* net 2 A
* net 4 NWELL,VDD
* net 5 Z
* net 7 PWELL,VSS
* device instance $1 r0 *1 0.2,0.995 PMOS_VTL
M$1 8 2 3 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.39,0.995 PMOS_VTL
M$2 4 1 8 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.58,0.995 PMOS_VTL
M$3 6 3 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $4 r0 *1 0.77,0.995 PMOS_VTL
M$4 5 2 6 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $5 r0 *1 0.96,0.995 PMOS_VTL
M$5 6 1 5 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $9 r0 *1 0.2,0.2975 NMOS_VTL
M$9 3 2 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $10 r0 *1 0.39,0.2975 NMOS_VTL
M$10 7 1 3 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.58,0.2975 NMOS_VTL
M$11 5 3 7 7 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $12 r0 *1 0.77,0.2975 NMOS_VTL
M$12 10 2 5 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.96,0.2975 NMOS_VTL
M$13 7 1 10 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 1.15,0.2975 NMOS_VTL
M$14 9 1 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 1.34,0.2975 NMOS_VTL
M$15 5 2 9 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
.ENDS XOR2_X2

* cell NOR3_X1
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NOR3_X1 1 2 3 4 5 6
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 8 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 7 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.2975 NMOS_VTL
M$4 6 1 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.36,0.2975 NMOS_VTL
M$5 4 2 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 3 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NOR3_X1

* cell AND3_X1
* pin A1
* pin A2
* pin A3
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND3_X1 1 2 3 5 6 7
* net 1 A1
* net 2 A2
* net 3 A3
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 7 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 5 1 4 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 4 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 4 3 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 7 4 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.17,0.195 NMOS_VTL
M$5 8 1 4 6 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $6 r0 *1 0.36,0.195 NMOS_VTL
M$6 9 2 8 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $7 r0 *1 0.55,0.195 NMOS_VTL
M$7 6 3 9 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $8 r0 *1 0.74,0.2975 NMOS_VTL
M$8 7 4 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AND3_X1

* cell AND3_X4
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT AND3_X4 1 2 3 5 6 7
* net 1 A3
* net 2 A2
* net 3 A1
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 6 6 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 6 2 4 6 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 4 3 6 6 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $7 r0 *1 1.31,0.995 PMOS_VTL
M$7 7 4 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $11 r0 *1 0.17,0.2975 NMOS_VTL
M$11 11 1 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $12 r0 *1 0.36,0.2975 NMOS_VTL
M$12 10 2 11 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.55,0.2975 NMOS_VTL
M$13 4 3 10 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 0.74,0.2975 NMOS_VTL
M$14 8 3 4 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 0.93,0.2975 NMOS_VTL
M$15 9 2 8 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 1.12,0.2975 NMOS_VTL
M$16 5 1 9 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $17 r0 *1 1.31,0.2975 NMOS_VTL
M$17 7 4 5 5 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS AND3_X4

* cell OR3_X4
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OR3_X4 1 2 3 5 6 7
* net 1 A3
* net 2 A2
* net 3 A1
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 0.205,0.995 PMOS_VTL
M$1 11 1 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.395,0.995 PMOS_VTL
M$2 10 2 11 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.585,0.995 PMOS_VTL
M$3 4 3 10 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.775,0.995 PMOS_VTL
M$4 9 3 4 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.965,0.995 PMOS_VTL
M$5 8 2 9 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.155,0.995 PMOS_VTL
M$6 6 1 8 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.345,0.995 PMOS_VTL
M$7 7 4 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.177975P AD=0.200025P PS=3.085U
+ PD=3.785U
* device instance $11 r0 *1 0.205,0.2975 NMOS_VTL
M$11 4 1 5 5 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $12 r0 *1 0.395,0.2975 NMOS_VTL
M$12 5 2 4 5 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $13 r0 *1 0.585,0.2975 NMOS_VTL
M$13 4 3 5 5 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $17 r0 *1 1.345,0.2975 NMOS_VTL
M$17 7 4 5 5 NMOS_VTL L=0.05U W=1.66U AS=0.1172375P AD=0.1317625P PS=2.225U
+ PD=2.71U
.ENDS OR3_X4

* cell OR3_X1
* pin A1
* pin A2
* pin A3
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OR3_X1 1 2 3 5 6 7
* net 1 A1
* net 2 A2
* net 3 A3
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 9 1 4 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 8 2 9 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 8 3 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 7 4 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.17,0.195 NMOS_VTL
M$5 5 1 4 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $6 r0 *1 0.36,0.195 NMOS_VTL
M$6 4 2 5 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $7 r0 *1 0.55,0.195 NMOS_VTL
M$7 5 3 4 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $8 r0 *1 0.74,0.2975 NMOS_VTL
M$8 7 4 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OR3_X1

* cell CLKBUF_X3
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT CLKBUF_X3 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 2 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=1.89U AS=0.1323P AD=0.15435P PS=2.31U PD=3.01U
* device instance $5 r0 *1 0.17,0.1875 NMOS_VTL
M$5 3 1 2 3 NMOS_VTL L=0.05U W=0.195U AS=0.020475P AD=0.01365P PS=0.6U PD=0.335U
* device instance $6 r0 *1 0.36,0.1875 NMOS_VTL
M$6 5 2 3 3 NMOS_VTL L=0.05U W=0.585U AS=0.04095P AD=0.047775P PS=1.005U
+ PD=1.27U
.ENDS CLKBUF_X3

* cell NOR2_X1
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NOR2_X1 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 6 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 5 2 6 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.185,0.2975 NMOS_VTL
M$3 5 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $4 r0 *1 0.375,0.2975 NMOS_VTL
M$4 3 2 5 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NOR2_X1

* cell NAND2_X2
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND2_X2 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 ZN
* device instance $1 r0 *1 0.195,0.995 PMOS_VTL
M$1 5 1 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.11025P PS=2.24U PD=2.24U
* device instance $2 r0 *1 0.385,0.995 PMOS_VTL
M$2 4 2 5 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $5 r0 *1 0.195,0.2975 NMOS_VTL
M$5 7 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.385,0.2975 NMOS_VTL
M$6 5 2 7 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.575,0.2975 NMOS_VTL
M$7 6 2 5 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.765,0.2975 NMOS_VTL
M$8 3 1 6 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND2_X2

* cell MUX2_X1
* pin A
* pin S
* pin B
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT MUX2_X1 1 2 3 5 6 8
* net 1 A
* net 2 S
* net 3 B
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 8 Z
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 6 2 4 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 9 1 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.55,1.1525 PMOS_VTL
M$3 7 2 9 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $4 r0 *1 0.74,1.1525 PMOS_VTL
M$4 10 4 7 6 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $5 r0 *1 0.93,1.1525 PMOS_VTL
M$5 10 3 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 8 7 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $7 r0 *1 0.17,0.195 NMOS_VTL
M$7 5 2 4 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $8 r0 *1 0.36,0.195 NMOS_VTL
M$8 12 1 5 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $9 r0 *1 0.55,0.195 NMOS_VTL
M$9 7 4 12 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $10 r0 *1 0.74,0.195 NMOS_VTL
M$10 11 2 7 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $11 r0 *1 0.93,0.195 NMOS_VTL
M$11 5 3 11 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
* device instance $12 r0 *1 1.12,0.2975 NMOS_VTL
M$12 8 7 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS MUX2_X1

* cell NAND3_X1
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND3_X1 1 2 3 4 5 6
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 6 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.2975 NMOS_VTL
M$4 8 1 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.36,0.2975 NMOS_VTL
M$5 7 2 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 3 7 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND3_X1

* cell OAI21_X2
* pin A
* pin B2
* pin B1
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT OAI21_X2 1 2 3 5 6 7
* net 1 A
* net 2 B2
* net 3 B1
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 1 5 5 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 8 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 7 3 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 9 3 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 5 2 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $7 r0 *1 0.17,0.2975 NMOS_VTL
M$7 6 1 4 6 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $9 r0 *1 0.55,0.2975 NMOS_VTL
M$9 7 2 4 6 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $10 r0 *1 0.74,0.2975 NMOS_VTL
M$10 4 3 7 6 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
.ENDS OAI21_X2

* cell OR3_X2
* pin A1
* pin A2
* pin A3
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OR3_X2 1 2 3 5 6 7
* net 1 A1
* net 2 A2
* net 3 A3
* net 5 PWELL,VSS
* net 6 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 9 1 4 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 8 2 9 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 8 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.74,0.995 PMOS_VTL
M$4 7 4 6 6 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $6 r0 *1 0.17,0.2975 NMOS_VTL
M$6 5 1 4 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $7 r0 *1 0.36,0.2975 NMOS_VTL
M$7 4 2 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $8 r0 *1 0.55,0.2975 NMOS_VTL
M$8 5 3 4 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.74,0.2975 NMOS_VTL
M$9 7 4 5 5 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
.ENDS OR3_X2

* cell XNOR2_X2
* pin A
* pin B
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT XNOR2_X2 2 3 4 5 7
* net 2 A
* net 3 B
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 7 ZN
* device instance $1 r0 *1 1.135,0.995 PMOS_VTL
M$1 7 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 1.325,0.995 PMOS_VTL
M$2 9 2 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 1.515,0.995 PMOS_VTL
M$3 5 3 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 1.705,0.995 PMOS_VTL
M$4 8 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $5 r0 *1 0.18,0.995 PMOS_VTL
M$5 7 1 5 5 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $7 r0 *1 0.56,0.995 PMOS_VTL
M$7 1 3 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 0.75,0.995 PMOS_VTL
M$8 5 2 1 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 1.135,0.2975 NMOS_VTL
M$9 6 2 7 4 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $11 r0 *1 1.515,0.2975 NMOS_VTL
M$11 6 3 7 4 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $13 r0 *1 0.18,0.2975 NMOS_VTL
M$13 6 1 4 4 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $15 r0 *1 0.56,0.2975 NMOS_VTL
M$15 10 3 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 0.75,0.2975 NMOS_VTL
M$16 1 2 10 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS XNOR2_X2

* cell AOI21_X4
* pin PWELL,VSS
* pin ZN
* pin A
* pin B2
* pin B1
* pin NWELL,VDD
.SUBCKT AOI21_X4 1 2 3 4 5 11
* net 1 PWELL,VSS
* net 2 ZN
* net 3 A
* net 4 B2
* net 5 B1
* net 11 NWELL,VDD
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 11 3 10 11 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.945,0.995 PMOS_VTL
M$5 2 4 10 11 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $6 r0 *1 1.135,0.995 PMOS_VTL
M$6 10 5 2 11 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.1764P PS=3.08U PD=3.08U
* device instance $13 r0 *1 0.185,0.2975 NMOS_VTL
M$13 2 3 1 1 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $17 r0 *1 0.945,0.2975 NMOS_VTL
M$17 8 4 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $18 r0 *1 1.135,0.2975 NMOS_VTL
M$18 2 5 8 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $19 r0 *1 1.325,0.2975 NMOS_VTL
M$19 9 5 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $20 r0 *1 1.515,0.2975 NMOS_VTL
M$20 1 4 9 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $21 r0 *1 1.705,0.2975 NMOS_VTL
M$21 6 4 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $22 r0 *1 1.895,0.2975 NMOS_VTL
M$22 2 5 6 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $23 r0 *1 2.085,0.2975 NMOS_VTL
M$23 7 5 2 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $24 r0 *1 2.275,0.2975 NMOS_VTL
M$24 1 4 7 1 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI21_X4

* cell MUX2_X2
* pin A
* pin B
* pin S
* pin NWELL,VDD
* pin PWELL,VSS
* pin Z
.SUBCKT MUX2_X2 1 2 3 6 7 8
* net 1 A
* net 2 B
* net 3 S
* net 6 NWELL,VDD
* net 7 PWELL,VSS
* net 8 Z
* device instance $1 r0 *1 1.16,0.995 PMOS_VTL
M$1 8 4 6 6 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.077175P PS=2.24U PD=1.54U
* device instance $3 r0 *1 1.54,1.1525 PMOS_VTL
M$3 9 3 6 6 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.033075P PS=0.77U
+ PD=0.84U
* device instance $4 r0 *1 0.215,0.995 PMOS_VTL
M$4 6 1 5 6 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $5 r0 *1 0.405,0.995 PMOS_VTL
M$5 5 9 6 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 0.595,0.995 PMOS_VTL
M$6 4 2 5 6 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.045675P PS=0.77U PD=0.775U
* device instance $7 r0 *1 0.79,0.995 PMOS_VTL
M$7 5 3 4 6 PMOS_VTL L=0.05U W=0.63U AS=0.045675P AD=0.0693P PS=0.775U PD=1.48U
* device instance $8 r0 *1 1.54,0.195 NMOS_VTL
M$8 9 3 7 7 NMOS_VTL L=0.05U W=0.21U AS=0.021875P AD=0.02205P PS=0.555U PD=0.63U
* device instance $9 r0 *1 1.16,0.2975 NMOS_VTL
M$9 8 4 7 7 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.050925P PS=1.595U
+ PD=1.11U
* device instance $11 r0 *1 0.215,0.2975 NMOS_VTL
M$11 11 1 4 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $12 r0 *1 0.405,0.2975 NMOS_VTL
M$12 7 9 11 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.595,0.2975 NMOS_VTL
M$13 10 2 7 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.0300875P PS=0.555U
+ PD=0.56U
* device instance $14 r0 *1 0.79,0.2975 NMOS_VTL
M$14 4 3 10 7 NMOS_VTL L=0.05U W=0.415U AS=0.0300875P AD=0.043575P PS=0.56U
+ PD=1.04U
.ENDS MUX2_X2

* cell INV_X4
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT INV_X4 1 2 3 4
* net 1 A
* net 2 PWELL,VSS
* net 3 NWELL,VDD
* net 4 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 3 3 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.19845P PS=3.78U PD=3.78U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 4 1 2 2 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.130725P PS=2.705U
+ PD=2.705U
.ENDS INV_X4

* cell AOI21_X1
* pin A
* pin B2
* pin B1
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT AOI21_X1 1 2 3 4 6 7
* net 1 A
* net 2 B2
* net 3 B1
* net 4 PWELL,VSS
* net 6 ZN
* net 7 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 6 2 5 7 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 5 3 6 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 7 1 5 7 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.21,0.2975 NMOS_VTL
M$4 8 2 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.4,0.2975 NMOS_VTL
M$5 6 3 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.59,0.2975 NMOS_VTL
M$6 4 1 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI21_X1

* cell XNOR2_X1
* pin A
* pin B
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT XNOR2_X1 1 2 4 5 7
* net 1 A
* net 2 B
* net 4 NWELL,VDD
* net 5 PWELL,VSS
* net 7 ZN
* device instance $1 r0 *1 0.18,1.1525 PMOS_VTL
M$1 3 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.37,1.1525 PMOS_VTL
M$2 3 2 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.0338625P AD=0.02205P PS=0.775U
+ PD=0.455U
* device instance $3 r0 *1 0.565,0.995 PMOS_VTL
M$3 7 3 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.0338625P AD=0.0441P PS=0.775U PD=0.77U
* device instance $4 r0 *1 0.755,0.995 PMOS_VTL
M$4 8 1 7 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.945,0.995 PMOS_VTL
M$5 4 2 8 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.18,0.195 NMOS_VTL
M$6 9 1 3 5 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $7 r0 *1 0.37,0.195 NMOS_VTL
M$7 5 2 9 5 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0224P PS=0.35U PD=0.56U
* device instance $8 r0 *1 0.565,0.2975 NMOS_VTL
M$8 6 3 5 5 NMOS_VTL L=0.05U W=0.415U AS=0.0224P AD=0.02905P PS=0.56U PD=0.555U
* device instance $9 r0 *1 0.755,0.2975 NMOS_VTL
M$9 7 1 6 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.945,0.2975 NMOS_VTL
M$10 6 2 7 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS XNOR2_X1

* cell AOI221_X2
* pin B1
* pin B2
* pin A
* pin C2
* pin C1
* pin ZN
* pin NWELL,VDD
* pin PWELL,VSS
.SUBCKT AOI221_X2 1 2 3 4 5 6 8 9
* net 1 B1
* net 2 B2
* net 3 A
* net 4 C2
* net 5 C1
* net 6 ZN
* net 8 NWELL,VDD
* net 9 PWELL,VSS
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 3 10 8 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.09135P PS=2.24U PD=1.55U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 8 1 7 8 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 7 2 8 8 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $7 r0 *1 1.32,0.995 PMOS_VTL
M$7 6 4 10 8 PMOS_VTL L=0.05U W=1.26U AS=0.09135P AD=0.11025P PS=1.55U PD=2.24U
* device instance $8 r0 *1 1.51,0.995 PMOS_VTL
M$8 10 5 6 8 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $11 r0 *1 0.17,0.2975 NMOS_VTL
M$11 6 3 9 9 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.060175P PS=1.595U
+ PD=1.12U
* device instance $12 r0 *1 0.36,0.2975 NMOS_VTL
M$12 14 1 6 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $13 r0 *1 0.55,0.2975 NMOS_VTL
M$13 9 2 14 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $14 r0 *1 0.74,0.2975 NMOS_VTL
M$14 13 2 9 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $15 r0 *1 0.93,0.2975 NMOS_VTL
M$15 6 1 13 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $17 r0 *1 1.32,0.2975 NMOS_VTL
M$17 12 4 9 9 NMOS_VTL L=0.05U W=0.415U AS=0.031125P AD=0.02905P PS=0.565U
+ PD=0.555U
* device instance $18 r0 *1 1.51,0.2975 NMOS_VTL
M$18 6 5 12 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $19 r0 *1 1.7,0.2975 NMOS_VTL
M$19 11 5 6 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $20 r0 *1 1.89,0.2975 NMOS_VTL
M$20 9 4 11 9 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI221_X2

* cell NOR2_X4
* pin A2
* pin A1
* pin ZN
* pin PWELL,VSS
* pin NWELL,VDD
.SUBCKT NOR2_X4 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 ZN
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 9 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 3 2 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 8 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 5 1 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 7 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.16,0.995 PMOS_VTL
M$6 3 2 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.35,0.995 PMOS_VTL
M$7 6 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.54,0.995 PMOS_VTL
M$8 5 1 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 0.21,0.2975 NMOS_VTL
M$9 3 1 4 4 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.130725P PS=2.705U
+ PD=2.705U
* device instance $10 r0 *1 0.4,0.2975 NMOS_VTL
M$10 4 2 3 4 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.1162P PS=2.22U PD=2.22U
.ENDS NOR2_X4

* cell NAND3_X2
* pin A3
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND3_X2 1 2 3 4 5 6
* net 1 A3
* net 2 A2
* net 3 A1
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 6 1 5 5 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.11025P PS=2.24U PD=2.24U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 5 2 6 5 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 6 3 5 5 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $7 r0 *1 0.21,0.2975 NMOS_VTL
M$7 10 1 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $8 r0 *1 0.4,0.2975 NMOS_VTL
M$8 9 2 10 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $9 r0 *1 0.59,0.2975 NMOS_VTL
M$9 6 3 9 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.78,0.2975 NMOS_VTL
M$10 8 3 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.97,0.2975 NMOS_VTL
M$11 7 2 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 1.16,0.2975 NMOS_VTL
M$12 4 1 7 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND3_X2

* cell OR2_X2
* pin A1
* pin A2
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OR2_X2 1 2 3 5 6
* net 1 A1
* net 2 A2
* net 3 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 1 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 4 5 5 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 4 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.36,0.2975 NMOS_VTL
M$6 3 2 4 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.55,0.2975 NMOS_VTL
M$7 6 4 3 3 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
.ENDS OR2_X2

* cell OAI21_X1
* pin B2
* pin B1
* pin A
* pin NWELL,VDD
* pin ZN
* pin PWELL,VSS
.SUBCKT OAI21_X1 1 2 3 5 6 7
* net 1 B2
* net 2 B1
* net 3 A
* net 5 NWELL,VDD
* net 6 ZN
* net 7 PWELL,VSS
* device instance $1 r0 *1 0.195,0.995 PMOS_VTL
M$1 8 1 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.385,0.995 PMOS_VTL
M$2 6 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.575,0.995 PMOS_VTL
M$3 5 3 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.195,0.2975 NMOS_VTL
M$4 6 1 4 7 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.385,0.2975 NMOS_VTL
M$5 4 2 6 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $6 r0 *1 0.575,0.2975 NMOS_VTL
M$6 7 3 4 7 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OAI21_X1

* cell NAND2_X4
* pin A2
* pin A1
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT NAND2_X4 1 2 4 5 6
* net 1 A2
* net 2 A1
* net 4 PWELL,VSS
* net 5 ZN
* net 6 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 5 1 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 5 2 6 6 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $9 r0 *1 0.21,0.2975 NMOS_VTL
M$9 4 1 3 4 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $13 r0 *1 0.97,0.2975 NMOS_VTL
M$13 5 2 3 4 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS NAND2_X4

* cell AOI21_X2
* pin A
* pin B2
* pin B1
* pin PWELL,VSS
* pin ZN
* pin NWELL,VDD
.SUBCKT AOI21_X2 1 2 3 4 6 7
* net 1 A
* net 2 B2
* net 3 B1
* net 4 PWELL,VSS
* net 6 ZN
* net 7 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 7 1 5 7 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 6 2 5 7 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 5 3 6 7 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.0882P PS=1.54U PD=1.54U
* device instance $7 r0 *1 0.21,0.2975 NMOS_VTL
M$7 6 1 4 4 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $9 r0 *1 0.59,0.2975 NMOS_VTL
M$9 9 2 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.78,0.2975 NMOS_VTL
M$10 6 3 9 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $11 r0 *1 0.97,0.2975 NMOS_VTL
M$11 8 3 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $12 r0 *1 1.16,0.2975 NMOS_VTL
M$12 4 2 8 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS AOI21_X2

* cell XOR2_X1
* pin A
* pin B
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT XOR2_X1 1 3 4 5 6
* net 1 A
* net 3 B
* net 4 PWELL,VSS
* net 5 NWELL,VDD
* net 6 Z
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 8 1 2 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 8 3 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.0338625P AD=0.02205P PS=0.775U
+ PD=0.455U
* device instance $3 r0 *1 0.555,0.995 PMOS_VTL
M$3 7 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0338625P AD=0.0441P PS=0.775U PD=0.77U
* device instance $4 r0 *1 0.745,0.995 PMOS_VTL
M$4 6 1 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.935,0.995 PMOS_VTL
M$5 7 3 6 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $6 r0 *1 0.17,0.195 NMOS_VTL
M$6 2 1 4 4 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $7 r0 *1 0.36,0.195 NMOS_VTL
M$7 4 3 2 4 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0224P PS=0.35U PD=0.56U
* device instance $8 r0 *1 0.555,0.2975 NMOS_VTL
M$8 6 2 4 4 NMOS_VTL L=0.05U W=0.415U AS=0.0224P AD=0.02905P PS=0.56U PD=0.555U
* device instance $9 r0 *1 0.745,0.2975 NMOS_VTL
M$9 9 1 6 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $10 r0 *1 0.935,0.2975 NMOS_VTL
M$10 4 3 9 4 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS XOR2_X1

* cell OAI221_X2
* pin C2
* pin C1
* pin B1
* pin B2
* pin A
* pin ZN
* pin PWELL,VSS
* pin NWELL,VDD
.SUBCKT OAI221_X2 1 2 3 4 5 7 9 10
* net 1 C2
* net 2 C1
* net 3 B1
* net 4 B2
* net 5 A
* net 7 ZN
* net 9 PWELL,VSS
* net 10 NWELL,VDD
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 12 1 10 10 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 7 2 12 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.59,0.995 PMOS_VTL
M$3 11 2 7 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $4 r0 *1 0.78,0.995 PMOS_VTL
M$4 10 1 11 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.97,0.995 PMOS_VTL
M$5 7 5 10 10 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $6 r0 *1 1.16,0.995 PMOS_VTL
M$6 14 3 7 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.35,0.995 PMOS_VTL
M$7 10 4 14 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.54,0.995 PMOS_VTL
M$8 13 4 10 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $9 r0 *1 1.73,0.995 PMOS_VTL
M$9 7 3 13 10 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $11 r0 *1 0.21,0.2975 NMOS_VTL
M$11 7 1 6 9 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $12 r0 *1 0.4,0.2975 NMOS_VTL
M$12 6 2 7 9 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $15 r0 *1 0.97,0.2975 NMOS_VTL
M$15 8 5 6 9 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
* device instance $16 r0 *1 1.16,0.2975 NMOS_VTL
M$16 9 3 8 9 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
* device instance $17 r0 *1 1.35,0.2975 NMOS_VTL
M$17 8 4 9 9 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.0581P PS=1.11U PD=1.11U
.ENDS OAI221_X2

* cell NAND2_X1
* pin A2
* pin A1
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT NAND2_X1 1 2 3 4 5
* net 1 A2
* net 2 A1
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 5 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.375,0.995 PMOS_VTL
M$2 4 2 5 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.185,0.2975 NMOS_VTL
M$3 6 1 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $4 r0 *1 0.375,0.2975 NMOS_VTL
M$4 5 2 6 3 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS NAND2_X1

* cell BUF_X1
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT BUF_X1 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 2 1 4 4 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.033075P PS=0.77U
+ PD=0.84U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $3 r0 *1 0.17,0.195 NMOS_VTL
M$3 3 1 2 3 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.021875P PS=0.63U PD=0.555U
* device instance $4 r0 *1 0.36,0.2975 NMOS_VTL
M$4 5 2 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS BUF_X1

* cell BUF_X2
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin Z
.SUBCKT BUF_X2 1 3 4 5
* net 1 A
* net 3 PWELL,VSS
* net 4 NWELL,VDD
* net 5 Z
* device instance $1 r0 *1 0.21,0.995 PMOS_VTL
M$1 4 1 2 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.4,0.995 PMOS_VTL
M$2 5 2 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $4 r0 *1 0.21,0.2975 NMOS_VTL
M$4 3 1 2 3 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $5 r0 *1 0.4,0.2975 NMOS_VTL
M$5 5 2 3 3 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
.ENDS BUF_X2

* cell HA_X1
* pin A
* pin B
* pin S
* pin NWELL,VDD
* pin PWELL,VSS
* pin CO
.SUBCKT HA_X1 1 2 4 5 6 9
* net 1 A
* net 2 B
* net 4 S
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 9 CO
* device instance $1 r0 *1 0.785,1.0275 PMOS_VTL
M$1 10 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.0338625P AD=0.02205P PS=0.775U
+ PD=0.455U
* device instance $2 r0 *1 0.975,1.0275 PMOS_VTL
M$2 7 1 10 5 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.033075P PS=0.455U
+ PD=0.84U
* device instance $3 r0 *1 0.21,0.995 PMOS_VTL
M$3 4 2 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $4 r0 *1 0.4,0.995 PMOS_VTL
M$4 3 1 4 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $5 r0 *1 0.59,0.995 PMOS_VTL
M$5 5 7 3 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0338625P PS=0.77U PD=0.775U
* device instance $6 r0 *1 1.345,1.0275 PMOS_VTL
M$6 8 1 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $7 r0 *1 1.535,1.0275 PMOS_VTL
M$7 8 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $8 r0 *1 1.725,0.995 PMOS_VTL
M$8 9 8 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $9 r0 *1 1.345,0.195 NMOS_VTL
M$9 12 1 8 6 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $10 r0 *1 1.535,0.195 NMOS_VTL
M$10 6 2 12 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
* device instance $11 r0 *1 1.725,0.2975 NMOS_VTL
M$11 9 8 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
* device instance $12 r0 *1 0.785,0.195 NMOS_VTL
M$12 7 2 6 6 NMOS_VTL L=0.05U W=0.21U AS=0.0224P AD=0.0147P PS=0.56U PD=0.35U
* device instance $13 r0 *1 0.975,0.195 NMOS_VTL
M$13 6 1 7 6 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.02205P PS=0.35U PD=0.63U
* device instance $14 r0 *1 0.21,0.2975 NMOS_VTL
M$14 11 2 6 6 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $15 r0 *1 0.4,0.2975 NMOS_VTL
M$15 4 1 11 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $16 r0 *1 0.59,0.2975 NMOS_VTL
M$16 6 7 4 6 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.0224P PS=0.555U PD=0.56U
.ENDS HA_X1

* cell FA_X1
* pin PWELL,VSS
* pin B
* pin CO
* pin S
* pin CI
* pin A
* pin NWELL,VDD
.SUBCKT FA_X1 1 2 3 8 11 12 14
* net 1 PWELL,VSS
* net 2 B
* net 3 CO
* net 8 S
* net 11 CI
* net 12 A
* net 14 NWELL,VDD
* device instance $1 r0 *1 0.385,1.0275 PMOS_VTL
M$1 17 2 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $2 r0 *1 0.575,1.0275 PMOS_VTL
M$2 4 12 17 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $3 r0 *1 0.765,1.0275 PMOS_VTL
M$3 15 11 4 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02265P PS=0.455U
+ PD=0.535U
* device instance $4 r0 *1 0.96,1.1025 PMOS_VTL
M$4 14 12 15 14 PMOS_VTL L=0.05U W=0.315U AS=0.02265P AD=0.02205P PS=0.535U
+ PD=0.455U
* device instance $5 r0 *1 1.15,1.1025 PMOS_VTL
M$5 15 2 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.033075P PS=0.455U
+ PD=0.84U
* device instance $6 r0 *1 0.195,0.995 PMOS_VTL
M$6 14 4 3 14 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.033075P PS=1.47U
+ PD=0.77U
* device instance $7 r0 *1 1.49,1.1525 PMOS_VTL
M$7 16 2 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $8 r0 *1 1.68,1.1525 PMOS_VTL
M$8 14 11 16 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $9 r0 *1 1.87,1.1525 PMOS_VTL
M$9 16 12 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $10 r0 *1 2.06,1.1525 PMOS_VTL
M$10 7 4 16 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.023625P PS=0.455U
+ PD=0.465U
* device instance $11 r0 *1 2.26,1.1525 PMOS_VTL
M$11 18 11 7 14 PMOS_VTL L=0.05U W=0.315U AS=0.023625P AD=0.02205P PS=0.465U
+ PD=0.455U
* device instance $12 r0 *1 2.45,1.1525 PMOS_VTL
M$12 19 2 18 14 PMOS_VTL L=0.05U W=0.315U AS=0.02205P AD=0.02205P PS=0.455U
+ PD=0.455U
* device instance $13 r0 *1 2.64,1.1525 PMOS_VTL
M$13 19 12 14 14 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $14 r0 *1 2.83,0.995 PMOS_VTL
M$14 8 7 14 14 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U
+ PD=1.47U
* device instance $15 r0 *1 0.385,0.32 NMOS_VTL
M$15 13 2 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.021875P AD=0.0147P PS=0.555U
+ PD=0.35U
* device instance $16 r0 *1 0.575,0.32 NMOS_VTL
M$16 4 12 13 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $17 r0 *1 0.765,0.32 NMOS_VTL
M$17 5 11 4 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.015225P PS=0.35U
+ PD=0.355U
* device instance $18 r0 *1 0.96,0.32 NMOS_VTL
M$18 1 12 5 1 NMOS_VTL L=0.05U W=0.21U AS=0.015225P AD=0.0147P PS=0.355U
+ PD=0.35U
* device instance $19 r0 *1 1.15,0.32 NMOS_VTL
M$19 5 2 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.02205P PS=0.35U PD=0.63U
* device instance $20 r0 *1 0.195,0.2975 NMOS_VTL
M$20 1 4 3 1 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.021875P PS=1.04U
+ PD=0.555U
* device instance $21 r0 *1 1.49,0.195 NMOS_VTL
M$21 6 2 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $22 r0 *1 1.68,0.195 NMOS_VTL
M$22 1 11 6 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $23 r0 *1 1.87,0.195 NMOS_VTL
M$23 6 12 1 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $24 r0 *1 2.06,0.195 NMOS_VTL
M$24 7 4 6 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.01575P PS=0.35U PD=0.36U
* device instance $25 r0 *1 2.26,0.195 NMOS_VTL
M$25 9 11 7 1 NMOS_VTL L=0.05U W=0.21U AS=0.01575P AD=0.0147P PS=0.36U PD=0.35U
* device instance $26 r0 *1 2.45,0.195 NMOS_VTL
M$26 10 2 9 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.0147P PS=0.35U PD=0.35U
* device instance $27 r0 *1 2.64,0.195 NMOS_VTL
M$27 1 12 10 1 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U
+ PD=0.555U
* device instance $28 r0 *1 2.83,0.2975 NMOS_VTL
M$28 8 7 1 1 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS FA_X1

* cell OAI21_X4
* pin A
* pin B2
* pin B1
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT OAI21_X4 1 2 3 5 6 7
* net 1 A
* net 2 B2
* net 3 B1
* net 5 NWELL,VDD
* net 6 PWELL,VSS
* net 7 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 7 1 5 5 PMOS_VTL L=0.05U W=2.52U AS=0.19845P AD=0.1764P PS=3.78U PD=3.08U
* device instance $5 r0 *1 0.93,0.995 PMOS_VTL
M$5 11 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $6 r0 *1 1.12,0.995 PMOS_VTL
M$6 7 3 11 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $7 r0 *1 1.31,0.995 PMOS_VTL
M$7 10 3 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $8 r0 *1 1.5,0.995 PMOS_VTL
M$8 5 2 10 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $9 r0 *1 1.69,0.995 PMOS_VTL
M$9 9 2 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $10 r0 *1 1.88,0.995 PMOS_VTL
M$10 7 3 9 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $11 r0 *1 2.07,0.995 PMOS_VTL
M$11 8 3 7 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $12 r0 *1 2.26,0.995 PMOS_VTL
M$12 5 2 8 5 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.06615P PS=0.77U PD=1.47U
* device instance $13 r0 *1 0.17,0.2975 NMOS_VTL
M$13 6 1 4 6 NMOS_VTL L=0.05U W=1.66U AS=0.130725P AD=0.1162P PS=2.705U PD=2.22U
* device instance $17 r0 *1 0.93,0.2975 NMOS_VTL
M$17 7 2 4 6 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
* device instance $18 r0 *1 1.12,0.2975 NMOS_VTL
M$18 4 3 7 6 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.1162P PS=2.22U PD=2.22U
.ENDS OAI21_X4

* cell OR2_X1
* pin A1
* pin A2
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT OR2_X1 1 2 3 5 6
* net 1 A1
* net 2 A2
* net 3 PWELL,VSS
* net 5 NWELL,VDD
* net 6 ZN
* device instance $1 r0 *1 0.17,1.1525 PMOS_VTL
M$1 7 1 4 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.84U
+ PD=0.455U
* device instance $2 r0 *1 0.36,1.1525 PMOS_VTL
M$2 7 2 5 5 PMOS_VTL L=0.05U W=0.315U AS=0.033075P AD=0.02205P PS=0.77U
+ PD=0.455U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 4 5 5 PMOS_VTL L=0.05U W=0.63U AS=0.033075P AD=0.06615P PS=0.77U PD=1.47U
* device instance $4 r0 *1 0.17,0.195 NMOS_VTL
M$4 4 1 3 3 NMOS_VTL L=0.05U W=0.21U AS=0.02205P AD=0.0147P PS=0.63U PD=0.35U
* device instance $5 r0 *1 0.36,0.195 NMOS_VTL
M$5 3 2 4 3 NMOS_VTL L=0.05U W=0.21U AS=0.0147P AD=0.021875P PS=0.35U PD=0.555U
* device instance $6 r0 *1 0.55,0.2975 NMOS_VTL
M$6 6 4 3 3 NMOS_VTL L=0.05U W=0.415U AS=0.021875P AD=0.043575P PS=0.555U
+ PD=1.04U
.ENDS OR2_X1

* cell INV_X2
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT INV_X2 1 2 3 4
* net 1 A
* net 2 PWELL,VSS
* net 3 NWELL,VDD
* net 4 ZN
* device instance $1 r0 *1 0.185,0.995 PMOS_VTL
M$1 4 1 3 3 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.11025P PS=2.24U PD=2.24U
* device instance $3 r0 *1 0.185,0.2975 NMOS_VTL
M$3 4 1 2 2 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.072625P PS=1.595U
+ PD=1.595U
.ENDS INV_X2

* cell AND2_X2
* pin A1
* pin A2
* pin NWELL,VDD
* pin PWELL,VSS
* pin ZN
.SUBCKT AND2_X2 1 2 4 5 6
* net 1 A1
* net 2 A2
* net 4 NWELL,VDD
* net 5 PWELL,VSS
* net 6 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 3 1 4 4 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.0441P PS=1.47U PD=0.77U
* device instance $2 r0 *1 0.36,0.995 PMOS_VTL
M$2 4 2 3 4 PMOS_VTL L=0.05U W=0.63U AS=0.0441P AD=0.0441P PS=0.77U PD=0.77U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 6 3 4 4 PMOS_VTL L=0.05U W=1.26U AS=0.0882P AD=0.11025P PS=1.54U PD=2.24U
* device instance $5 r0 *1 0.17,0.2975 NMOS_VTL
M$5 7 1 3 5 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.02905P PS=1.04U
+ PD=0.555U
* device instance $6 r0 *1 0.36,0.2975 NMOS_VTL
M$6 5 2 7 5 NMOS_VTL L=0.05U W=0.415U AS=0.02905P AD=0.02905P PS=0.555U
+ PD=0.555U
* device instance $7 r0 *1 0.55,0.2975 NMOS_VTL
M$7 6 3 5 5 NMOS_VTL L=0.05U W=0.83U AS=0.0581P AD=0.072625P PS=1.11U PD=1.595U
.ENDS AND2_X2

* cell INV_X1
* pin A
* pin PWELL,VSS
* pin NWELL,VDD
* pin ZN
.SUBCKT INV_X1 1 2 3 4
* net 1 A
* net 2 PWELL,VSS
* net 3 NWELL,VDD
* net 4 ZN
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 4 1 3 3 PMOS_VTL L=0.05U W=0.63U AS=0.06615P AD=0.06615P PS=1.47U PD=1.47U
* device instance $2 r0 *1 0.17,0.2975 NMOS_VTL
M$2 4 1 2 2 NMOS_VTL L=0.05U W=0.415U AS=0.043575P AD=0.043575P PS=1.04U
+ PD=1.04U
.ENDS INV_X1

* cell BUF_X4
* pin A
* pin NWELL,VDD
* pin Z
* pin PWELL,VSS
.SUBCKT BUF_X4 1 3 4 5
* net 1 A
* net 3 NWELL,VDD
* net 4 Z
* net 5 PWELL,VSS
* device instance $1 r0 *1 0.17,0.995 PMOS_VTL
M$1 2 1 3 3 PMOS_VTL L=0.05U W=1.26U AS=0.11025P AD=0.0882P PS=2.24U PD=1.54U
* device instance $3 r0 *1 0.55,0.995 PMOS_VTL
M$3 4 2 3 3 PMOS_VTL L=0.05U W=2.52U AS=0.1764P AD=0.19845P PS=3.08U PD=3.78U
* device instance $7 r0 *1 0.17,0.2975 NMOS_VTL
M$7 2 1 5 5 NMOS_VTL L=0.05U W=0.83U AS=0.072625P AD=0.0581P PS=1.595U PD=1.11U
* device instance $9 r0 *1 0.55,0.2975 NMOS_VTL
M$9 4 2 5 5 NMOS_VTL L=0.05U W=1.66U AS=0.1162P AD=0.130725P PS=2.22U PD=2.705U
.ENDS BUF_X4
