module parameterized_sync_reset_counter (clk,
    enable,
    sync_rst,
    tc,
    count);
 input clk;
 input enable;
 input sync_rst;
 output tc;
 output [7:0] count;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;
 wire _30_;
 wire _31_;
 wire _32_;
 wire _33_;
 wire _34_;
 wire _35_;
 wire _36_;
 wire _37_;
 wire _38_;
 wire _39_;
 wire _40_;
 wire _41_;
 wire _42_;
 wire _43_;
 wire _44_;
 wire _45_;
 wire _46_;
 wire _47_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 CLKBUF_X3 _48_ (.A(sync_rst),
    .Z(_08_));
 BUF_X4 _49_ (.A(enable),
    .Z(_09_));
 INV_X1 _50_ (.A(_09_),
    .ZN(_10_));
 NAND2_X1 _51_ (.A1(net1),
    .A2(_10_),
    .ZN(_11_));
 INV_X1 _52_ (.A(net8),
    .ZN(_12_));
 BUF_X2 _53_ (.A(net4),
    .Z(_13_));
 BUF_X2 _54_ (.A(net5),
    .Z(_14_));
 NAND4_X2 _55_ (.A1(_13_),
    .A2(net6),
    .A3(_14_),
    .A4(net7),
    .ZN(_15_));
 BUF_X2 _56_ (.A(net3),
    .Z(_16_));
 NAND2_X1 _57_ (.A1(_16_),
    .A2(_46_),
    .ZN(_17_));
 NOR3_X1 _58_ (.A1(_12_),
    .A2(_15_),
    .A3(_17_),
    .ZN(net9));
 OR3_X1 _59_ (.A1(net1),
    .A2(_10_),
    .A3(_08_),
    .ZN(_18_));
 OAI22_X1 _60_ (.A1(_08_),
    .A2(_11_),
    .B1(net9),
    .B2(_18_),
    .ZN(_00_));
 NAND2_X1 _61_ (.A1(_09_),
    .A2(_47_),
    .ZN(_19_));
 NAND2_X1 _62_ (.A1(net2),
    .A2(_10_),
    .ZN(_20_));
 AOI21_X1 _63_ (.A(_08_),
    .B1(_19_),
    .B2(_20_),
    .ZN(_01_));
 NAND2_X1 _64_ (.A1(_46_),
    .A2(_09_),
    .ZN(_21_));
 XOR2_X1 _65_ (.A(_16_),
    .B(_21_),
    .Z(_22_));
 NOR2_X1 _66_ (.A1(_08_),
    .A2(_22_),
    .ZN(_02_));
 NAND3_X2 _67_ (.A1(_16_),
    .A2(_46_),
    .A3(_09_),
    .ZN(_23_));
 NOR3_X2 _68_ (.A1(_12_),
    .A2(_15_),
    .A3(_23_),
    .ZN(_24_));
 NAND4_X2 _69_ (.A1(_16_),
    .A2(net1),
    .A3(net2),
    .A4(_09_),
    .ZN(_25_));
 XOR2_X1 _70_ (.A(_13_),
    .B(_25_),
    .Z(_26_));
 NOR3_X1 _71_ (.A1(_08_),
    .A2(_24_),
    .A3(_26_),
    .ZN(_03_));
 NAND4_X1 _72_ (.A1(_13_),
    .A2(_16_),
    .A3(_46_),
    .A4(_09_),
    .ZN(_27_));
 XOR2_X1 _73_ (.A(_14_),
    .B(_27_),
    .Z(_28_));
 NOR2_X1 _74_ (.A1(_08_),
    .A2(_28_),
    .ZN(_04_));
 NAND2_X1 _75_ (.A1(_13_),
    .A2(_14_),
    .ZN(_29_));
 OAI21_X1 _76_ (.A(net6),
    .B1(_29_),
    .B2(_25_),
    .ZN(_30_));
 OR3_X1 _77_ (.A1(net6),
    .A2(_29_),
    .A3(_25_),
    .ZN(_31_));
 AOI211_X2 _78_ (.A(_08_),
    .B(_24_),
    .C1(_30_),
    .C2(_31_),
    .ZN(_05_));
 NAND3_X1 _79_ (.A1(_13_),
    .A2(net6),
    .A3(_14_),
    .ZN(_32_));
 OAI21_X1 _80_ (.A(net7),
    .B1(_32_),
    .B2(_23_),
    .ZN(_33_));
 OR3_X1 _81_ (.A1(net7),
    .A2(_32_),
    .A3(_23_),
    .ZN(_34_));
 AOI21_X1 _82_ (.A(_08_),
    .B1(_33_),
    .B2(_34_),
    .ZN(_06_));
 NOR2_X1 _83_ (.A1(_12_),
    .A2(_15_),
    .ZN(_35_));
 NAND2_X1 _84_ (.A1(_23_),
    .A2(_25_),
    .ZN(_36_));
 OR2_X1 _85_ (.A1(_15_),
    .A2(_25_),
    .ZN(_37_));
 AOI221_X1 _86_ (.A(_08_),
    .B1(_35_),
    .B2(_36_),
    .C1(_37_),
    .C2(_12_),
    .ZN(_07_));
 HA_X1 _87_ (.A(net1),
    .B(net2),
    .CO(_46_),
    .S(_47_));
 DFF_X2 \counter_reg[0]$_SDFFE_PP0P_  (.D(_00_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net1),
    .QN(_45_));
 DFF_X2 \counter_reg[1]$_SDFFE_PP0P_  (.D(_01_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net2),
    .QN(_44_));
 DFF_X1 \counter_reg[2]$_SDFFE_PP0P_  (.D(_02_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net3),
    .QN(_43_));
 DFF_X1 \counter_reg[3]$_SDFFE_PP0P_  (.D(_03_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net4),
    .QN(_42_));
 DFF_X1 \counter_reg[4]$_SDFFE_PP0P_  (.D(_04_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net5),
    .QN(_41_));
 DFF_X2 \counter_reg[5]$_SDFFE_PP0P_  (.D(_05_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net6),
    .QN(_40_));
 DFF_X2 \counter_reg[6]$_SDFFE_PP0P_  (.D(_06_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net7),
    .QN(_39_));
 DFF_X1 \counter_reg[7]$_SDFFE_PP0P_  (.D(_07_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net8),
    .QN(_38_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_59 ();
 BUF_X1 output1 (.A(net1),
    .Z(count[0]));
 BUF_X1 output2 (.A(net2),
    .Z(count[1]));
 BUF_X1 output3 (.A(net3),
    .Z(count[2]));
 BUF_X1 output4 (.A(net4),
    .Z(count[3]));
 BUF_X1 output5 (.A(net5),
    .Z(count[4]));
 BUF_X1 output6 (.A(net6),
    .Z(count[5]));
 BUF_X1 output7 (.A(net7),
    .Z(count[6]));
 BUF_X1 output8 (.A(net8),
    .Z(count[7]));
 BUF_X1 output9 (.A(net9),
    .Z(tc));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X16 FILLER_0_65 ();
 FILLCELL_X8 FILLER_0_81 ();
 FILLCELL_X4 FILLER_0_89 ();
 FILLCELL_X2 FILLER_0_96 ();
 FILLCELL_X1 FILLER_0_98 ();
 FILLCELL_X32 FILLER_0_102 ();
 FILLCELL_X32 FILLER_0_134 ();
 FILLCELL_X32 FILLER_0_166 ();
 FILLCELL_X16 FILLER_0_198 ();
 FILLCELL_X8 FILLER_0_214 ();
 FILLCELL_X4 FILLER_0_222 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X1 FILLER_1_225 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X1 FILLER_2_225 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X1 FILLER_3_225 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X1 FILLER_4_225 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X1 FILLER_5_225 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X1 FILLER_6_225 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X1 FILLER_7_225 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X1 FILLER_8_225 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X1 FILLER_9_225 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X8 FILLER_10_33 ();
 FILLCELL_X4 FILLER_10_41 ();
 FILLCELL_X1 FILLER_10_45 ();
 FILLCELL_X8 FILLER_10_63 ();
 FILLCELL_X4 FILLER_10_71 ();
 FILLCELL_X2 FILLER_10_75 ();
 FILLCELL_X1 FILLER_10_77 ();
 FILLCELL_X32 FILLER_10_95 ();
 FILLCELL_X32 FILLER_10_127 ();
 FILLCELL_X32 FILLER_10_159 ();
 FILLCELL_X32 FILLER_10_191 ();
 FILLCELL_X2 FILLER_10_223 ();
 FILLCELL_X1 FILLER_10_225 ();
 FILLCELL_X32 FILLER_11_13 ();
 FILLCELL_X2 FILLER_11_45 ();
 FILLCELL_X1 FILLER_11_47 ();
 FILLCELL_X8 FILLER_11_51 ();
 FILLCELL_X2 FILLER_11_59 ();
 FILLCELL_X8 FILLER_11_65 ();
 FILLCELL_X4 FILLER_11_73 ();
 FILLCELL_X8 FILLER_11_80 ();
 FILLCELL_X2 FILLER_11_88 ();
 FILLCELL_X1 FILLER_11_90 ();
 FILLCELL_X32 FILLER_11_95 ();
 FILLCELL_X32 FILLER_11_127 ();
 FILLCELL_X32 FILLER_11_159 ();
 FILLCELL_X32 FILLER_11_191 ();
 FILLCELL_X2 FILLER_11_223 ();
 FILLCELL_X1 FILLER_11_225 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X8 FILLER_12_33 ();
 FILLCELL_X2 FILLER_12_41 ();
 FILLCELL_X1 FILLER_12_43 ();
 FILLCELL_X16 FILLER_12_50 ();
 FILLCELL_X4 FILLER_12_66 ();
 FILLCELL_X2 FILLER_12_70 ();
 FILLCELL_X1 FILLER_12_72 ();
 FILLCELL_X8 FILLER_12_79 ();
 FILLCELL_X2 FILLER_12_87 ();
 FILLCELL_X1 FILLER_12_89 ();
 FILLCELL_X32 FILLER_12_113 ();
 FILLCELL_X32 FILLER_12_145 ();
 FILLCELL_X8 FILLER_12_177 ();
 FILLCELL_X4 FILLER_12_185 ();
 FILLCELL_X32 FILLER_12_192 ();
 FILLCELL_X2 FILLER_12_224 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X8 FILLER_13_33 ();
 FILLCELL_X2 FILLER_13_41 ();
 FILLCELL_X1 FILLER_13_43 ();
 FILLCELL_X16 FILLER_13_47 ();
 FILLCELL_X8 FILLER_13_68 ();
 FILLCELL_X4 FILLER_13_76 ();
 FILLCELL_X32 FILLER_13_93 ();
 FILLCELL_X32 FILLER_13_125 ();
 FILLCELL_X32 FILLER_13_157 ();
 FILLCELL_X8 FILLER_13_189 ();
 FILLCELL_X2 FILLER_13_197 ();
 FILLCELL_X1 FILLER_13_199 ();
 FILLCELL_X16 FILLER_13_203 ();
 FILLCELL_X4 FILLER_13_219 ();
 FILLCELL_X2 FILLER_13_223 ();
 FILLCELL_X1 FILLER_13_225 ();
 FILLCELL_X4 FILLER_14_1 ();
 FILLCELL_X2 FILLER_14_5 ();
 FILLCELL_X1 FILLER_14_7 ();
 FILLCELL_X2 FILLER_14_11 ();
 FILLCELL_X1 FILLER_14_13 ();
 FILLCELL_X2 FILLER_14_21 ();
 FILLCELL_X1 FILLER_14_23 ();
 FILLCELL_X4 FILLER_14_27 ();
 FILLCELL_X2 FILLER_14_31 ();
 FILLCELL_X16 FILLER_14_43 ();
 FILLCELL_X4 FILLER_14_71 ();
 FILLCELL_X8 FILLER_14_84 ();
 FILLCELL_X2 FILLER_14_92 ();
 FILLCELL_X1 FILLER_14_94 ();
 FILLCELL_X32 FILLER_14_103 ();
 FILLCELL_X32 FILLER_14_135 ();
 FILLCELL_X32 FILLER_14_167 ();
 FILLCELL_X16 FILLER_14_199 ();
 FILLCELL_X8 FILLER_14_215 ();
 FILLCELL_X2 FILLER_14_223 ();
 FILLCELL_X1 FILLER_14_225 ();
 FILLCELL_X8 FILLER_15_1 ();
 FILLCELL_X2 FILLER_15_9 ();
 FILLCELL_X1 FILLER_15_11 ();
 FILLCELL_X8 FILLER_15_42 ();
 FILLCELL_X2 FILLER_15_50 ();
 FILLCELL_X16 FILLER_15_55 ();
 FILLCELL_X2 FILLER_15_71 ();
 FILLCELL_X1 FILLER_15_73 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X32 FILLER_15_161 ();
 FILLCELL_X32 FILLER_15_193 ();
 FILLCELL_X1 FILLER_15_225 ();
 FILLCELL_X1 FILLER_16_1 ();
 FILLCELL_X4 FILLER_16_5 ();
 FILLCELL_X1 FILLER_16_9 ();
 FILLCELL_X16 FILLER_16_18 ();
 FILLCELL_X2 FILLER_16_34 ();
 FILLCELL_X8 FILLER_16_41 ();
 FILLCELL_X4 FILLER_16_49 ();
 FILLCELL_X1 FILLER_16_53 ();
 FILLCELL_X1 FILLER_16_64 ();
 FILLCELL_X4 FILLER_16_69 ();
 FILLCELL_X4 FILLER_16_80 ();
 FILLCELL_X32 FILLER_16_98 ();
 FILLCELL_X32 FILLER_16_130 ();
 FILLCELL_X32 FILLER_16_162 ();
 FILLCELL_X32 FILLER_16_194 ();
 FILLCELL_X8 FILLER_17_1 ();
 FILLCELL_X2 FILLER_17_9 ();
 FILLCELL_X32 FILLER_17_16 ();
 FILLCELL_X8 FILLER_17_48 ();
 FILLCELL_X4 FILLER_17_56 ();
 FILLCELL_X8 FILLER_17_66 ();
 FILLCELL_X4 FILLER_17_74 ();
 FILLCELL_X1 FILLER_17_78 ();
 FILLCELL_X2 FILLER_17_85 ();
 FILLCELL_X1 FILLER_17_87 ();
 FILLCELL_X4 FILLER_17_92 ();
 FILLCELL_X1 FILLER_17_96 ();
 FILLCELL_X32 FILLER_17_101 ();
 FILLCELL_X32 FILLER_17_133 ();
 FILLCELL_X32 FILLER_17_165 ();
 FILLCELL_X16 FILLER_17_197 ();
 FILLCELL_X8 FILLER_17_213 ();
 FILLCELL_X4 FILLER_17_221 ();
 FILLCELL_X1 FILLER_17_225 ();
 FILLCELL_X1 FILLER_18_1 ();
 FILLCELL_X4 FILLER_18_5 ();
 FILLCELL_X1 FILLER_18_9 ();
 FILLCELL_X16 FILLER_18_29 ();
 FILLCELL_X8 FILLER_18_45 ();
 FILLCELL_X4 FILLER_18_53 ();
 FILLCELL_X2 FILLER_18_57 ();
 FILLCELL_X8 FILLER_18_78 ();
 FILLCELL_X1 FILLER_18_86 ();
 FILLCELL_X32 FILLER_18_104 ();
 FILLCELL_X32 FILLER_18_136 ();
 FILLCELL_X16 FILLER_18_168 ();
 FILLCELL_X4 FILLER_18_184 ();
 FILLCELL_X32 FILLER_18_191 ();
 FILLCELL_X2 FILLER_18_223 ();
 FILLCELL_X1 FILLER_18_225 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X32 FILLER_19_193 ();
 FILLCELL_X1 FILLER_19_225 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X32 FILLER_20_193 ();
 FILLCELL_X1 FILLER_20_225 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X32 FILLER_21_193 ();
 FILLCELL_X1 FILLER_21_225 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X32 FILLER_22_193 ();
 FILLCELL_X1 FILLER_22_225 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X32 FILLER_23_193 ();
 FILLCELL_X1 FILLER_23_225 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X32 FILLER_24_193 ();
 FILLCELL_X1 FILLER_24_225 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X32 FILLER_25_193 ();
 FILLCELL_X1 FILLER_25_225 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X32 FILLER_26_193 ();
 FILLCELL_X1 FILLER_26_225 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X1 FILLER_27_225 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X1 FILLER_28_225 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X16 FILLER_29_65 ();
 FILLCELL_X4 FILLER_29_81 ();
 FILLCELL_X1 FILLER_29_85 ();
 FILLCELL_X32 FILLER_29_89 ();
 FILLCELL_X32 FILLER_29_121 ();
 FILLCELL_X32 FILLER_29_153 ();
 FILLCELL_X32 FILLER_29_185 ();
 FILLCELL_X8 FILLER_29_217 ();
 FILLCELL_X1 FILLER_29_225 ();
endmodule
