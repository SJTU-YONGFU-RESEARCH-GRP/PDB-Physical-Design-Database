module wishbone_master (clk,
    read_done,
    read_err,
    read_req,
    rst_n,
    wb_ack_i,
    wb_cyc_o,
    wb_err_i,
    wb_rty_i,
    wb_stb_o,
    wb_we_o,
    write_done,
    write_err,
    write_req,
    read_addr,
    read_data,
    read_sel,
    wb_adr_o,
    wb_dat_i,
    wb_dat_o,
    wb_sel_o,
    wb_tgd_i,
    wb_tgd_o,
    write_addr,
    write_data,
    write_sel);
 input clk;
 output read_done;
 output read_err;
 input read_req;
 input rst_n;
 input wb_ack_i;
 output wb_cyc_o;
 input wb_err_i;
 input wb_rty_i;
 output wb_stb_o;
 output wb_we_o;
 output write_done;
 output write_err;
 input write_req;
 input [31:0] read_addr;
 output [31:0] read_data;
 input [3:0] read_sel;
 output [31:0] wb_adr_o;
 input [31:0] wb_dat_i;
 output [31:0] wb_dat_o;
 output [3:0] wb_sel_o;
 input [0:0] wb_tgd_i;
 output [0:0] wb_tgd_o;
 input [31:0] write_addr;
 input [31:0] write_data;
 input [3:0] write_sel;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire net23;
 wire net22;
 wire _125_;
 wire net21;
 wire net20;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire net19;
 wire net18;
 wire net17;
 wire _135_;
 wire _136_;
 wire _137_;
 wire net16;
 wire _139_;
 wire _140_;
 wire net15;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire net14;
 wire net13;
 wire _174_;
 wire net12;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire net11;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire net10;
 wire _195_;
 wire _196_;
 wire _197_;
 wire net9;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire net8;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire net7;
 wire _218_;
 wire _219_;
 wire _220_;
 wire net6;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire net5;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire net4;
 wire net3;
 wire net2;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire \retry_count[0] ;
 wire \retry_count[1] ;
 wire \retry_count[2] ;
 wire \retry_count[3] ;
 wire \state[0] ;
 wire \state[1] ;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net260;
 wire net247;
 wire net248;
 wire net249;
 wire net1;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire clknet_0_clk;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net261;

 sky130_fd_sc_hd__clkdlybuf4s50_1 input24 (.A(read_addr[2]),
    .X(net23));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input23 (.A(read_addr[29]),
    .X(net22));
 sky130_fd_sc_hd__nor2_1 _273_ (.A(net33),
    .B(net260),
    .Y(_125_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input22 (.A(read_addr[28]),
    .X(net21));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input21 (.A(read_addr[27]),
    .X(net20));
 sky130_fd_sc_hd__nor4b_4 _276_ (.A(net39),
    .B(net73),
    .C(net72),
    .D_N(_003_),
    .Y(_128_));
 sky130_fd_sc_hd__nor2b_1 _277_ (.A(\retry_count[3] ),
    .B_N(_006_),
    .Y(_129_));
 sky130_fd_sc_hd__nor3_1 _278_ (.A(_002_),
    .B(_128_),
    .C(_129_),
    .Y(_130_));
 sky130_fd_sc_hd__a21oi_1 _279_ (.A1(_002_),
    .A2(_125_),
    .B1(_130_),
    .Y(_265_));
 sky130_fd_sc_hd__inv_1 _280_ (.A(\state[0] ),
    .Y(_000_));
 sky130_fd_sc_hd__inv_1 _281_ (.A(\retry_count[0] ),
    .Y(_007_));
 sky130_fd_sc_hd__inv_1 _282_ (.A(\state[1] ),
    .Y(_001_));
 sky130_fd_sc_hd__inv_1 _283_ (.A(\retry_count[1] ),
    .Y(_008_));
 sky130_fd_sc_hd__nand2_2 _284_ (.A(net39),
    .B(_004_),
    .Y(_131_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input20 (.A(read_addr[26]),
    .X(net19));
 sky130_fd_sc_hd__mux2_2 _286_ (.A0(net40),
    .A1(net143),
    .S(_131_),
    .X(_012_));
 sky130_fd_sc_hd__mux2_2 _287_ (.A0(net41),
    .A1(net144),
    .S(_131_),
    .X(_013_));
 sky130_fd_sc_hd__mux2_2 _288_ (.A0(net42),
    .A1(net145),
    .S(_131_),
    .X(_014_));
 sky130_fd_sc_hd__mux2_2 _289_ (.A0(net43),
    .A1(net146),
    .S(_131_),
    .X(_015_));
 sky130_fd_sc_hd__mux2_2 _290_ (.A0(net44),
    .A1(net147),
    .S(_131_),
    .X(_016_));
 sky130_fd_sc_hd__mux2_2 _291_ (.A0(net45),
    .A1(net148),
    .S(_131_),
    .X(_017_));
 sky130_fd_sc_hd__mux2_2 _292_ (.A0(net46),
    .A1(net149),
    .S(_131_),
    .X(_018_));
 sky130_fd_sc_hd__mux2_2 _293_ (.A0(net47),
    .A1(net150),
    .S(_131_),
    .X(_019_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input19 (.A(read_addr[25]),
    .X(net18));
 sky130_fd_sc_hd__mux2_2 _295_ (.A0(net48),
    .A1(net151),
    .S(_131_),
    .X(_020_));
 sky130_fd_sc_hd__mux2_2 _296_ (.A0(net49),
    .A1(net152),
    .S(_131_),
    .X(_021_));
 sky130_fd_sc_hd__mux2_2 _297_ (.A0(net50),
    .A1(net153),
    .S(_131_),
    .X(_022_));
 sky130_fd_sc_hd__mux2_2 _298_ (.A0(net51),
    .A1(net154),
    .S(_131_),
    .X(_023_));
 sky130_fd_sc_hd__mux2_2 _299_ (.A0(net52),
    .A1(net155),
    .S(_131_),
    .X(_024_));
 sky130_fd_sc_hd__mux2_2 _300_ (.A0(net53),
    .A1(net156),
    .S(_131_),
    .X(_025_));
 sky130_fd_sc_hd__mux2_2 _301_ (.A0(net54),
    .A1(net157),
    .S(_131_),
    .X(_026_));
 sky130_fd_sc_hd__mux2_2 _302_ (.A0(net55),
    .A1(net158),
    .S(_131_),
    .X(_027_));
 sky130_fd_sc_hd__mux2_2 _303_ (.A0(net56),
    .A1(net159),
    .S(_131_),
    .X(_028_));
 sky130_fd_sc_hd__mux2_2 _304_ (.A0(net57),
    .A1(net160),
    .S(_131_),
    .X(_029_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input18 (.A(read_addr[24]),
    .X(net17));
 sky130_fd_sc_hd__mux2_2 _306_ (.A0(net58),
    .A1(net161),
    .S(_131_),
    .X(_030_));
 sky130_fd_sc_hd__mux2_2 _307_ (.A0(net59),
    .A1(net162),
    .S(_131_),
    .X(_031_));
 sky130_fd_sc_hd__mux2_2 _308_ (.A0(net60),
    .A1(net163),
    .S(_131_),
    .X(_032_));
 sky130_fd_sc_hd__mux2_2 _309_ (.A0(net61),
    .A1(net164),
    .S(_131_),
    .X(_033_));
 sky130_fd_sc_hd__mux2_2 _310_ (.A0(net62),
    .A1(net165),
    .S(_131_),
    .X(_034_));
 sky130_fd_sc_hd__mux2_2 _311_ (.A0(net63),
    .A1(net166),
    .S(_131_),
    .X(_035_));
 sky130_fd_sc_hd__mux2_2 _312_ (.A0(net64),
    .A1(net167),
    .S(_131_),
    .X(_036_));
 sky130_fd_sc_hd__mux2_2 _313_ (.A0(net65),
    .A1(net168),
    .S(_131_),
    .X(_037_));
 sky130_fd_sc_hd__mux2_2 _314_ (.A0(net66),
    .A1(net169),
    .S(_131_),
    .X(_038_));
 sky130_fd_sc_hd__mux2_2 _315_ (.A0(net67),
    .A1(net170),
    .S(_131_),
    .X(_039_));
 sky130_fd_sc_hd__mux2_2 _316_ (.A0(net68),
    .A1(net171),
    .S(_131_),
    .X(_040_));
 sky130_fd_sc_hd__mux2_2 _317_ (.A0(net69),
    .A1(net172),
    .S(_131_),
    .X(_041_));
 sky130_fd_sc_hd__mux2_2 _318_ (.A0(net70),
    .A1(net173),
    .S(_131_),
    .X(_042_));
 sky130_fd_sc_hd__mux2_2 _319_ (.A0(net71),
    .A1(net174),
    .S(_131_),
    .X(_043_));
 sky130_fd_sc_hd__inv_1 _320_ (.A(net33),
    .Y(_135_));
 sky130_fd_sc_hd__o21ai_1 _321_ (.A1(_135_),
    .A2(net260),
    .B1(_002_),
    .Y(_136_));
 sky130_fd_sc_hd__a21oi_1 _322_ (.A1(net39),
    .A2(_136_),
    .B1(net175),
    .Y(_137_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input17 (.A(read_addr[23]),
    .X(net16));
 sky130_fd_sc_hd__nand3b_1 _324_ (.A_N(net260),
    .B(_002_),
    .C(net33),
    .Y(_139_));
 sky130_fd_sc_hd__a21oi_1 _325_ (.A1(net175),
    .A2(_139_),
    .B1(_004_),
    .Y(_140_));
 sky130_fd_sc_hd__nor2_1 _326_ (.A(_137_),
    .B(_140_),
    .Y(_044_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input16 (.A(read_addr[22]),
    .X(net15));
 sky130_fd_sc_hd__nor3_1 _328_ (.A(_006_),
    .B(_005_),
    .C(_004_),
    .Y(_142_));
 sky130_fd_sc_hd__inv_1 _329_ (.A(\retry_count[3] ),
    .Y(_143_));
 sky130_fd_sc_hd__o21ai_0 _330_ (.A1(_143_),
    .A2(net247),
    .B1(_006_),
    .Y(_144_));
 sky130_fd_sc_hd__nor2_1 _331_ (.A(net39),
    .B(net72),
    .Y(_145_));
 sky130_fd_sc_hd__a21oi_1 _332_ (.A1(_004_),
    .A2(_145_),
    .B1(_005_),
    .Y(_146_));
 sky130_fd_sc_hd__a41oi_1 _333_ (.A1(_131_),
    .A2(_136_),
    .A3(_144_),
    .A4(_146_),
    .B1(net176),
    .Y(_147_));
 sky130_fd_sc_hd__a31oi_1 _334_ (.A1(_131_),
    .A2(_136_),
    .A3(_142_),
    .B1(_147_),
    .Y(_045_));
 sky130_fd_sc_hd__nand2_1 _335_ (.A(net73),
    .B(_145_),
    .Y(_148_));
 sky130_fd_sc_hd__a21oi_1 _336_ (.A1(_003_),
    .A2(_148_),
    .B1(_006_),
    .Y(_149_));
 sky130_fd_sc_hd__nor3b_2 _337_ (.A(net39),
    .B(net72),
    .C_N(net73),
    .Y(_150_));
 sky130_fd_sc_hd__nand3b_1 _338_ (.A_N(_006_),
    .B(_003_),
    .C(_150_),
    .Y(_151_));
 sky130_fd_sc_hd__mux2i_1 _339_ (.A0(_149_),
    .A1(_151_),
    .S(_007_),
    .Y(_046_));
 sky130_fd_sc_hd__inv_1 _340_ (.A(_010_),
    .Y(_152_));
 sky130_fd_sc_hd__o22ai_1 _341_ (.A1(_008_),
    .A2(_149_),
    .B1(_151_),
    .B2(_152_),
    .Y(_047_));
 sky130_fd_sc_hd__nand2_1 _342_ (.A(_011_),
    .B(_150_),
    .Y(_153_));
 sky130_fd_sc_hd__nor2_1 _343_ (.A(_006_),
    .B(\retry_count[2] ),
    .Y(_154_));
 sky130_fd_sc_hd__nand2_1 _344_ (.A(_003_),
    .B(_154_),
    .Y(_155_));
 sky130_fd_sc_hd__a21oi_1 _345_ (.A1(_003_),
    .A2(_153_),
    .B1(_006_),
    .Y(_156_));
 sky130_fd_sc_hd__inv_1 _346_ (.A(\retry_count[2] ),
    .Y(_157_));
 sky130_fd_sc_hd__o22ai_1 _347_ (.A1(_153_),
    .A2(_155_),
    .B1(_156_),
    .B2(_157_),
    .Y(_048_));
 sky130_fd_sc_hd__nand4_1 _348_ (.A(\retry_count[2] ),
    .B(\retry_count[0] ),
    .C(\retry_count[1] ),
    .D(_150_),
    .Y(_158_));
 sky130_fd_sc_hd__nor2_1 _349_ (.A(_006_),
    .B(\retry_count[3] ),
    .Y(_159_));
 sky130_fd_sc_hd__nand2_1 _350_ (.A(_003_),
    .B(_159_),
    .Y(_160_));
 sky130_fd_sc_hd__a21oi_1 _351_ (.A1(_003_),
    .A2(_158_),
    .B1(_006_),
    .Y(_161_));
 sky130_fd_sc_hd__o22ai_1 _352_ (.A1(_158_),
    .A2(_160_),
    .B1(_161_),
    .B2(_143_),
    .Y(_049_));
 sky130_fd_sc_hd__a221oi_1 _353_ (.A1(_003_),
    .A2(_145_),
    .B1(_129_),
    .B2(net247),
    .C1(_002_),
    .Y(_162_));
 sky130_fd_sc_hd__nor2b_1 _354_ (.A(net260),
    .B_N(_002_),
    .Y(_163_));
 sky130_fd_sc_hd__a21o_1 _355_ (.A1(_002_),
    .A2(_125_),
    .B1(_128_),
    .X(_164_));
 sky130_fd_sc_hd__nand2_1 _356_ (.A(\state[0] ),
    .B(_164_),
    .Y(_165_));
 sky130_fd_sc_hd__o31ai_1 _357_ (.A1(_128_),
    .A2(_162_),
    .A3(_163_),
    .B1(_165_),
    .Y(_050_));
 sky130_fd_sc_hd__inv_1 _358_ (.A(net247),
    .Y(_166_));
 sky130_fd_sc_hd__a221oi_1 _359_ (.A1(_003_),
    .A2(_145_),
    .B1(_129_),
    .B2(_166_),
    .C1(_002_),
    .Y(_167_));
 sky130_fd_sc_hd__nand2_2 _360_ (.A(net260),
    .B(_002_),
    .Y(_168_));
 sky130_fd_sc_hd__nand2b_1 _361_ (.A_N(_164_),
    .B(net257),
    .Y(_169_));
 sky130_fd_sc_hd__nand2_1 _362_ (.A(\state[1] ),
    .B(_164_),
    .Y(_170_));
 sky130_fd_sc_hd__o21ai_0 _363_ (.A1(_167_),
    .A2(_169_),
    .B1(_170_),
    .Y(_051_));
 sky130_fd_sc_hd__o21ai_4 _364_ (.A1(net33),
    .A2(net260),
    .B1(_002_),
    .Y(_171_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input15 (.A(read_addr[21]),
    .X(net14));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input14 (.A(read_addr[20]),
    .X(net13));
 sky130_fd_sc_hd__mux2i_1 _367_ (.A0(net1),
    .A1(net74),
    .S(net260),
    .Y(_174_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input13 (.A(read_addr[1]),
    .X(net12));
 sky130_fd_sc_hd__nand2_1 _369_ (.A(net177),
    .B(net256),
    .Y(_176_));
 sky130_fd_sc_hd__o21ai_0 _370_ (.A1(net256),
    .A2(_174_),
    .B1(_176_),
    .Y(_052_));
 sky130_fd_sc_hd__mux2i_1 _371_ (.A0(net2),
    .A1(net75),
    .S(net260),
    .Y(_177_));
 sky130_fd_sc_hd__nand2_1 _372_ (.A(net178),
    .B(net256),
    .Y(_178_));
 sky130_fd_sc_hd__o21ai_0 _373_ (.A1(net256),
    .A2(_177_),
    .B1(_178_),
    .Y(_053_));
 sky130_fd_sc_hd__mux2i_1 _374_ (.A0(net3),
    .A1(net76),
    .S(net260),
    .Y(_179_));
 sky130_fd_sc_hd__nand2_1 _375_ (.A(net179),
    .B(net256),
    .Y(_180_));
 sky130_fd_sc_hd__o21ai_0 _376_ (.A1(net256),
    .A2(_179_),
    .B1(_180_),
    .Y(_054_));
 sky130_fd_sc_hd__mux2i_1 _377_ (.A0(net4),
    .A1(net77),
    .S(net260),
    .Y(_181_));
 sky130_fd_sc_hd__nand2_1 _378_ (.A(net180),
    .B(net256),
    .Y(_182_));
 sky130_fd_sc_hd__o21ai_0 _379_ (.A1(net256),
    .A2(_181_),
    .B1(_182_),
    .Y(_055_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input12 (.A(read_addr[19]),
    .X(net11));
 sky130_fd_sc_hd__mux2i_1 _381_ (.A0(net5),
    .A1(net78),
    .S(net260),
    .Y(_184_));
 sky130_fd_sc_hd__nand2_1 _382_ (.A(net181),
    .B(net256),
    .Y(_185_));
 sky130_fd_sc_hd__o21ai_1 _383_ (.A1(net256),
    .A2(_184_),
    .B1(_185_),
    .Y(_056_));
 sky130_fd_sc_hd__mux2i_1 _384_ (.A0(net6),
    .A1(net79),
    .S(net260),
    .Y(_186_));
 sky130_fd_sc_hd__nand2_1 _385_ (.A(net182),
    .B(net256),
    .Y(_187_));
 sky130_fd_sc_hd__o21ai_0 _386_ (.A1(net256),
    .A2(_186_),
    .B1(_187_),
    .Y(_057_));
 sky130_fd_sc_hd__mux2i_1 _387_ (.A0(net7),
    .A1(net80),
    .S(net260),
    .Y(_188_));
 sky130_fd_sc_hd__nand2_1 _388_ (.A(net183),
    .B(net256),
    .Y(_189_));
 sky130_fd_sc_hd__o21ai_0 _389_ (.A1(net256),
    .A2(_188_),
    .B1(_189_),
    .Y(_058_));
 sky130_fd_sc_hd__mux2i_1 _390_ (.A0(net8),
    .A1(net81),
    .S(net260),
    .Y(_190_));
 sky130_fd_sc_hd__nand2_1 _391_ (.A(net184),
    .B(net256),
    .Y(_191_));
 sky130_fd_sc_hd__o21ai_0 _392_ (.A1(net256),
    .A2(_190_),
    .B1(_191_),
    .Y(_059_));
 sky130_fd_sc_hd__mux2i_1 _393_ (.A0(net9),
    .A1(net82),
    .S(net260),
    .Y(_192_));
 sky130_fd_sc_hd__nand2_1 _394_ (.A(net185),
    .B(net256),
    .Y(_193_));
 sky130_fd_sc_hd__o21ai_0 _395_ (.A1(net256),
    .A2(_192_),
    .B1(_193_),
    .Y(_060_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input11 (.A(read_addr[18]),
    .X(net10));
 sky130_fd_sc_hd__mux2i_1 _397_ (.A0(net10),
    .A1(net83),
    .S(net260),
    .Y(_195_));
 sky130_fd_sc_hd__nand2_1 _398_ (.A(net186),
    .B(net256),
    .Y(_196_));
 sky130_fd_sc_hd__o21ai_1 _399_ (.A1(net256),
    .A2(_195_),
    .B1(_196_),
    .Y(_061_));
 sky130_fd_sc_hd__mux2i_1 _400_ (.A0(net11),
    .A1(net84),
    .S(net260),
    .Y(_197_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input10 (.A(read_addr[17]),
    .X(net9));
 sky130_fd_sc_hd__nand2_1 _402_ (.A(net187),
    .B(net256),
    .Y(_199_));
 sky130_fd_sc_hd__o21ai_1 _403_ (.A1(net256),
    .A2(_197_),
    .B1(_199_),
    .Y(_062_));
 sky130_fd_sc_hd__mux2i_1 _404_ (.A0(net12),
    .A1(net85),
    .S(net260),
    .Y(_200_));
 sky130_fd_sc_hd__nand2_1 _405_ (.A(net188),
    .B(net256),
    .Y(_201_));
 sky130_fd_sc_hd__o21ai_1 _406_ (.A1(net256),
    .A2(_200_),
    .B1(_201_),
    .Y(_063_));
 sky130_fd_sc_hd__mux2i_1 _407_ (.A0(net13),
    .A1(net86),
    .S(net260),
    .Y(_202_));
 sky130_fd_sc_hd__nand2_1 _408_ (.A(net189),
    .B(net256),
    .Y(_203_));
 sky130_fd_sc_hd__o21ai_0 _409_ (.A1(net256),
    .A2(_202_),
    .B1(_203_),
    .Y(_064_));
 sky130_fd_sc_hd__mux2i_1 _410_ (.A0(net14),
    .A1(net87),
    .S(net260),
    .Y(_204_));
 sky130_fd_sc_hd__nand2_1 _411_ (.A(net190),
    .B(net256),
    .Y(_205_));
 sky130_fd_sc_hd__o21ai_0 _412_ (.A1(net256),
    .A2(_204_),
    .B1(_205_),
    .Y(_065_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input9 (.A(read_addr[16]),
    .X(net8));
 sky130_fd_sc_hd__mux2i_1 _414_ (.A0(net15),
    .A1(net88),
    .S(net260),
    .Y(_207_));
 sky130_fd_sc_hd__nand2_1 _415_ (.A(net191),
    .B(net256),
    .Y(_208_));
 sky130_fd_sc_hd__o21ai_1 _416_ (.A1(net256),
    .A2(_207_),
    .B1(_208_),
    .Y(_066_));
 sky130_fd_sc_hd__mux2i_1 _417_ (.A0(net16),
    .A1(net89),
    .S(net260),
    .Y(_209_));
 sky130_fd_sc_hd__nand2_1 _418_ (.A(net192),
    .B(net256),
    .Y(_210_));
 sky130_fd_sc_hd__o21ai_0 _419_ (.A1(net256),
    .A2(_209_),
    .B1(_210_),
    .Y(_067_));
 sky130_fd_sc_hd__mux2i_1 _420_ (.A0(net17),
    .A1(net90),
    .S(net260),
    .Y(_211_));
 sky130_fd_sc_hd__nand2_1 _421_ (.A(net193),
    .B(net256),
    .Y(_212_));
 sky130_fd_sc_hd__o21ai_1 _422_ (.A1(net256),
    .A2(_211_),
    .B1(_212_),
    .Y(_068_));
 sky130_fd_sc_hd__mux2i_1 _423_ (.A0(net18),
    .A1(net91),
    .S(net260),
    .Y(_213_));
 sky130_fd_sc_hd__nand2_1 _424_ (.A(net194),
    .B(net256),
    .Y(_214_));
 sky130_fd_sc_hd__o21ai_0 _425_ (.A1(net256),
    .A2(_213_),
    .B1(_214_),
    .Y(_069_));
 sky130_fd_sc_hd__mux2i_1 _426_ (.A0(net19),
    .A1(net92),
    .S(net260),
    .Y(_215_));
 sky130_fd_sc_hd__nand2_1 _427_ (.A(net195),
    .B(net256),
    .Y(_216_));
 sky130_fd_sc_hd__o21ai_1 _428_ (.A1(net256),
    .A2(_215_),
    .B1(_216_),
    .Y(_070_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input8 (.A(read_addr[15]),
    .X(net7));
 sky130_fd_sc_hd__mux2i_1 _430_ (.A0(net20),
    .A1(net93),
    .S(net260),
    .Y(_218_));
 sky130_fd_sc_hd__nand2_1 _431_ (.A(net196),
    .B(net256),
    .Y(_219_));
 sky130_fd_sc_hd__o21ai_0 _432_ (.A1(net256),
    .A2(_218_),
    .B1(_219_),
    .Y(_071_));
 sky130_fd_sc_hd__mux2i_1 _433_ (.A0(net21),
    .A1(net94),
    .S(net260),
    .Y(_220_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input7 (.A(read_addr[14]),
    .X(net6));
 sky130_fd_sc_hd__nand2_1 _435_ (.A(net197),
    .B(net256),
    .Y(_222_));
 sky130_fd_sc_hd__o21ai_0 _436_ (.A1(net256),
    .A2(_220_),
    .B1(_222_),
    .Y(_072_));
 sky130_fd_sc_hd__mux2i_1 _437_ (.A0(net22),
    .A1(net95),
    .S(net260),
    .Y(_223_));
 sky130_fd_sc_hd__nand2_1 _438_ (.A(net198),
    .B(net256),
    .Y(_224_));
 sky130_fd_sc_hd__o21ai_0 _439_ (.A1(net256),
    .A2(_223_),
    .B1(_224_),
    .Y(_073_));
 sky130_fd_sc_hd__mux2i_1 _440_ (.A0(net23),
    .A1(net96),
    .S(net260),
    .Y(_225_));
 sky130_fd_sc_hd__nand2_1 _441_ (.A(net199),
    .B(net256),
    .Y(_226_));
 sky130_fd_sc_hd__o21ai_0 _442_ (.A1(net256),
    .A2(_225_),
    .B1(_226_),
    .Y(_074_));
 sky130_fd_sc_hd__mux2i_1 _443_ (.A0(net24),
    .A1(net97),
    .S(net260),
    .Y(_227_));
 sky130_fd_sc_hd__nand2_1 _444_ (.A(net200),
    .B(net256),
    .Y(_228_));
 sky130_fd_sc_hd__o21ai_0 _445_ (.A1(net256),
    .A2(_227_),
    .B1(_228_),
    .Y(_075_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input6 (.A(read_addr[13]),
    .X(net5));
 sky130_fd_sc_hd__mux2i_1 _447_ (.A0(net25),
    .A1(net98),
    .S(net260),
    .Y(_230_));
 sky130_fd_sc_hd__nand2_1 _448_ (.A(net201),
    .B(net256),
    .Y(_231_));
 sky130_fd_sc_hd__o21ai_0 _449_ (.A1(net256),
    .A2(_230_),
    .B1(_231_),
    .Y(_076_));
 sky130_fd_sc_hd__mux2i_1 _450_ (.A0(net26),
    .A1(net99),
    .S(net260),
    .Y(_232_));
 sky130_fd_sc_hd__nand2_1 _451_ (.A(net202),
    .B(net256),
    .Y(_233_));
 sky130_fd_sc_hd__o21ai_0 _452_ (.A1(net256),
    .A2(_232_),
    .B1(_233_),
    .Y(_077_));
 sky130_fd_sc_hd__mux2i_1 _453_ (.A0(net27),
    .A1(net100),
    .S(net260),
    .Y(_234_));
 sky130_fd_sc_hd__nand2_1 _454_ (.A(net203),
    .B(net256),
    .Y(_235_));
 sky130_fd_sc_hd__o21ai_0 _455_ (.A1(net256),
    .A2(_234_),
    .B1(_235_),
    .Y(_078_));
 sky130_fd_sc_hd__mux2i_1 _456_ (.A0(net28),
    .A1(net101),
    .S(net260),
    .Y(_236_));
 sky130_fd_sc_hd__nand2_1 _457_ (.A(net204),
    .B(net256),
    .Y(_237_));
 sky130_fd_sc_hd__o21ai_0 _458_ (.A1(net256),
    .A2(_236_),
    .B1(_237_),
    .Y(_079_));
 sky130_fd_sc_hd__mux2i_1 _459_ (.A0(net29),
    .A1(net102),
    .S(net260),
    .Y(_238_));
 sky130_fd_sc_hd__nand2_1 _460_ (.A(net205),
    .B(net256),
    .Y(_239_));
 sky130_fd_sc_hd__o21ai_0 _461_ (.A1(net256),
    .A2(_238_),
    .B1(_239_),
    .Y(_080_));
 sky130_fd_sc_hd__mux2i_1 _462_ (.A0(net30),
    .A1(net103),
    .S(net260),
    .Y(_240_));
 sky130_fd_sc_hd__nand2_1 _463_ (.A(net206),
    .B(net256),
    .Y(_241_));
 sky130_fd_sc_hd__o21ai_0 _464_ (.A1(net256),
    .A2(_240_),
    .B1(_241_),
    .Y(_081_));
 sky130_fd_sc_hd__mux2i_1 _465_ (.A0(net31),
    .A1(net104),
    .S(net260),
    .Y(_242_));
 sky130_fd_sc_hd__nand2_1 _466_ (.A(net207),
    .B(net256),
    .Y(_243_));
 sky130_fd_sc_hd__o21ai_0 _467_ (.A1(net256),
    .A2(_242_),
    .B1(_243_),
    .Y(_082_));
 sky130_fd_sc_hd__mux2i_1 _468_ (.A0(net32),
    .A1(net105),
    .S(net260),
    .Y(_244_));
 sky130_fd_sc_hd__nand2_1 _469_ (.A(net208),
    .B(net256),
    .Y(_245_));
 sky130_fd_sc_hd__o21ai_0 _470_ (.A1(net256),
    .A2(_244_),
    .B1(_245_),
    .Y(_083_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input5 (.A(read_addr[12]),
    .X(net4));
 sky130_fd_sc_hd__mux2_4 _472_ (.A0(net106),
    .A1(net210),
    .S(net257),
    .X(_084_));
 sky130_fd_sc_hd__mux2_4 _473_ (.A0(net107),
    .A1(net211),
    .S(net257),
    .X(_085_));
 sky130_fd_sc_hd__mux2_4 _474_ (.A0(net108),
    .A1(net212),
    .S(net257),
    .X(_086_));
 sky130_fd_sc_hd__mux2_4 _475_ (.A0(net109),
    .A1(net213),
    .S(net257),
    .X(_087_));
 sky130_fd_sc_hd__mux2_4 _476_ (.A0(net110),
    .A1(net214),
    .S(net257),
    .X(_088_));
 sky130_fd_sc_hd__mux2_4 _477_ (.A0(net111),
    .A1(net215),
    .S(net257),
    .X(_089_));
 sky130_fd_sc_hd__mux2_4 _478_ (.A0(net112),
    .A1(net216),
    .S(net257),
    .X(_090_));
 sky130_fd_sc_hd__mux2_4 _479_ (.A0(net113),
    .A1(net217),
    .S(net257),
    .X(_091_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input4 (.A(read_addr[11]),
    .X(net3));
 sky130_fd_sc_hd__mux2_4 _481_ (.A0(net114),
    .A1(net218),
    .S(net257),
    .X(_092_));
 sky130_fd_sc_hd__mux2_4 _482_ (.A0(net115),
    .A1(net219),
    .S(net257),
    .X(_093_));
 sky130_fd_sc_hd__mux2_4 _483_ (.A0(net116),
    .A1(net220),
    .S(net257),
    .X(_094_));
 sky130_fd_sc_hd__mux2_4 _484_ (.A0(net117),
    .A1(net221),
    .S(net257),
    .X(_095_));
 sky130_fd_sc_hd__mux2_4 _485_ (.A0(net118),
    .A1(net222),
    .S(net257),
    .X(_096_));
 sky130_fd_sc_hd__mux2_4 _486_ (.A0(net119),
    .A1(net223),
    .S(net257),
    .X(_097_));
 sky130_fd_sc_hd__mux2_4 _487_ (.A0(net120),
    .A1(net224),
    .S(net257),
    .X(_098_));
 sky130_fd_sc_hd__mux2_4 _488_ (.A0(net121),
    .A1(net225),
    .S(net257),
    .X(_099_));
 sky130_fd_sc_hd__mux2_4 _489_ (.A0(net122),
    .A1(net226),
    .S(net257),
    .X(_100_));
 sky130_fd_sc_hd__mux2_4 _490_ (.A0(net123),
    .A1(net227),
    .S(net257),
    .X(_101_));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input3 (.A(read_addr[10]),
    .X(net2));
 sky130_fd_sc_hd__mux2_4 _492_ (.A0(net124),
    .A1(net228),
    .S(net257),
    .X(_102_));
 sky130_fd_sc_hd__mux2_4 _493_ (.A0(net125),
    .A1(net229),
    .S(net257),
    .X(_103_));
 sky130_fd_sc_hd__mux2_4 _494_ (.A0(net126),
    .A1(net230),
    .S(net257),
    .X(_104_));
 sky130_fd_sc_hd__mux2_4 _495_ (.A0(net127),
    .A1(net231),
    .S(net257),
    .X(_105_));
 sky130_fd_sc_hd__mux2_4 _496_ (.A0(net128),
    .A1(net232),
    .S(net257),
    .X(_106_));
 sky130_fd_sc_hd__mux2_4 _497_ (.A0(net129),
    .A1(net233),
    .S(net257),
    .X(_107_));
 sky130_fd_sc_hd__mux2_4 _498_ (.A0(net130),
    .A1(net234),
    .S(net257),
    .X(_108_));
 sky130_fd_sc_hd__mux2_4 _499_ (.A0(net131),
    .A1(net235),
    .S(net257),
    .X(_109_));
 sky130_fd_sc_hd__mux2_4 _500_ (.A0(net132),
    .A1(net236),
    .S(net257),
    .X(_110_));
 sky130_fd_sc_hd__mux2_4 _501_ (.A0(net133),
    .A1(net237),
    .S(net257),
    .X(_111_));
 sky130_fd_sc_hd__mux2_2 _502_ (.A0(net134),
    .A1(net238),
    .S(net257),
    .X(_112_));
 sky130_fd_sc_hd__mux2_2 _503_ (.A0(net135),
    .A1(net239),
    .S(net257),
    .X(_113_));
 sky130_fd_sc_hd__mux2_2 _504_ (.A0(net136),
    .A1(net240),
    .S(net257),
    .X(_114_));
 sky130_fd_sc_hd__mux2_2 _505_ (.A0(net137),
    .A1(net241),
    .S(net257),
    .X(_115_));
 sky130_fd_sc_hd__mux2i_1 _506_ (.A0(net34),
    .A1(net139),
    .S(net260),
    .Y(_249_));
 sky130_fd_sc_hd__nand2_1 _507_ (.A(net242),
    .B(net256),
    .Y(_250_));
 sky130_fd_sc_hd__o21ai_0 _508_ (.A1(net256),
    .A2(_249_),
    .B1(_250_),
    .Y(_116_));
 sky130_fd_sc_hd__mux2i_1 _509_ (.A0(net35),
    .A1(net140),
    .S(net260),
    .Y(_251_));
 sky130_fd_sc_hd__nand2_1 _510_ (.A(net243),
    .B(net256),
    .Y(_252_));
 sky130_fd_sc_hd__o21ai_0 _511_ (.A1(net256),
    .A2(_251_),
    .B1(_252_),
    .Y(_117_));
 sky130_fd_sc_hd__mux2i_1 _512_ (.A0(net36),
    .A1(net141),
    .S(net260),
    .Y(_253_));
 sky130_fd_sc_hd__nand2_1 _513_ (.A(net244),
    .B(net256),
    .Y(_254_));
 sky130_fd_sc_hd__o21ai_0 _514_ (.A1(net256),
    .A2(_253_),
    .B1(_254_),
    .Y(_118_));
 sky130_fd_sc_hd__mux2i_1 _515_ (.A0(net37),
    .A1(net142),
    .S(net260),
    .Y(_255_));
 sky130_fd_sc_hd__nand2_1 _516_ (.A(net245),
    .B(net256),
    .Y(_256_));
 sky130_fd_sc_hd__o21ai_0 _517_ (.A1(net256),
    .A2(_255_),
    .B1(_256_),
    .Y(_119_));
 sky130_fd_sc_hd__and2_1 _518_ (.A(net33),
    .B(_002_),
    .X(_257_));
 sky130_fd_sc_hd__o21ai_0 _519_ (.A1(_166_),
    .A2(_257_),
    .B1(net257),
    .Y(_120_));
 sky130_fd_sc_hd__mux2i_1 _520_ (.A0(net248),
    .A1(_005_),
    .S(net260),
    .Y(_258_));
 sky130_fd_sc_hd__a21oi_1 _521_ (.A1(net39),
    .A2(_005_),
    .B1(net248),
    .Y(_259_));
 sky130_fd_sc_hd__a21oi_1 _522_ (.A1(_002_),
    .A2(_258_),
    .B1(_259_),
    .Y(_121_));
 sky130_fd_sc_hd__nand2_1 _523_ (.A(\retry_count[3] ),
    .B(net247),
    .Y(_260_));
 sky130_fd_sc_hd__nand2b_1 _524_ (.A_N(net39),
    .B(net72),
    .Y(_261_));
 sky130_fd_sc_hd__a221oi_2 _525_ (.A1(_006_),
    .A2(_260_),
    .B1(_261_),
    .B2(_005_),
    .C1(_163_),
    .Y(_262_));
 sky130_fd_sc_hd__nor2_1 _526_ (.A(net249),
    .B(_262_),
    .Y(_263_));
 sky130_fd_sc_hd__a211oi_1 _527_ (.A1(net249),
    .A2(net257),
    .B1(_006_),
    .C1(_005_),
    .Y(_264_));
 sky130_fd_sc_hd__nor2_1 _528_ (.A(_263_),
    .B(_264_),
    .Y(_122_));
 sky130_fd_sc_hd__ha_1 _529_ (.A(_000_),
    .B(_001_),
    .COUT(_002_),
    .SUM(_003_));
 sky130_fd_sc_hd__ha_1 _530_ (.A(_000_),
    .B(\state[1] ),
    .COUT(_004_),
    .SUM(_266_));
 sky130_fd_sc_hd__ha_1 _531_ (.A(\state[0] ),
    .B(_001_),
    .COUT(_005_),
    .SUM(_267_));
 sky130_fd_sc_hd__ha_1 _532_ (.A(\state[0] ),
    .B(\state[1] ),
    .COUT(_006_),
    .SUM(_268_));
 sky130_fd_sc_hd__ha_1 _533_ (.A(_007_),
    .B(_008_),
    .COUT(_009_),
    .SUM(_010_));
 sky130_fd_sc_hd__ha_1 _534_ (.A(\retry_count[0] ),
    .B(\retry_count[1] ),
    .COUT(_011_),
    .SUM(_269_));
 sky130_fd_sc_hd__buf_4 place261 (.A(net138),
    .X(net260));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input2 (.A(read_addr[0]),
    .X(net1));
 sky130_fd_sc_hd__dfrtp_1 \read_data[0]$_DFFE_PN0P_  (.D(_012_),
    .Q(net143),
    .RESET_B(net258),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[10]$_DFFE_PN0P_  (.D(_013_),
    .Q(net144),
    .RESET_B(net258),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[11]$_DFFE_PN0P_  (.D(_014_),
    .Q(net145),
    .RESET_B(net259),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[12]$_DFFE_PN0P_  (.D(_015_),
    .Q(net146),
    .RESET_B(net259),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[13]$_DFFE_PN0P_  (.D(_016_),
    .Q(net147),
    .RESET_B(net258),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[14]$_DFFE_PN0P_  (.D(_017_),
    .Q(net148),
    .RESET_B(net259),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[15]$_DFFE_PN0P_  (.D(_018_),
    .Q(net149),
    .RESET_B(net259),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[16]$_DFFE_PN0P_  (.D(_019_),
    .Q(net150),
    .RESET_B(net258),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[17]$_DFFE_PN0P_  (.D(_020_),
    .Q(net151),
    .RESET_B(net38),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[18]$_DFFE_PN0P_  (.D(_021_),
    .Q(net152),
    .RESET_B(net38),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[19]$_DFFE_PN0P_  (.D(_022_),
    .Q(net153),
    .RESET_B(net38),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[1]$_DFFE_PN0P_  (.D(_023_),
    .Q(net154),
    .RESET_B(net38),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[20]$_DFFE_PN0P_  (.D(_024_),
    .Q(net155),
    .RESET_B(net38),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[21]$_DFFE_PN0P_  (.D(_025_),
    .Q(net156),
    .RESET_B(net38),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[22]$_DFFE_PN0P_  (.D(_026_),
    .Q(net157),
    .RESET_B(net38),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[23]$_DFFE_PN0P_  (.D(_027_),
    .Q(net158),
    .RESET_B(net38),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[24]$_DFFE_PN0P_  (.D(_028_),
    .Q(net159),
    .RESET_B(net38),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[25]$_DFFE_PN0P_  (.D(_029_),
    .Q(net160),
    .RESET_B(net38),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[26]$_DFFE_PN0P_  (.D(_030_),
    .Q(net161),
    .RESET_B(net38),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[27]$_DFFE_PN0P_  (.D(_031_),
    .Q(net162),
    .RESET_B(net38),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[28]$_DFFE_PN0P_  (.D(_032_),
    .Q(net163),
    .RESET_B(net38),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[29]$_DFFE_PN0P_  (.D(_033_),
    .Q(net164),
    .RESET_B(net38),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[2]$_DFFE_PN0P_  (.D(_034_),
    .Q(net165),
    .RESET_B(net38),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[30]$_DFFE_PN0P_  (.D(_035_),
    .Q(net166),
    .RESET_B(net38),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[31]$_DFFE_PN0P_  (.D(_036_),
    .Q(net167),
    .RESET_B(net38),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[3]$_DFFE_PN0P_  (.D(_037_),
    .Q(net168),
    .RESET_B(net38),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[4]$_DFFE_PN0P_  (.D(_038_),
    .Q(net169),
    .RESET_B(net38),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[5]$_DFFE_PN0P_  (.D(_039_),
    .Q(net170),
    .RESET_B(net38),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[6]$_DFFE_PN0P_  (.D(_040_),
    .Q(net171),
    .RESET_B(net258),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[7]$_DFFE_PN0P_  (.D(_041_),
    .Q(net172),
    .RESET_B(net258),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[8]$_DFFE_PN0P_  (.D(_042_),
    .Q(net173),
    .RESET_B(net258),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[9]$_DFFE_PN0P_  (.D(_043_),
    .Q(net174),
    .RESET_B(net258),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_done$_DFFE_PN0P_  (.D(_044_),
    .Q(net175),
    .RESET_B(net258),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_err$_DFFE_PN0P_  (.D(_045_),
    .Q(net176),
    .RESET_B(net258),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \retry_count[0]$_DFFE_PN0P_  (.D(_046_),
    .Q(\retry_count[0] ),
    .RESET_B(net258),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \retry_count[1]$_DFFE_PN0P_  (.D(_047_),
    .Q(\retry_count[1] ),
    .RESET_B(net258),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \retry_count[2]$_DFFE_PN0P_  (.D(_048_),
    .Q(\retry_count[2] ),
    .RESET_B(net258),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \retry_count[3]$_DFFE_PN0P_  (.D(_049_),
    .Q(\retry_count[3] ),
    .RESET_B(net258),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \state[0]$_DFFE_PN0P_  (.D(_050_),
    .Q(\state[0] ),
    .RESET_B(net258),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \state[1]$_DFFE_PN0P_  (.D(_051_),
    .Q(\state[1] ),
    .RESET_B(net258),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[0]$_DFFE_PN0P_  (.D(_052_),
    .Q(net177),
    .RESET_B(net259),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[10]$_DFFE_PN0P_  (.D(_053_),
    .Q(net178),
    .RESET_B(net259),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[11]$_DFFE_PN0P_  (.D(_054_),
    .Q(net179),
    .RESET_B(net259),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[12]$_DFFE_PN0P_  (.D(_055_),
    .Q(net180),
    .RESET_B(net259),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[13]$_DFFE_PN0P_  (.D(_056_),
    .Q(net181),
    .RESET_B(net259),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[14]$_DFFE_PN0P_  (.D(_057_),
    .Q(net182),
    .RESET_B(net259),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[15]$_DFFE_PN0P_  (.D(_058_),
    .Q(net183),
    .RESET_B(net259),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[16]$_DFFE_PN0P_  (.D(_059_),
    .Q(net184),
    .RESET_B(net259),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[17]$_DFFE_PN0P_  (.D(_060_),
    .Q(net185),
    .RESET_B(net259),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[18]$_DFFE_PN0P_  (.D(_061_),
    .Q(net186),
    .RESET_B(net259),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[19]$_DFFE_PN0P_  (.D(_062_),
    .Q(net187),
    .RESET_B(net259),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[1]$_DFFE_PN0P_  (.D(_063_),
    .Q(net188),
    .RESET_B(net259),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[20]$_DFFE_PN0P_  (.D(_064_),
    .Q(net189),
    .RESET_B(net259),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[21]$_DFFE_PN0P_  (.D(_065_),
    .Q(net190),
    .RESET_B(net259),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[22]$_DFFE_PN0P_  (.D(_066_),
    .Q(net191),
    .RESET_B(net259),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[23]$_DFFE_PN0P_  (.D(_067_),
    .Q(net192),
    .RESET_B(net259),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[24]$_DFFE_PN0P_  (.D(_068_),
    .Q(net193),
    .RESET_B(net259),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[25]$_DFFE_PN0P_  (.D(_069_),
    .Q(net194),
    .RESET_B(net259),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[26]$_DFFE_PN0P_  (.D(_070_),
    .Q(net195),
    .RESET_B(net259),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[27]$_DFFE_PN0P_  (.D(_071_),
    .Q(net196),
    .RESET_B(net259),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[28]$_DFFE_PN0P_  (.D(_072_),
    .Q(net197),
    .RESET_B(net259),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[29]$_DFFE_PN0P_  (.D(_073_),
    .Q(net198),
    .RESET_B(net259),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[2]$_DFFE_PN0P_  (.D(_074_),
    .Q(net199),
    .RESET_B(net259),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[30]$_DFFE_PN0P_  (.D(_075_),
    .Q(net200),
    .RESET_B(net259),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[31]$_DFFE_PN0P_  (.D(_076_),
    .Q(net201),
    .RESET_B(net259),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[3]$_DFFE_PN0P_  (.D(_077_),
    .Q(net202),
    .RESET_B(net259),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[4]$_DFFE_PN0P_  (.D(_078_),
    .Q(net203),
    .RESET_B(net259),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[5]$_DFFE_PN0P_  (.D(_079_),
    .Q(net204),
    .RESET_B(net259),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[6]$_DFFE_PN0P_  (.D(_080_),
    .Q(net205),
    .RESET_B(net259),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[7]$_DFFE_PN0P_  (.D(_081_),
    .Q(net206),
    .RESET_B(net259),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[8]$_DFFE_PN0P_  (.D(_082_),
    .Q(net207),
    .RESET_B(net259),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[9]$_DFFE_PN0P_  (.D(_083_),
    .Q(net208),
    .RESET_B(net259),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[0]$_DFFE_PN0P_  (.D(_084_),
    .Q(net210),
    .RESET_B(net38),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[10]$_DFFE_PN0P_  (.D(_085_),
    .Q(net211),
    .RESET_B(net258),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[11]$_DFFE_PN0P_  (.D(_086_),
    .Q(net212),
    .RESET_B(net258),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[12]$_DFFE_PN0P_  (.D(_087_),
    .Q(net213),
    .RESET_B(net258),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[13]$_DFFE_PN0P_  (.D(_088_),
    .Q(net214),
    .RESET_B(net258),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[14]$_DFFE_PN0P_  (.D(_089_),
    .Q(net215),
    .RESET_B(net258),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[15]$_DFFE_PN0P_  (.D(_090_),
    .Q(net216),
    .RESET_B(net258),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[16]$_DFFE_PN0P_  (.D(_091_),
    .Q(net217),
    .RESET_B(net258),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[17]$_DFFE_PN0P_  (.D(_092_),
    .Q(net218),
    .RESET_B(net38),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[18]$_DFFE_PN0P_  (.D(_093_),
    .Q(net219),
    .RESET_B(net38),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[19]$_DFFE_PN0P_  (.D(_094_),
    .Q(net220),
    .RESET_B(net38),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[1]$_DFFE_PN0P_  (.D(_095_),
    .Q(net221),
    .RESET_B(net259),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[20]$_DFFE_PN0P_  (.D(_096_),
    .Q(net222),
    .RESET_B(net259),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[21]$_DFFE_PN0P_  (.D(_097_),
    .Q(net223),
    .RESET_B(net259),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[22]$_DFFE_PN0P_  (.D(_098_),
    .Q(net224),
    .RESET_B(net38),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[23]$_DFFE_PN0P_  (.D(_099_),
    .Q(net225),
    .RESET_B(net259),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[24]$_DFFE_PN0P_  (.D(_100_),
    .Q(net226),
    .RESET_B(net38),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[25]$_DFFE_PN0P_  (.D(_101_),
    .Q(net227),
    .RESET_B(net38),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[26]$_DFFE_PN0P_  (.D(_102_),
    .Q(net228),
    .RESET_B(net258),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[27]$_DFFE_PN0P_  (.D(_103_),
    .Q(net229),
    .RESET_B(net258),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[28]$_DFFE_PN0P_  (.D(_104_),
    .Q(net230),
    .RESET_B(net38),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[29]$_DFFE_PN0P_  (.D(_105_),
    .Q(net231),
    .RESET_B(net38),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[2]$_DFFE_PN0P_  (.D(_106_),
    .Q(net232),
    .RESET_B(net258),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[30]$_DFFE_PN0P_  (.D(_107_),
    .Q(net233),
    .RESET_B(net258),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[31]$_DFFE_PN0P_  (.D(_108_),
    .Q(net234),
    .RESET_B(net258),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[3]$_DFFE_PN0P_  (.D(_109_),
    .Q(net235),
    .RESET_B(net258),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[4]$_DFFE_PN0P_  (.D(_110_),
    .Q(net236),
    .RESET_B(net38),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[5]$_DFFE_PN0P_  (.D(_111_),
    .Q(net237),
    .RESET_B(net258),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[6]$_DFFE_PN0P_  (.D(_112_),
    .Q(net238),
    .RESET_B(net38),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[7]$_DFFE_PN0P_  (.D(_113_),
    .Q(net239),
    .RESET_B(net38),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[8]$_DFFE_PN0P_  (.D(_114_),
    .Q(net240),
    .RESET_B(net38),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[9]$_DFFE_PN0P_  (.D(_115_),
    .Q(net241),
    .RESET_B(net38),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_sel_o[0]$_DFFE_PN0P_  (.D(_116_),
    .Q(net242),
    .RESET_B(net259),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_sel_o[1]$_DFFE_PN0P_  (.D(_117_),
    .Q(net243),
    .RESET_B(net259),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_sel_o[2]$_DFFE_PN0P_  (.D(_118_),
    .Q(net244),
    .RESET_B(net259),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_sel_o[3]$_DFFE_PN0P_  (.D(_119_),
    .Q(net245),
    .RESET_B(net259),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_stb_o$_DFF_PN0_  (.D(_265_),
    .Q(net209),
    .RESET_B(net259),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_we_o$_DFFE_PN0P_  (.D(_120_),
    .Q(net247),
    .RESET_B(net258),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \write_done$_DFFE_PN0P_  (.D(_121_),
    .Q(net248),
    .RESET_B(net258),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \write_err$_DFFE_PN0P_  (.D(_122_),
    .Q(net249),
    .RESET_B(net258),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__conb_1 _537__1 (.LO(wb_tgd_o[0]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input25 (.A(read_addr[30]),
    .X(net24));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input26 (.A(read_addr[31]),
    .X(net25));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input27 (.A(read_addr[3]),
    .X(net26));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input28 (.A(read_addr[4]),
    .X(net27));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input29 (.A(read_addr[5]),
    .X(net28));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input30 (.A(read_addr[6]),
    .X(net29));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input31 (.A(read_addr[7]),
    .X(net30));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input32 (.A(read_addr[8]),
    .X(net31));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input33 (.A(read_addr[9]),
    .X(net32));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input34 (.A(read_req),
    .X(net33));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input35 (.A(read_sel[0]),
    .X(net34));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input36 (.A(read_sel[1]),
    .X(net35));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input37 (.A(read_sel[2]),
    .X(net36));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input38 (.A(read_sel[3]),
    .X(net37));
 sky130_fd_sc_hd__buf_4 input39 (.A(net261),
    .X(net38));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input40 (.A(wb_ack_i),
    .X(net39));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input41 (.A(wb_dat_i[0]),
    .X(net40));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input42 (.A(wb_dat_i[10]),
    .X(net41));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input43 (.A(wb_dat_i[11]),
    .X(net42));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input44 (.A(wb_dat_i[12]),
    .X(net43));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input45 (.A(wb_dat_i[13]),
    .X(net44));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input46 (.A(wb_dat_i[14]),
    .X(net45));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input47 (.A(wb_dat_i[15]),
    .X(net46));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input48 (.A(wb_dat_i[16]),
    .X(net47));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input49 (.A(wb_dat_i[17]),
    .X(net48));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input50 (.A(wb_dat_i[18]),
    .X(net49));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input51 (.A(wb_dat_i[19]),
    .X(net50));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input52 (.A(wb_dat_i[1]),
    .X(net51));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input53 (.A(wb_dat_i[20]),
    .X(net52));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input54 (.A(wb_dat_i[21]),
    .X(net53));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input55 (.A(wb_dat_i[22]),
    .X(net54));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input56 (.A(wb_dat_i[23]),
    .X(net55));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input57 (.A(wb_dat_i[24]),
    .X(net56));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input58 (.A(wb_dat_i[25]),
    .X(net57));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input59 (.A(wb_dat_i[26]),
    .X(net58));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input60 (.A(wb_dat_i[27]),
    .X(net59));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input61 (.A(wb_dat_i[28]),
    .X(net60));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input62 (.A(wb_dat_i[29]),
    .X(net61));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input63 (.A(wb_dat_i[2]),
    .X(net62));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input64 (.A(wb_dat_i[30]),
    .X(net63));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input65 (.A(wb_dat_i[31]),
    .X(net64));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input66 (.A(wb_dat_i[3]),
    .X(net65));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input67 (.A(wb_dat_i[4]),
    .X(net66));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input68 (.A(wb_dat_i[5]),
    .X(net67));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input69 (.A(wb_dat_i[6]),
    .X(net68));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input70 (.A(wb_dat_i[7]),
    .X(net69));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input71 (.A(wb_dat_i[8]),
    .X(net70));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input72 (.A(wb_dat_i[9]),
    .X(net71));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input73 (.A(wb_err_i),
    .X(net72));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input74 (.A(wb_rty_i),
    .X(net73));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input75 (.A(write_addr[0]),
    .X(net74));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input76 (.A(write_addr[10]),
    .X(net75));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input77 (.A(write_addr[11]),
    .X(net76));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input78 (.A(write_addr[12]),
    .X(net77));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input79 (.A(write_addr[13]),
    .X(net78));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input80 (.A(write_addr[14]),
    .X(net79));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input81 (.A(write_addr[15]),
    .X(net80));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input82 (.A(write_addr[16]),
    .X(net81));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input83 (.A(write_addr[17]),
    .X(net82));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input84 (.A(write_addr[18]),
    .X(net83));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input85 (.A(write_addr[19]),
    .X(net84));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input86 (.A(write_addr[1]),
    .X(net85));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input87 (.A(write_addr[20]),
    .X(net86));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input88 (.A(write_addr[21]),
    .X(net87));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input89 (.A(write_addr[22]),
    .X(net88));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input90 (.A(write_addr[23]),
    .X(net89));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input91 (.A(write_addr[24]),
    .X(net90));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input92 (.A(write_addr[25]),
    .X(net91));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input93 (.A(write_addr[26]),
    .X(net92));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input94 (.A(write_addr[27]),
    .X(net93));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input95 (.A(write_addr[28]),
    .X(net94));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input96 (.A(write_addr[29]),
    .X(net95));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input97 (.A(write_addr[2]),
    .X(net96));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input98 (.A(write_addr[30]),
    .X(net97));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input99 (.A(write_addr[31]),
    .X(net98));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input100 (.A(write_addr[3]),
    .X(net99));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input101 (.A(write_addr[4]),
    .X(net100));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input102 (.A(write_addr[5]),
    .X(net101));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input103 (.A(write_addr[6]),
    .X(net102));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input104 (.A(write_addr[7]),
    .X(net103));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input105 (.A(write_addr[8]),
    .X(net104));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input106 (.A(write_addr[9]),
    .X(net105));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input107 (.A(write_data[0]),
    .X(net106));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input108 (.A(write_data[10]),
    .X(net107));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input109 (.A(write_data[11]),
    .X(net108));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input110 (.A(write_data[12]),
    .X(net109));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input111 (.A(write_data[13]),
    .X(net110));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input112 (.A(write_data[14]),
    .X(net111));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input113 (.A(write_data[15]),
    .X(net112));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input114 (.A(write_data[16]),
    .X(net113));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input115 (.A(write_data[17]),
    .X(net114));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input116 (.A(write_data[18]),
    .X(net115));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input117 (.A(write_data[19]),
    .X(net116));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input118 (.A(write_data[1]),
    .X(net117));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input119 (.A(write_data[20]),
    .X(net118));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input120 (.A(write_data[21]),
    .X(net119));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input121 (.A(write_data[22]),
    .X(net120));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input122 (.A(write_data[23]),
    .X(net121));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input123 (.A(write_data[24]),
    .X(net122));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input124 (.A(write_data[25]),
    .X(net123));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input125 (.A(write_data[26]),
    .X(net124));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input126 (.A(write_data[27]),
    .X(net125));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input127 (.A(write_data[28]),
    .X(net126));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input128 (.A(write_data[29]),
    .X(net127));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input129 (.A(write_data[2]),
    .X(net128));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input130 (.A(write_data[30]),
    .X(net129));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input131 (.A(write_data[31]),
    .X(net130));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input132 (.A(write_data[3]),
    .X(net131));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input133 (.A(write_data[4]),
    .X(net132));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input134 (.A(write_data[5]),
    .X(net133));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input135 (.A(write_data[6]),
    .X(net134));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input136 (.A(write_data[7]),
    .X(net135));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input137 (.A(write_data[8]),
    .X(net136));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input138 (.A(write_data[9]),
    .X(net137));
 sky130_fd_sc_hd__buf_2 input139 (.A(write_req),
    .X(net138));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input140 (.A(write_sel[0]),
    .X(net139));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input141 (.A(write_sel[1]),
    .X(net140));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input142 (.A(write_sel[2]),
    .X(net141));
 sky130_fd_sc_hd__clkdlybuf4s50_1 input143 (.A(write_sel[3]),
    .X(net142));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output144 (.A(net143),
    .X(read_data[0]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output145 (.A(net144),
    .X(read_data[10]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output146 (.A(net145),
    .X(read_data[11]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output147 (.A(net146),
    .X(read_data[12]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output148 (.A(net147),
    .X(read_data[13]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output149 (.A(net148),
    .X(read_data[14]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output150 (.A(net149),
    .X(read_data[15]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output151 (.A(net150),
    .X(read_data[16]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output152 (.A(net151),
    .X(read_data[17]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output153 (.A(net152),
    .X(read_data[18]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output154 (.A(net153),
    .X(read_data[19]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output155 (.A(net154),
    .X(read_data[1]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output156 (.A(net155),
    .X(read_data[20]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output157 (.A(net156),
    .X(read_data[21]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output158 (.A(net157),
    .X(read_data[22]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output159 (.A(net158),
    .X(read_data[23]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output160 (.A(net159),
    .X(read_data[24]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output161 (.A(net160),
    .X(read_data[25]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output162 (.A(net161),
    .X(read_data[26]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output163 (.A(net162),
    .X(read_data[27]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output164 (.A(net163),
    .X(read_data[28]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output165 (.A(net164),
    .X(read_data[29]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output166 (.A(net165),
    .X(read_data[2]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output167 (.A(net166),
    .X(read_data[30]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output168 (.A(net167),
    .X(read_data[31]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output169 (.A(net168),
    .X(read_data[3]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output170 (.A(net169),
    .X(read_data[4]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output171 (.A(net170),
    .X(read_data[5]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output172 (.A(net171),
    .X(read_data[6]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output173 (.A(net172),
    .X(read_data[7]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output174 (.A(net173),
    .X(read_data[8]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output175 (.A(net174),
    .X(read_data[9]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output176 (.A(net175),
    .X(read_done));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output177 (.A(net176),
    .X(read_err));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output178 (.A(net177),
    .X(wb_adr_o[0]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output179 (.A(net178),
    .X(wb_adr_o[10]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output180 (.A(net179),
    .X(wb_adr_o[11]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output181 (.A(net180),
    .X(wb_adr_o[12]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output182 (.A(net181),
    .X(wb_adr_o[13]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output183 (.A(net182),
    .X(wb_adr_o[14]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output184 (.A(net183),
    .X(wb_adr_o[15]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output185 (.A(net184),
    .X(wb_adr_o[16]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output186 (.A(net185),
    .X(wb_adr_o[17]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output187 (.A(net186),
    .X(wb_adr_o[18]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output188 (.A(net187),
    .X(wb_adr_o[19]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output189 (.A(net188),
    .X(wb_adr_o[1]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output190 (.A(net189),
    .X(wb_adr_o[20]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output191 (.A(net190),
    .X(wb_adr_o[21]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output192 (.A(net191),
    .X(wb_adr_o[22]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output193 (.A(net192),
    .X(wb_adr_o[23]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output194 (.A(net193),
    .X(wb_adr_o[24]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output195 (.A(net194),
    .X(wb_adr_o[25]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output196 (.A(net195),
    .X(wb_adr_o[26]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output197 (.A(net196),
    .X(wb_adr_o[27]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output198 (.A(net197),
    .X(wb_adr_o[28]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output199 (.A(net198),
    .X(wb_adr_o[29]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output200 (.A(net199),
    .X(wb_adr_o[2]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output201 (.A(net200),
    .X(wb_adr_o[30]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output202 (.A(net201),
    .X(wb_adr_o[31]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output203 (.A(net202),
    .X(wb_adr_o[3]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output204 (.A(net203),
    .X(wb_adr_o[4]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output205 (.A(net204),
    .X(wb_adr_o[5]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output206 (.A(net205),
    .X(wb_adr_o[6]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output207 (.A(net206),
    .X(wb_adr_o[7]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output208 (.A(net207),
    .X(wb_adr_o[8]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output209 (.A(net208),
    .X(wb_adr_o[9]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output210 (.A(net209),
    .X(wb_cyc_o));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output211 (.A(net210),
    .X(wb_dat_o[0]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output212 (.A(net211),
    .X(wb_dat_o[10]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output213 (.A(net212),
    .X(wb_dat_o[11]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output214 (.A(net213),
    .X(wb_dat_o[12]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output215 (.A(net214),
    .X(wb_dat_o[13]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output216 (.A(net215),
    .X(wb_dat_o[14]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output217 (.A(net216),
    .X(wb_dat_o[15]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output218 (.A(net217),
    .X(wb_dat_o[16]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output219 (.A(net218),
    .X(wb_dat_o[17]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output220 (.A(net219),
    .X(wb_dat_o[18]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output221 (.A(net220),
    .X(wb_dat_o[19]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output222 (.A(net221),
    .X(wb_dat_o[1]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output223 (.A(net222),
    .X(wb_dat_o[20]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output224 (.A(net223),
    .X(wb_dat_o[21]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output225 (.A(net224),
    .X(wb_dat_o[22]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output226 (.A(net225),
    .X(wb_dat_o[23]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output227 (.A(net226),
    .X(wb_dat_o[24]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output228 (.A(net227),
    .X(wb_dat_o[25]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output229 (.A(net228),
    .X(wb_dat_o[26]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output230 (.A(net229),
    .X(wb_dat_o[27]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output231 (.A(net230),
    .X(wb_dat_o[28]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output232 (.A(net231),
    .X(wb_dat_o[29]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output233 (.A(net232),
    .X(wb_dat_o[2]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output234 (.A(net233),
    .X(wb_dat_o[30]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output235 (.A(net234),
    .X(wb_dat_o[31]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output236 (.A(net235),
    .X(wb_dat_o[3]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output237 (.A(net236),
    .X(wb_dat_o[4]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output238 (.A(net237),
    .X(wb_dat_o[5]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output239 (.A(net238),
    .X(wb_dat_o[6]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output240 (.A(net239),
    .X(wb_dat_o[7]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output241 (.A(net240),
    .X(wb_dat_o[8]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output242 (.A(net241),
    .X(wb_dat_o[9]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output243 (.A(net242),
    .X(wb_sel_o[0]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output244 (.A(net243),
    .X(wb_sel_o[1]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output245 (.A(net244),
    .X(wb_sel_o[2]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output246 (.A(net245),
    .X(wb_sel_o[3]));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output247 (.A(net209),
    .X(wb_stb_o));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output248 (.A(net247),
    .X(wb_we_o));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output249 (.A(net248),
    .X(write_done));
 sky130_fd_sc_hd__clkdlybuf4s50_1 output250 (.A(net249),
    .X(write_err));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__buf_4 place257 (.A(_171_),
    .X(net256));
 sky130_fd_sc_hd__buf_4 place258 (.A(_168_),
    .X(net257));
 sky130_fd_sc_hd__buf_4 place259 (.A(net38),
    .X(net258));
 sky130_fd_sc_hd__buf_4 place260 (.A(net38),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkinv_4 clkload0 (.A(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload1 (.A(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkinv_2 clkload2 (.A(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__inv_8 clkload3 (.A(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkinv_4 clkload4 (.A(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkinv_4 clkload5 (.A(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload6 (.A(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(rst_n),
    .X(net261));
endmodule
