module true_random_generator (clk,
    data_valid,
    enable,
    entropy_low,
    read_next,
    rst_n,
    test_failed,
    random_data);
 input clk;
 output data_valid;
 input enable;
 output entropy_low;
 input read_next;
 input rst_n;
 output test_failed;
 output [31:0] random_data;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire \entropy_pool2[0] ;
 wire \entropy_pool2[10] ;
 wire \entropy_pool2[11] ;
 wire \entropy_pool2[12] ;
 wire \entropy_pool2[13] ;
 wire \entropy_pool2[14] ;
 wire \entropy_pool2[15] ;
 wire \entropy_pool2[16] ;
 wire \entropy_pool2[17] ;
 wire \entropy_pool2[18] ;
 wire \entropy_pool2[19] ;
 wire \entropy_pool2[1] ;
 wire \entropy_pool2[20] ;
 wire \entropy_pool2[21] ;
 wire \entropy_pool2[22] ;
 wire \entropy_pool2[23] ;
 wire \entropy_pool2[24] ;
 wire \entropy_pool2[25] ;
 wire \entropy_pool2[26] ;
 wire \entropy_pool2[27] ;
 wire \entropy_pool2[28] ;
 wire \entropy_pool2[29] ;
 wire \entropy_pool2[2] ;
 wire \entropy_pool2[30] ;
 wire \entropy_pool2[31] ;
 wire \entropy_pool2[3] ;
 wire \entropy_pool2[4] ;
 wire \entropy_pool2[5] ;
 wire \entropy_pool2[6] ;
 wire \entropy_pool2[7] ;
 wire \entropy_pool2[8] ;
 wire \entropy_pool2[9] ;
 wire \entropy_pool[0] ;
 wire \entropy_pool[10] ;
 wire \entropy_pool[11] ;
 wire \entropy_pool[12] ;
 wire \entropy_pool[13] ;
 wire \entropy_pool[14] ;
 wire \entropy_pool[15] ;
 wire \entropy_pool[16] ;
 wire \entropy_pool[17] ;
 wire \entropy_pool[18] ;
 wire \entropy_pool[19] ;
 wire \entropy_pool[1] ;
 wire \entropy_pool[20] ;
 wire \entropy_pool[21] ;
 wire \entropy_pool[22] ;
 wire \entropy_pool[23] ;
 wire \entropy_pool[24] ;
 wire \entropy_pool[25] ;
 wire \entropy_pool[26] ;
 wire \entropy_pool[27] ;
 wire \entropy_pool[28] ;
 wire \entropy_pool[29] ;
 wire \entropy_pool[2] ;
 wire \entropy_pool[30] ;
 wire \entropy_pool[31] ;
 wire \entropy_pool[3] ;
 wire \entropy_pool[4] ;
 wire \entropy_pool[5] ;
 wire \entropy_pool[6] ;
 wire \entropy_pool[7] ;
 wire \entropy_pool[8] ;
 wire \entropy_pool[9] ;
 wire \gen_ring_osc.init_osc ;
 wire \gen_ring_osc.inv_chain[1] ;
 wire \gen_ring_osc.toggle_sampling ;
 wire \health_counter[0] ;
 wire \health_counter[1] ;
 wire \health_counter[2] ;
 wire \health_counter[3] ;
 wire \health_counter[4] ;
 wire \health_counter[5] ;
 wire \health_counter[6] ;
 wire \health_counter[7] ;
 wire \lfsr_reg[0] ;
 wire \lfsr_reg[10] ;
 wire \lfsr_reg[11] ;
 wire \lfsr_reg[12] ;
 wire \lfsr_reg[13] ;
 wire \lfsr_reg[14] ;
 wire \lfsr_reg[15] ;
 wire \lfsr_reg[16] ;
 wire \lfsr_reg[17] ;
 wire \lfsr_reg[18] ;
 wire \lfsr_reg[19] ;
 wire \lfsr_reg[1] ;
 wire \lfsr_reg[20] ;
 wire \lfsr_reg[21] ;
 wire \lfsr_reg[22] ;
 wire \lfsr_reg[23] ;
 wire \lfsr_reg[24] ;
 wire \lfsr_reg[25] ;
 wire \lfsr_reg[26] ;
 wire \lfsr_reg[27] ;
 wire \lfsr_reg[28] ;
 wire \lfsr_reg[29] ;
 wire \lfsr_reg[2] ;
 wire \lfsr_reg[30] ;
 wire \lfsr_reg[31] ;
 wire \lfsr_reg[3] ;
 wire \lfsr_reg[4] ;
 wire \lfsr_reg[5] ;
 wire \lfsr_reg[6] ;
 wire \lfsr_reg[7] ;
 wire \lfsr_reg[8] ;
 wire \lfsr_reg[9] ;
 wire \mixed_output[0] ;
 wire \mixed_output[10] ;
 wire \mixed_output[11] ;
 wire \mixed_output[12] ;
 wire \mixed_output[13] ;
 wire \mixed_output[14] ;
 wire \mixed_output[15] ;
 wire \mixed_output[16] ;
 wire \mixed_output[17] ;
 wire \mixed_output[18] ;
 wire \mixed_output[19] ;
 wire \mixed_output[1] ;
 wire \mixed_output[20] ;
 wire \mixed_output[21] ;
 wire \mixed_output[22] ;
 wire \mixed_output[23] ;
 wire \mixed_output[24] ;
 wire \mixed_output[25] ;
 wire \mixed_output[26] ;
 wire \mixed_output[27] ;
 wire \mixed_output[28] ;
 wire \mixed_output[29] ;
 wire \mixed_output[2] ;
 wire \mixed_output[30] ;
 wire \mixed_output[31] ;
 wire \mixed_output[3] ;
 wire \mixed_output[4] ;
 wire \mixed_output[5] ;
 wire \mixed_output[6] ;
 wire \mixed_output[7] ;
 wire \mixed_output[8] ;
 wire \mixed_output[9] ;
 wire \state[0] ;
 wire \state[1] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sky130_fd_sc_hd__nor2b_2 _0576_ (.A(\state[0] ),
    .B_N(\state[1] ),
    .Y(_0141_));
 sky130_fd_sc_hd__clkbuf_2 _0577_ (.A(_0141_),
    .X(_0142_));
 sky130_fd_sc_hd__and2_0 _0578_ (.A(\mixed_output[1] ),
    .B(_0142_),
    .X(net15));
 sky130_fd_sc_hd__and2_0 _0579_ (.A(\mixed_output[0] ),
    .B(_0142_),
    .X(net4));
 sky130_fd_sc_hd__and2_0 _0580_ (.A(\mixed_output[3] ),
    .B(_0142_),
    .X(net29));
 sky130_fd_sc_hd__and2_0 _0581_ (.A(\mixed_output[2] ),
    .B(_0141_),
    .X(net26));
 sky130_fd_sc_hd__and2_0 _0582_ (.A(\mixed_output[5] ),
    .B(_0142_),
    .X(net31));
 sky130_fd_sc_hd__and2_0 _0583_ (.A(\mixed_output[4] ),
    .B(_0142_),
    .X(net30));
 sky130_fd_sc_hd__and2_0 _0584_ (.A(\mixed_output[7] ),
    .B(_0142_),
    .X(net33));
 sky130_fd_sc_hd__and2_0 _0585_ (.A(\mixed_output[6] ),
    .B(_0142_),
    .X(net32));
 sky130_fd_sc_hd__and2_0 _0586_ (.A(\mixed_output[9] ),
    .B(_0142_),
    .X(net35));
 sky130_fd_sc_hd__and2_0 _0587_ (.A(\mixed_output[8] ),
    .B(_0142_),
    .X(net34));
 sky130_fd_sc_hd__and2_0 _0588_ (.A(\mixed_output[11] ),
    .B(_0142_),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 _0589_ (.A(_0141_),
    .X(_0143_));
 sky130_fd_sc_hd__and2_0 _0590_ (.A(\mixed_output[10] ),
    .B(_0143_),
    .X(net5));
 sky130_fd_sc_hd__and2_0 _0591_ (.A(\mixed_output[13] ),
    .B(_0143_),
    .X(net8));
 sky130_fd_sc_hd__and2_0 _0592_ (.A(\mixed_output[12] ),
    .B(_0143_),
    .X(net7));
 sky130_fd_sc_hd__and2_0 _0593_ (.A(\mixed_output[15] ),
    .B(_0143_),
    .X(net10));
 sky130_fd_sc_hd__and2_0 _0594_ (.A(\mixed_output[14] ),
    .B(_0143_),
    .X(net9));
 sky130_fd_sc_hd__and2_0 _0595_ (.A(\mixed_output[17] ),
    .B(_0143_),
    .X(net12));
 sky130_fd_sc_hd__and2_0 _0596_ (.A(\mixed_output[16] ),
    .B(_0143_),
    .X(net11));
 sky130_fd_sc_hd__and2_0 _0597_ (.A(\mixed_output[19] ),
    .B(_0143_),
    .X(net14));
 sky130_fd_sc_hd__and2_0 _0598_ (.A(\mixed_output[18] ),
    .B(_0143_),
    .X(net13));
 sky130_fd_sc_hd__and2_0 _0599_ (.A(\mixed_output[21] ),
    .B(_0143_),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 _0600_ (.A(_0141_),
    .X(_0144_));
 sky130_fd_sc_hd__and2_0 _0601_ (.A(\mixed_output[20] ),
    .B(_0144_),
    .X(net16));
 sky130_fd_sc_hd__and2_0 _0602_ (.A(\mixed_output[23] ),
    .B(_0144_),
    .X(net19));
 sky130_fd_sc_hd__and2_0 _0603_ (.A(\mixed_output[22] ),
    .B(_0144_),
    .X(net18));
 sky130_fd_sc_hd__and2_0 _0604_ (.A(\mixed_output[25] ),
    .B(_0144_),
    .X(net21));
 sky130_fd_sc_hd__and2_0 _0605_ (.A(\mixed_output[24] ),
    .B(_0144_),
    .X(net20));
 sky130_fd_sc_hd__and2_0 _0606_ (.A(\mixed_output[27] ),
    .B(_0144_),
    .X(net23));
 sky130_fd_sc_hd__and2_0 _0607_ (.A(\mixed_output[26] ),
    .B(_0144_),
    .X(net22));
 sky130_fd_sc_hd__and2_0 _0608_ (.A(\mixed_output[29] ),
    .B(_0144_),
    .X(net25));
 sky130_fd_sc_hd__and2_0 _0609_ (.A(\mixed_output[28] ),
    .B(_0144_),
    .X(net24));
 sky130_fd_sc_hd__and2_0 _0610_ (.A(\mixed_output[31] ),
    .B(_0144_),
    .X(net28));
 sky130_fd_sc_hd__and2_0 _0611_ (.A(\mixed_output[30] ),
    .B(_0141_),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 _0612_ (.A(rst_n),
    .X(_0145_));
 sky130_fd_sc_hd__inv_1 _0613_ (.A(_0145_),
    .Y(_0146_));
 sky130_fd_sc_hd__clkbuf_4 _0614_ (.A(_0146_),
    .X(_0147_));
 sky130_fd_sc_hd__clkbuf_4 _0615_ (.A(_0147_),
    .X(_0000_));
 sky130_fd_sc_hd__inv_1 _0616_ (.A(\health_counter[0] ),
    .Y(_0570_));
 sky130_fd_sc_hd__inv_1 _0617_ (.A(\health_counter[1] ),
    .Y(_0571_));
 sky130_fd_sc_hd__or2_0 _0618_ (.A(\gen_ring_osc.init_osc ),
    .B(\gen_ring_osc.inv_chain[1] ),
    .X(\gen_ring_osc.inv_chain[1] ));
 sky130_fd_sc_hd__nand3b_4 _0619_ (.A_N(\state[0] ),
    .B(\state[1] ),
    .C(_0145_),
    .Y(_0148_));
 sky130_fd_sc_hd__inv_1 _0620_ (.A(_0148_),
    .Y(_0149_));
 sky130_fd_sc_hd__buf_2 _0621_ (.A(_0149_),
    .X(_0001_));
 sky130_fd_sc_hd__clkbuf_4 _0622_ (.A(_0145_),
    .X(_0150_));
 sky130_fd_sc_hd__clkbuf_4 _0623_ (.A(_0150_),
    .X(_0151_));
 sky130_fd_sc_hd__clkbuf_2 _0624_ (.A(enable),
    .X(_0152_));
 sky130_fd_sc_hd__nor2b_2 _0625_ (.A(\state[1] ),
    .B_N(\state[0] ),
    .Y(_0153_));
 sky130_fd_sc_hd__nand2_1 _0626_ (.A(_0152_),
    .B(_0153_),
    .Y(_0154_));
 sky130_fd_sc_hd__buf_2 _0627_ (.A(_0154_),
    .X(_0155_));
 sky130_fd_sc_hd__buf_2 _0628_ (.A(_0155_),
    .X(_0156_));
 sky130_fd_sc_hd__nand2_1 _0629_ (.A(\entropy_pool2[0] ),
    .B(_0156_),
    .Y(_0157_));
 sky130_fd_sc_hd__and2_0 _0630_ (.A(_0152_),
    .B(_0153_),
    .X(_0158_));
 sky130_fd_sc_hd__buf_2 _0631_ (.A(_0158_),
    .X(_0159_));
 sky130_fd_sc_hd__buf_2 _0632_ (.A(_0159_),
    .X(_0160_));
 sky130_fd_sc_hd__nand2_1 _0633_ (.A(\entropy_pool2[1] ),
    .B(_0160_),
    .Y(_0161_));
 sky130_fd_sc_hd__nand3_1 _0634_ (.A(_0151_),
    .B(_0157_),
    .C(_0161_),
    .Y(_0002_));
 sky130_fd_sc_hd__nand2_1 _0635_ (.A(\entropy_pool2[10] ),
    .B(_0156_),
    .Y(_0162_));
 sky130_fd_sc_hd__nand2_1 _0636_ (.A(\entropy_pool2[11] ),
    .B(_0160_),
    .Y(_0163_));
 sky130_fd_sc_hd__nand3_1 _0637_ (.A(_0151_),
    .B(_0162_),
    .C(_0163_),
    .Y(_0003_));
 sky130_fd_sc_hd__nand2_1 _0638_ (.A(\entropy_pool2[11] ),
    .B(_0156_),
    .Y(_0164_));
 sky130_fd_sc_hd__nand2_1 _0639_ (.A(\entropy_pool2[12] ),
    .B(_0160_),
    .Y(_0165_));
 sky130_fd_sc_hd__nand3_1 _0640_ (.A(_0151_),
    .B(_0164_),
    .C(_0165_),
    .Y(_0004_));
 sky130_fd_sc_hd__buf_2 _0641_ (.A(_0150_),
    .X(_0166_));
 sky130_fd_sc_hd__nand2_1 _0642_ (.A(\entropy_pool2[12] ),
    .B(_0156_),
    .Y(_0167_));
 sky130_fd_sc_hd__nand2_1 _0643_ (.A(\entropy_pool2[13] ),
    .B(_0160_),
    .Y(_0168_));
 sky130_fd_sc_hd__nand3_1 _0644_ (.A(_0166_),
    .B(_0167_),
    .C(_0168_),
    .Y(_0005_));
 sky130_fd_sc_hd__nand2_1 _0645_ (.A(\entropy_pool2[13] ),
    .B(_0156_),
    .Y(_0169_));
 sky130_fd_sc_hd__nand2_1 _0646_ (.A(\entropy_pool2[14] ),
    .B(_0160_),
    .Y(_0170_));
 sky130_fd_sc_hd__nand3_1 _0647_ (.A(_0166_),
    .B(_0169_),
    .C(_0170_),
    .Y(_0006_));
 sky130_fd_sc_hd__nand2_1 _0648_ (.A(\entropy_pool2[14] ),
    .B(_0156_),
    .Y(_0171_));
 sky130_fd_sc_hd__nand2_1 _0649_ (.A(\entropy_pool2[15] ),
    .B(_0160_),
    .Y(_0172_));
 sky130_fd_sc_hd__nand3_1 _0650_ (.A(_0166_),
    .B(_0171_),
    .C(_0172_),
    .Y(_0007_));
 sky130_fd_sc_hd__nand2_1 _0651_ (.A(\entropy_pool2[15] ),
    .B(_0156_),
    .Y(_0173_));
 sky130_fd_sc_hd__nand2_1 _0652_ (.A(\entropy_pool2[16] ),
    .B(_0160_),
    .Y(_0174_));
 sky130_fd_sc_hd__nand3_1 _0653_ (.A(_0166_),
    .B(_0173_),
    .C(_0174_),
    .Y(_0008_));
 sky130_fd_sc_hd__nand2_1 _0654_ (.A(\entropy_pool2[16] ),
    .B(_0156_),
    .Y(_0175_));
 sky130_fd_sc_hd__nand2_1 _0655_ (.A(\entropy_pool2[17] ),
    .B(_0160_),
    .Y(_0176_));
 sky130_fd_sc_hd__nand3_1 _0656_ (.A(_0166_),
    .B(_0175_),
    .C(_0176_),
    .Y(_0009_));
 sky130_fd_sc_hd__nand2_1 _0657_ (.A(\entropy_pool2[17] ),
    .B(_0156_),
    .Y(_0177_));
 sky130_fd_sc_hd__nand2_1 _0658_ (.A(\entropy_pool2[18] ),
    .B(_0160_),
    .Y(_0178_));
 sky130_fd_sc_hd__nand3_1 _0659_ (.A(_0166_),
    .B(_0177_),
    .C(_0178_),
    .Y(_0010_));
 sky130_fd_sc_hd__nand2_1 _0660_ (.A(\entropy_pool2[18] ),
    .B(_0156_),
    .Y(_0179_));
 sky130_fd_sc_hd__nand2_1 _0661_ (.A(\entropy_pool2[19] ),
    .B(_0160_),
    .Y(_0180_));
 sky130_fd_sc_hd__nand3_1 _0662_ (.A(_0166_),
    .B(_0179_),
    .C(_0180_),
    .Y(_0011_));
 sky130_fd_sc_hd__buf_2 _0663_ (.A(_0155_),
    .X(_0181_));
 sky130_fd_sc_hd__nand2_1 _0664_ (.A(\entropy_pool2[19] ),
    .B(_0181_),
    .Y(_0182_));
 sky130_fd_sc_hd__buf_2 _0665_ (.A(_0159_),
    .X(_0183_));
 sky130_fd_sc_hd__nand2_1 _0666_ (.A(\entropy_pool2[20] ),
    .B(_0183_),
    .Y(_0184_));
 sky130_fd_sc_hd__nand3_1 _0667_ (.A(_0166_),
    .B(_0182_),
    .C(_0184_),
    .Y(_0012_));
 sky130_fd_sc_hd__nand2_1 _0668_ (.A(\entropy_pool2[1] ),
    .B(_0181_),
    .Y(_0185_));
 sky130_fd_sc_hd__nand2_1 _0669_ (.A(\entropy_pool2[2] ),
    .B(_0183_),
    .Y(_0186_));
 sky130_fd_sc_hd__nand3_1 _0670_ (.A(_0166_),
    .B(_0185_),
    .C(_0186_),
    .Y(_0013_));
 sky130_fd_sc_hd__nand2_1 _0671_ (.A(\entropy_pool2[20] ),
    .B(_0181_),
    .Y(_0187_));
 sky130_fd_sc_hd__nand2_1 _0672_ (.A(\entropy_pool2[21] ),
    .B(_0183_),
    .Y(_0188_));
 sky130_fd_sc_hd__nand3_1 _0673_ (.A(_0166_),
    .B(_0187_),
    .C(_0188_),
    .Y(_0014_));
 sky130_fd_sc_hd__buf_2 _0674_ (.A(_0150_),
    .X(_0189_));
 sky130_fd_sc_hd__nand2_1 _0675_ (.A(\entropy_pool2[21] ),
    .B(_0181_),
    .Y(_0190_));
 sky130_fd_sc_hd__nand2_1 _0676_ (.A(\entropy_pool2[22] ),
    .B(_0183_),
    .Y(_0191_));
 sky130_fd_sc_hd__nand3_1 _0677_ (.A(_0189_),
    .B(_0190_),
    .C(_0191_),
    .Y(_0015_));
 sky130_fd_sc_hd__nand2_1 _0678_ (.A(\entropy_pool2[22] ),
    .B(_0181_),
    .Y(_0192_));
 sky130_fd_sc_hd__nand2_1 _0679_ (.A(\entropy_pool2[23] ),
    .B(_0183_),
    .Y(_0193_));
 sky130_fd_sc_hd__nand3_1 _0680_ (.A(_0189_),
    .B(_0192_),
    .C(_0193_),
    .Y(_0016_));
 sky130_fd_sc_hd__nand2_1 _0681_ (.A(\entropy_pool2[23] ),
    .B(_0181_),
    .Y(_0194_));
 sky130_fd_sc_hd__nand2_1 _0682_ (.A(\entropy_pool2[24] ),
    .B(_0183_),
    .Y(_0195_));
 sky130_fd_sc_hd__nand3_1 _0683_ (.A(_0189_),
    .B(_0194_),
    .C(_0195_),
    .Y(_0017_));
 sky130_fd_sc_hd__nand2_1 _0684_ (.A(\entropy_pool2[24] ),
    .B(_0181_),
    .Y(_0196_));
 sky130_fd_sc_hd__nand2_1 _0685_ (.A(\entropy_pool2[25] ),
    .B(_0183_),
    .Y(_0197_));
 sky130_fd_sc_hd__nand3_1 _0686_ (.A(_0189_),
    .B(_0196_),
    .C(_0197_),
    .Y(_0018_));
 sky130_fd_sc_hd__nand2_1 _0687_ (.A(\entropy_pool2[25] ),
    .B(_0181_),
    .Y(_0198_));
 sky130_fd_sc_hd__nand2_1 _0688_ (.A(\entropy_pool2[26] ),
    .B(_0183_),
    .Y(_0199_));
 sky130_fd_sc_hd__nand3_1 _0689_ (.A(_0189_),
    .B(_0198_),
    .C(_0199_),
    .Y(_0019_));
 sky130_fd_sc_hd__nand2_1 _0690_ (.A(\entropy_pool2[26] ),
    .B(_0181_),
    .Y(_0200_));
 sky130_fd_sc_hd__nand2_1 _0691_ (.A(\entropy_pool2[27] ),
    .B(_0183_),
    .Y(_0201_));
 sky130_fd_sc_hd__nand3_1 _0692_ (.A(_0189_),
    .B(_0200_),
    .C(_0201_),
    .Y(_0020_));
 sky130_fd_sc_hd__nand2_1 _0693_ (.A(\entropy_pool2[27] ),
    .B(_0181_),
    .Y(_0202_));
 sky130_fd_sc_hd__nand2_1 _0694_ (.A(\entropy_pool2[28] ),
    .B(_0183_),
    .Y(_0203_));
 sky130_fd_sc_hd__nand3_1 _0695_ (.A(_0189_),
    .B(_0202_),
    .C(_0203_),
    .Y(_0021_));
 sky130_fd_sc_hd__buf_2 _0696_ (.A(_0155_),
    .X(_0204_));
 sky130_fd_sc_hd__nand2_1 _0697_ (.A(\entropy_pool2[28] ),
    .B(_0204_),
    .Y(_0205_));
 sky130_fd_sc_hd__buf_2 _0698_ (.A(_0159_),
    .X(_0206_));
 sky130_fd_sc_hd__nand2_1 _0699_ (.A(\entropy_pool2[29] ),
    .B(_0206_),
    .Y(_0207_));
 sky130_fd_sc_hd__nand3_1 _0700_ (.A(_0189_),
    .B(_0205_),
    .C(_0207_),
    .Y(_0022_));
 sky130_fd_sc_hd__nand2_1 _0701_ (.A(\entropy_pool2[29] ),
    .B(_0204_),
    .Y(_0208_));
 sky130_fd_sc_hd__nand2_1 _0702_ (.A(\entropy_pool2[30] ),
    .B(_0206_),
    .Y(_0209_));
 sky130_fd_sc_hd__nand3_1 _0703_ (.A(_0189_),
    .B(_0208_),
    .C(_0209_),
    .Y(_0023_));
 sky130_fd_sc_hd__nand2_1 _0704_ (.A(\entropy_pool2[2] ),
    .B(_0204_),
    .Y(_0210_));
 sky130_fd_sc_hd__nand2_1 _0705_ (.A(\entropy_pool2[3] ),
    .B(_0206_),
    .Y(_0211_));
 sky130_fd_sc_hd__nand3_1 _0706_ (.A(_0189_),
    .B(_0210_),
    .C(_0211_),
    .Y(_0024_));
 sky130_fd_sc_hd__buf_2 _0707_ (.A(_0150_),
    .X(_0212_));
 sky130_fd_sc_hd__nand2_1 _0708_ (.A(\entropy_pool2[30] ),
    .B(_0204_),
    .Y(_0213_));
 sky130_fd_sc_hd__nand2_1 _0709_ (.A(\entropy_pool2[31] ),
    .B(_0206_),
    .Y(_0214_));
 sky130_fd_sc_hd__nand3_1 _0710_ (.A(_0212_),
    .B(_0213_),
    .C(_0214_),
    .Y(_0025_));
 sky130_fd_sc_hd__buf_2 _0711_ (.A(_0154_),
    .X(_0215_));
 sky130_fd_sc_hd__xnor2_1 _0712_ (.A(\entropy_pool2[0] ),
    .B(\gen_ring_osc.toggle_sampling ),
    .Y(_0216_));
 sky130_fd_sc_hd__nand2_1 _0713_ (.A(\entropy_pool2[31] ),
    .B(_0215_),
    .Y(_0217_));
 sky130_fd_sc_hd__o211ai_1 _0714_ (.A1(_0215_),
    .A2(_0216_),
    .B1(_0217_),
    .C1(_0212_),
    .Y(_0026_));
 sky130_fd_sc_hd__nand2_1 _0715_ (.A(\entropy_pool2[3] ),
    .B(_0204_),
    .Y(_0218_));
 sky130_fd_sc_hd__nand2_1 _0716_ (.A(\entropy_pool2[4] ),
    .B(_0206_),
    .Y(_0219_));
 sky130_fd_sc_hd__nand3_1 _0717_ (.A(_0212_),
    .B(_0218_),
    .C(_0219_),
    .Y(_0027_));
 sky130_fd_sc_hd__nand2_1 _0718_ (.A(\entropy_pool2[4] ),
    .B(_0204_),
    .Y(_0220_));
 sky130_fd_sc_hd__nand2_1 _0719_ (.A(\entropy_pool2[5] ),
    .B(_0206_),
    .Y(_0221_));
 sky130_fd_sc_hd__nand3_1 _0720_ (.A(_0212_),
    .B(_0220_),
    .C(_0221_),
    .Y(_0028_));
 sky130_fd_sc_hd__nand2_1 _0721_ (.A(\entropy_pool2[5] ),
    .B(_0204_),
    .Y(_0222_));
 sky130_fd_sc_hd__nand2_1 _0722_ (.A(\entropy_pool2[6] ),
    .B(_0206_),
    .Y(_0223_));
 sky130_fd_sc_hd__nand3_1 _0723_ (.A(_0212_),
    .B(_0222_),
    .C(_0223_),
    .Y(_0029_));
 sky130_fd_sc_hd__nand2_1 _0724_ (.A(\entropy_pool2[6] ),
    .B(_0204_),
    .Y(_0224_));
 sky130_fd_sc_hd__nand2_1 _0725_ (.A(\entropy_pool2[7] ),
    .B(_0206_),
    .Y(_0225_));
 sky130_fd_sc_hd__nand3_1 _0726_ (.A(_0212_),
    .B(_0224_),
    .C(_0225_),
    .Y(_0030_));
 sky130_fd_sc_hd__nand2_1 _0727_ (.A(\entropy_pool2[7] ),
    .B(_0204_),
    .Y(_0226_));
 sky130_fd_sc_hd__nand2_1 _0728_ (.A(\entropy_pool2[8] ),
    .B(_0206_),
    .Y(_0227_));
 sky130_fd_sc_hd__nand3_1 _0729_ (.A(_0212_),
    .B(_0226_),
    .C(_0227_),
    .Y(_0031_));
 sky130_fd_sc_hd__nand2_1 _0730_ (.A(\entropy_pool2[8] ),
    .B(_0204_),
    .Y(_0228_));
 sky130_fd_sc_hd__nand2_1 _0731_ (.A(\entropy_pool2[9] ),
    .B(_0206_),
    .Y(_0229_));
 sky130_fd_sc_hd__nand3_1 _0732_ (.A(_0212_),
    .B(_0228_),
    .C(_0229_),
    .Y(_0032_));
 sky130_fd_sc_hd__nand2_1 _0733_ (.A(\entropy_pool2[9] ),
    .B(_0215_),
    .Y(_0230_));
 sky130_fd_sc_hd__buf_4 _0734_ (.A(_0159_),
    .X(_0231_));
 sky130_fd_sc_hd__nand2_1 _0735_ (.A(\entropy_pool2[10] ),
    .B(_0231_),
    .Y(_0232_));
 sky130_fd_sc_hd__nand3_1 _0736_ (.A(_0212_),
    .B(_0230_),
    .C(_0232_),
    .Y(_0033_));
 sky130_fd_sc_hd__xnor2_1 _0737_ (.A(\entropy_pool[31] ),
    .B(\gen_ring_osc.toggle_sampling ),
    .Y(_0233_));
 sky130_fd_sc_hd__nand2_1 _0738_ (.A(\entropy_pool[0] ),
    .B(_0215_),
    .Y(_0234_));
 sky130_fd_sc_hd__o211ai_1 _0739_ (.A1(_0215_),
    .A2(_0233_),
    .B1(_0234_),
    .C1(_0212_),
    .Y(_0034_));
 sky130_fd_sc_hd__nand2_1 _0740_ (.A(\entropy_pool[9] ),
    .B(_0231_),
    .Y(_0235_));
 sky130_fd_sc_hd__nand2_1 _0741_ (.A(\entropy_pool[10] ),
    .B(_0215_),
    .Y(_0236_));
 sky130_fd_sc_hd__clkbuf_4 _0742_ (.A(_0146_),
    .X(_0237_));
 sky130_fd_sc_hd__a21oi_1 _0743_ (.A1(_0235_),
    .A2(_0236_),
    .B1(_0237_),
    .Y(_0035_));
 sky130_fd_sc_hd__nand2_1 _0744_ (.A(\entropy_pool[10] ),
    .B(_0231_),
    .Y(_0238_));
 sky130_fd_sc_hd__nand2_1 _0745_ (.A(\entropy_pool[11] ),
    .B(_0215_),
    .Y(_0239_));
 sky130_fd_sc_hd__a21oi_1 _0746_ (.A1(_0238_),
    .A2(_0239_),
    .B1(_0237_),
    .Y(_0036_));
 sky130_fd_sc_hd__nand2_1 _0747_ (.A(\entropy_pool[11] ),
    .B(_0231_),
    .Y(_0240_));
 sky130_fd_sc_hd__nand2_1 _0748_ (.A(\entropy_pool[12] ),
    .B(_0215_),
    .Y(_0241_));
 sky130_fd_sc_hd__a21oi_1 _0749_ (.A1(_0240_),
    .A2(_0241_),
    .B1(_0237_),
    .Y(_0037_));
 sky130_fd_sc_hd__nand2_1 _0750_ (.A(\entropy_pool[12] ),
    .B(_0231_),
    .Y(_0242_));
 sky130_fd_sc_hd__nand2_1 _0751_ (.A(\entropy_pool[13] ),
    .B(_0215_),
    .Y(_0243_));
 sky130_fd_sc_hd__buf_2 _0752_ (.A(_0147_),
    .X(_0244_));
 sky130_fd_sc_hd__a21oi_1 _0753_ (.A1(_0242_),
    .A2(_0243_),
    .B1(_0244_),
    .Y(_0038_));
 sky130_fd_sc_hd__nand2_1 _0754_ (.A(\entropy_pool[13] ),
    .B(_0231_),
    .Y(_0245_));
 sky130_fd_sc_hd__nand2_1 _0755_ (.A(\entropy_pool[14] ),
    .B(_0215_),
    .Y(_0246_));
 sky130_fd_sc_hd__a21oi_1 _0756_ (.A1(_0245_),
    .A2(_0246_),
    .B1(_0244_),
    .Y(_0039_));
 sky130_fd_sc_hd__nand2_1 _0757_ (.A(\entropy_pool[14] ),
    .B(_0231_),
    .Y(_0247_));
 sky130_fd_sc_hd__buf_2 _0758_ (.A(_0155_),
    .X(_0248_));
 sky130_fd_sc_hd__nand2_1 _0759_ (.A(\entropy_pool[15] ),
    .B(_0248_),
    .Y(_0249_));
 sky130_fd_sc_hd__a21oi_1 _0760_ (.A1(_0247_),
    .A2(_0249_),
    .B1(_0244_),
    .Y(_0040_));
 sky130_fd_sc_hd__nand2_1 _0761_ (.A(\entropy_pool[15] ),
    .B(_0231_),
    .Y(_0250_));
 sky130_fd_sc_hd__nand2_1 _0762_ (.A(\entropy_pool[16] ),
    .B(_0248_),
    .Y(_0251_));
 sky130_fd_sc_hd__a21oi_1 _0763_ (.A1(_0250_),
    .A2(_0251_),
    .B1(_0244_),
    .Y(_0041_));
 sky130_fd_sc_hd__nand2_1 _0764_ (.A(\entropy_pool[16] ),
    .B(_0231_),
    .Y(_0252_));
 sky130_fd_sc_hd__nand2_1 _0765_ (.A(\entropy_pool[17] ),
    .B(_0248_),
    .Y(_0253_));
 sky130_fd_sc_hd__a21oi_1 _0766_ (.A1(_0252_),
    .A2(_0253_),
    .B1(_0244_),
    .Y(_0042_));
 sky130_fd_sc_hd__nand2_1 _0767_ (.A(\entropy_pool[17] ),
    .B(_0231_),
    .Y(_0254_));
 sky130_fd_sc_hd__nand2_1 _0768_ (.A(\entropy_pool[18] ),
    .B(_0248_),
    .Y(_0255_));
 sky130_fd_sc_hd__a21oi_1 _0769_ (.A1(_0254_),
    .A2(_0255_),
    .B1(_0244_),
    .Y(_0043_));
 sky130_fd_sc_hd__buf_4 _0770_ (.A(_0159_),
    .X(_0256_));
 sky130_fd_sc_hd__nand2_1 _0771_ (.A(\entropy_pool[18] ),
    .B(_0256_),
    .Y(_0257_));
 sky130_fd_sc_hd__nand2_1 _0772_ (.A(\entropy_pool[19] ),
    .B(_0248_),
    .Y(_0258_));
 sky130_fd_sc_hd__a21oi_1 _0773_ (.A1(_0257_),
    .A2(_0258_),
    .B1(_0244_),
    .Y(_0044_));
 sky130_fd_sc_hd__nand2_1 _0774_ (.A(\entropy_pool[0] ),
    .B(_0256_),
    .Y(_0259_));
 sky130_fd_sc_hd__nand2_1 _0775_ (.A(\entropy_pool[1] ),
    .B(_0248_),
    .Y(_0260_));
 sky130_fd_sc_hd__a21oi_1 _0776_ (.A1(_0259_),
    .A2(_0260_),
    .B1(_0244_),
    .Y(_0045_));
 sky130_fd_sc_hd__nand2_1 _0777_ (.A(\entropy_pool[19] ),
    .B(_0256_),
    .Y(_0261_));
 sky130_fd_sc_hd__nand2_1 _0778_ (.A(\entropy_pool[20] ),
    .B(_0248_),
    .Y(_0262_));
 sky130_fd_sc_hd__a21oi_1 _0779_ (.A1(_0261_),
    .A2(_0262_),
    .B1(_0244_),
    .Y(_0046_));
 sky130_fd_sc_hd__nand2_1 _0780_ (.A(\entropy_pool[20] ),
    .B(_0256_),
    .Y(_0263_));
 sky130_fd_sc_hd__nand2_1 _0781_ (.A(\entropy_pool[21] ),
    .B(_0248_),
    .Y(_0264_));
 sky130_fd_sc_hd__a21oi_1 _0782_ (.A1(_0263_),
    .A2(_0264_),
    .B1(_0244_),
    .Y(_0047_));
 sky130_fd_sc_hd__nand2_1 _0783_ (.A(\entropy_pool[21] ),
    .B(_0256_),
    .Y(_0265_));
 sky130_fd_sc_hd__nand2_1 _0784_ (.A(\entropy_pool[22] ),
    .B(_0248_),
    .Y(_0266_));
 sky130_fd_sc_hd__clkbuf_4 _0785_ (.A(_0146_),
    .X(_0267_));
 sky130_fd_sc_hd__a21oi_1 _0786_ (.A1(_0265_),
    .A2(_0266_),
    .B1(_0267_),
    .Y(_0048_));
 sky130_fd_sc_hd__nand2_1 _0787_ (.A(\entropy_pool[22] ),
    .B(_0256_),
    .Y(_0268_));
 sky130_fd_sc_hd__nand2_1 _0788_ (.A(\entropy_pool[23] ),
    .B(_0248_),
    .Y(_0269_));
 sky130_fd_sc_hd__a21oi_1 _0789_ (.A1(_0268_),
    .A2(_0269_),
    .B1(_0267_),
    .Y(_0049_));
 sky130_fd_sc_hd__nand2_1 _0790_ (.A(\entropy_pool[23] ),
    .B(_0256_),
    .Y(_0270_));
 sky130_fd_sc_hd__clkbuf_4 _0791_ (.A(_0154_),
    .X(_0271_));
 sky130_fd_sc_hd__nand2_1 _0792_ (.A(\entropy_pool[24] ),
    .B(_0271_),
    .Y(_0272_));
 sky130_fd_sc_hd__a21oi_1 _0793_ (.A1(_0270_),
    .A2(_0272_),
    .B1(_0267_),
    .Y(_0050_));
 sky130_fd_sc_hd__nand2_1 _0794_ (.A(\entropy_pool[24] ),
    .B(_0256_),
    .Y(_0273_));
 sky130_fd_sc_hd__nand2_1 _0795_ (.A(\entropy_pool[25] ),
    .B(_0271_),
    .Y(_0274_));
 sky130_fd_sc_hd__a21oi_1 _0796_ (.A1(_0273_),
    .A2(_0274_),
    .B1(_0267_),
    .Y(_0051_));
 sky130_fd_sc_hd__nand2_1 _0797_ (.A(\entropy_pool[25] ),
    .B(_0256_),
    .Y(_0275_));
 sky130_fd_sc_hd__nand2_1 _0798_ (.A(\entropy_pool[26] ),
    .B(_0271_),
    .Y(_0276_));
 sky130_fd_sc_hd__a21oi_1 _0799_ (.A1(_0275_),
    .A2(_0276_),
    .B1(_0267_),
    .Y(_0052_));
 sky130_fd_sc_hd__nand2_1 _0800_ (.A(\entropy_pool[26] ),
    .B(_0256_),
    .Y(_0277_));
 sky130_fd_sc_hd__nand2_1 _0801_ (.A(\entropy_pool[27] ),
    .B(_0271_),
    .Y(_0278_));
 sky130_fd_sc_hd__a21oi_1 _0802_ (.A1(_0277_),
    .A2(_0278_),
    .B1(_0267_),
    .Y(_0053_));
 sky130_fd_sc_hd__buf_4 _0803_ (.A(_0159_),
    .X(_0279_));
 sky130_fd_sc_hd__nand2_1 _0804_ (.A(\entropy_pool[27] ),
    .B(_0279_),
    .Y(_0280_));
 sky130_fd_sc_hd__nand2_1 _0805_ (.A(\entropy_pool[28] ),
    .B(_0271_),
    .Y(_0281_));
 sky130_fd_sc_hd__a21oi_1 _0806_ (.A1(_0280_),
    .A2(_0281_),
    .B1(_0267_),
    .Y(_0054_));
 sky130_fd_sc_hd__nand2_1 _0807_ (.A(\entropy_pool[28] ),
    .B(_0279_),
    .Y(_0282_));
 sky130_fd_sc_hd__nand2_1 _0808_ (.A(\entropy_pool[29] ),
    .B(_0271_),
    .Y(_0283_));
 sky130_fd_sc_hd__a21oi_1 _0809_ (.A1(_0282_),
    .A2(_0283_),
    .B1(_0267_),
    .Y(_0055_));
 sky130_fd_sc_hd__nand2_1 _0810_ (.A(\entropy_pool[1] ),
    .B(_0279_),
    .Y(_0284_));
 sky130_fd_sc_hd__nand2_1 _0811_ (.A(\entropy_pool[2] ),
    .B(_0271_),
    .Y(_0285_));
 sky130_fd_sc_hd__a21oi_1 _0812_ (.A1(_0284_),
    .A2(_0285_),
    .B1(_0267_),
    .Y(_0056_));
 sky130_fd_sc_hd__nand2_1 _0813_ (.A(\entropy_pool[29] ),
    .B(_0279_),
    .Y(_0286_));
 sky130_fd_sc_hd__nand2_1 _0814_ (.A(\entropy_pool[30] ),
    .B(_0271_),
    .Y(_0287_));
 sky130_fd_sc_hd__a21oi_1 _0815_ (.A1(_0286_),
    .A2(_0287_),
    .B1(_0267_),
    .Y(_0057_));
 sky130_fd_sc_hd__nand2_1 _0816_ (.A(\entropy_pool[30] ),
    .B(_0279_),
    .Y(_0288_));
 sky130_fd_sc_hd__nand2_1 _0817_ (.A(\entropy_pool[31] ),
    .B(_0271_),
    .Y(_0289_));
 sky130_fd_sc_hd__a21oi_1 _0818_ (.A1(_0288_),
    .A2(_0289_),
    .B1(_0147_),
    .Y(_0058_));
 sky130_fd_sc_hd__nand2_1 _0819_ (.A(\entropy_pool[2] ),
    .B(_0279_),
    .Y(_0290_));
 sky130_fd_sc_hd__nand2_1 _0820_ (.A(\entropy_pool[3] ),
    .B(_0271_),
    .Y(_0291_));
 sky130_fd_sc_hd__a21oi_1 _0821_ (.A1(_0290_),
    .A2(_0291_),
    .B1(_0147_),
    .Y(_0059_));
 sky130_fd_sc_hd__nand2_1 _0822_ (.A(\entropy_pool[3] ),
    .B(_0279_),
    .Y(_0292_));
 sky130_fd_sc_hd__nand2_1 _0823_ (.A(\entropy_pool[4] ),
    .B(_0155_),
    .Y(_0293_));
 sky130_fd_sc_hd__a21oi_1 _0824_ (.A1(_0292_),
    .A2(_0293_),
    .B1(_0147_),
    .Y(_0060_));
 sky130_fd_sc_hd__nand2_1 _0825_ (.A(\entropy_pool[4] ),
    .B(_0279_),
    .Y(_0294_));
 sky130_fd_sc_hd__nand2_1 _0826_ (.A(\entropy_pool[5] ),
    .B(_0155_),
    .Y(_0295_));
 sky130_fd_sc_hd__a21oi_1 _0827_ (.A1(_0294_),
    .A2(_0295_),
    .B1(_0147_),
    .Y(_0061_));
 sky130_fd_sc_hd__nand2_1 _0828_ (.A(\entropy_pool[5] ),
    .B(_0279_),
    .Y(_0296_));
 sky130_fd_sc_hd__nand2_1 _0829_ (.A(\entropy_pool[6] ),
    .B(_0155_),
    .Y(_0297_));
 sky130_fd_sc_hd__a21oi_1 _0830_ (.A1(_0296_),
    .A2(_0297_),
    .B1(_0147_),
    .Y(_0062_));
 sky130_fd_sc_hd__nand2_1 _0831_ (.A(\entropy_pool[6] ),
    .B(_0279_),
    .Y(_0298_));
 sky130_fd_sc_hd__nand2_1 _0832_ (.A(\entropy_pool[7] ),
    .B(_0155_),
    .Y(_0299_));
 sky130_fd_sc_hd__a21oi_1 _0833_ (.A1(_0298_),
    .A2(_0299_),
    .B1(_0147_),
    .Y(_0063_));
 sky130_fd_sc_hd__nand2_1 _0834_ (.A(\entropy_pool[7] ),
    .B(_0159_),
    .Y(_0300_));
 sky130_fd_sc_hd__nand2_1 _0835_ (.A(\entropy_pool[8] ),
    .B(_0155_),
    .Y(_0301_));
 sky130_fd_sc_hd__a21oi_1 _0836_ (.A1(_0300_),
    .A2(_0301_),
    .B1(_0147_),
    .Y(_0064_));
 sky130_fd_sc_hd__nand2_1 _0837_ (.A(\entropy_pool[8] ),
    .B(_0159_),
    .Y(_0302_));
 sky130_fd_sc_hd__nand2_1 _0838_ (.A(\entropy_pool[9] ),
    .B(_0155_),
    .Y(_0303_));
 sky130_fd_sc_hd__a21oi_1 _0839_ (.A1(_0302_),
    .A2(_0303_),
    .B1(_0147_),
    .Y(_0065_));
 sky130_fd_sc_hd__buf_4 _0840_ (.A(_0152_),
    .X(_0304_));
 sky130_fd_sc_hd__mux2i_1 _0841_ (.A0(\gen_ring_osc.toggle_sampling ),
    .A1(\gen_ring_osc.inv_chain[1] ),
    .S(_0304_),
    .Y(_0305_));
 sky130_fd_sc_hd__nor2_1 _0842_ (.A(_0000_),
    .B(_0305_),
    .Y(_0066_));
 sky130_fd_sc_hd__buf_2 _0843_ (.A(\state[1] ),
    .X(_0306_));
 sky130_fd_sc_hd__mux2i_1 _0844_ (.A0(_0306_),
    .A1(_0153_),
    .S(_0570_),
    .Y(_0307_));
 sky130_fd_sc_hd__nor2_1 _0845_ (.A(_0000_),
    .B(_0307_),
    .Y(_0067_));
 sky130_fd_sc_hd__a22oi_1 _0846_ (.A1(_0306_),
    .A2(\health_counter[1] ),
    .B1(_0573_),
    .B2(_0153_),
    .Y(_0308_));
 sky130_fd_sc_hd__nor2_1 _0847_ (.A(_0000_),
    .B(_0308_),
    .Y(_0068_));
 sky130_fd_sc_hd__o21ai_2 _0848_ (.A1(\state[0] ),
    .A2(_0306_),
    .B1(_0145_),
    .Y(_0309_));
 sky130_fd_sc_hd__nor2b_1 _0849_ (.A(_0306_),
    .B_N(_0574_),
    .Y(_0310_));
 sky130_fd_sc_hd__xnor2_1 _0850_ (.A(\health_counter[2] ),
    .B(_0310_),
    .Y(_0311_));
 sky130_fd_sc_hd__nor2_1 _0851_ (.A(_0309_),
    .B(_0311_),
    .Y(_0069_));
 sky130_fd_sc_hd__nand4b_1 _0852_ (.A_N(_0306_),
    .B(\health_counter[2] ),
    .C(\health_counter[0] ),
    .D(\health_counter[1] ),
    .Y(_0312_));
 sky130_fd_sc_hd__xor2_1 _0853_ (.A(\health_counter[3] ),
    .B(_0312_),
    .X(_0313_));
 sky130_fd_sc_hd__nor2_1 _0854_ (.A(_0309_),
    .B(_0313_),
    .Y(_0070_));
 sky130_fd_sc_hd__nand4b_1 _0855_ (.A_N(_0306_),
    .B(\health_counter[3] ),
    .C(\health_counter[2] ),
    .D(_0574_),
    .Y(_0314_));
 sky130_fd_sc_hd__xor2_1 _0856_ (.A(\health_counter[4] ),
    .B(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__nor2_1 _0857_ (.A(_0309_),
    .B(_0315_),
    .Y(_0071_));
 sky130_fd_sc_hd__and4b_1 _0858_ (.A_N(\state[1] ),
    .B(\health_counter[4] ),
    .C(\health_counter[3] ),
    .D(\health_counter[2] ),
    .X(_0316_));
 sky130_fd_sc_hd__nand3_1 _0859_ (.A(\health_counter[0] ),
    .B(\health_counter[1] ),
    .C(_0316_),
    .Y(_0317_));
 sky130_fd_sc_hd__xor2_1 _0860_ (.A(\health_counter[5] ),
    .B(_0317_),
    .X(_0318_));
 sky130_fd_sc_hd__nor2_1 _0861_ (.A(_0309_),
    .B(_0318_),
    .Y(_0072_));
 sky130_fd_sc_hd__nand3_1 _0862_ (.A(\health_counter[5] ),
    .B(_0574_),
    .C(_0316_),
    .Y(_0319_));
 sky130_fd_sc_hd__xor2_1 _0863_ (.A(\health_counter[6] ),
    .B(_0319_),
    .X(_0320_));
 sky130_fd_sc_hd__nor2_1 _0864_ (.A(_0309_),
    .B(_0320_),
    .Y(_0073_));
 sky130_fd_sc_hd__and3_1 _0865_ (.A(\health_counter[6] ),
    .B(\health_counter[0] ),
    .C(\health_counter[1] ),
    .X(_0321_));
 sky130_fd_sc_hd__nand3_1 _0866_ (.A(\health_counter[5] ),
    .B(_0316_),
    .C(_0321_),
    .Y(_0322_));
 sky130_fd_sc_hd__xor2_1 _0867_ (.A(\health_counter[7] ),
    .B(_0322_),
    .X(_0323_));
 sky130_fd_sc_hd__nor2_1 _0868_ (.A(_0309_),
    .B(_0323_),
    .Y(_0074_));
 sky130_fd_sc_hd__buf_2 _0869_ (.A(_0150_),
    .X(_0324_));
 sky130_fd_sc_hd__buf_2 _0870_ (.A(\lfsr_reg[31] ),
    .X(_0325_));
 sky130_fd_sc_hd__clkbuf_4 _0871_ (.A(_0152_),
    .X(_0326_));
 sky130_fd_sc_hd__mux2i_1 _0872_ (.A0(\lfsr_reg[0] ),
    .A1(_0325_),
    .S(_0326_),
    .Y(_0327_));
 sky130_fd_sc_hd__nand2_1 _0873_ (.A(_0324_),
    .B(_0327_),
    .Y(_0075_));
 sky130_fd_sc_hd__mux2i_1 _0874_ (.A0(\lfsr_reg[10] ),
    .A1(\lfsr_reg[9] ),
    .S(_0304_),
    .Y(_0328_));
 sky130_fd_sc_hd__nor2_1 _0875_ (.A(_0000_),
    .B(_0328_),
    .Y(_0076_));
 sky130_fd_sc_hd__xnor2_1 _0876_ (.A(\lfsr_reg[30] ),
    .B(\lfsr_reg[10] ),
    .Y(_0329_));
 sky130_fd_sc_hd__nand2_1 _0877_ (.A(_0326_),
    .B(_0329_),
    .Y(_0330_));
 sky130_fd_sc_hd__o21ai_0 _0878_ (.A1(_0326_),
    .A2(\lfsr_reg[11] ),
    .B1(_0330_),
    .Y(_0331_));
 sky130_fd_sc_hd__nand2_1 _0879_ (.A(_0324_),
    .B(_0331_),
    .Y(_0077_));
 sky130_fd_sc_hd__mux2i_1 _0880_ (.A0(\lfsr_reg[12] ),
    .A1(\lfsr_reg[11] ),
    .S(_0304_),
    .Y(_0332_));
 sky130_fd_sc_hd__nor2_1 _0881_ (.A(_0000_),
    .B(_0332_),
    .Y(_0078_));
 sky130_fd_sc_hd__buf_4 _0882_ (.A(_0152_),
    .X(_0333_));
 sky130_fd_sc_hd__mux2i_1 _0883_ (.A0(\lfsr_reg[13] ),
    .A1(\lfsr_reg[12] ),
    .S(_0333_),
    .Y(_0334_));
 sky130_fd_sc_hd__nand2_1 _0884_ (.A(_0324_),
    .B(_0334_),
    .Y(_0079_));
 sky130_fd_sc_hd__mux2i_1 _0885_ (.A0(\lfsr_reg[14] ),
    .A1(\lfsr_reg[13] ),
    .S(_0333_),
    .Y(_0335_));
 sky130_fd_sc_hd__nand2_1 _0886_ (.A(_0324_),
    .B(_0335_),
    .Y(_0080_));
 sky130_fd_sc_hd__mux2i_1 _0887_ (.A0(\lfsr_reg[15] ),
    .A1(\lfsr_reg[14] ),
    .S(_0333_),
    .Y(_0336_));
 sky130_fd_sc_hd__nand2_1 _0888_ (.A(_0324_),
    .B(_0336_),
    .Y(_0081_));
 sky130_fd_sc_hd__xnor2_1 _0889_ (.A(\lfsr_reg[28] ),
    .B(\lfsr_reg[15] ),
    .Y(_0337_));
 sky130_fd_sc_hd__nand2_1 _0890_ (.A(_0326_),
    .B(_0337_),
    .Y(_0338_));
 sky130_fd_sc_hd__o21ai_0 _0891_ (.A1(_0326_),
    .A2(\lfsr_reg[16] ),
    .B1(_0338_),
    .Y(_0339_));
 sky130_fd_sc_hd__nand2_1 _0892_ (.A(_0324_),
    .B(_0339_),
    .Y(_0082_));
 sky130_fd_sc_hd__mux2i_1 _0893_ (.A0(\lfsr_reg[17] ),
    .A1(\lfsr_reg[16] ),
    .S(_0304_),
    .Y(_0340_));
 sky130_fd_sc_hd__nor2_1 _0894_ (.A(_0000_),
    .B(_0340_),
    .Y(_0083_));
 sky130_fd_sc_hd__mux2i_1 _0895_ (.A0(\lfsr_reg[18] ),
    .A1(\lfsr_reg[17] ),
    .S(_0333_),
    .Y(_0341_));
 sky130_fd_sc_hd__nand2_1 _0896_ (.A(_0324_),
    .B(_0341_),
    .Y(_0084_));
 sky130_fd_sc_hd__mux2i_1 _0897_ (.A0(\lfsr_reg[19] ),
    .A1(\lfsr_reg[18] ),
    .S(_0333_),
    .Y(_0342_));
 sky130_fd_sc_hd__nand2_1 _0898_ (.A(_0324_),
    .B(_0342_),
    .Y(_0085_));
 sky130_fd_sc_hd__mux2i_1 _0899_ (.A0(\lfsr_reg[1] ),
    .A1(\lfsr_reg[0] ),
    .S(_0304_),
    .Y(_0343_));
 sky130_fd_sc_hd__nor2_1 _0900_ (.A(_0000_),
    .B(_0343_),
    .Y(_0086_));
 sky130_fd_sc_hd__mux2i_1 _0901_ (.A0(\lfsr_reg[20] ),
    .A1(\lfsr_reg[19] ),
    .S(_0304_),
    .Y(_0344_));
 sky130_fd_sc_hd__nor2_1 _0902_ (.A(_0000_),
    .B(_0344_),
    .Y(_0087_));
 sky130_fd_sc_hd__mux2i_1 _0903_ (.A0(\lfsr_reg[21] ),
    .A1(\lfsr_reg[20] ),
    .S(_0304_),
    .Y(_0345_));
 sky130_fd_sc_hd__nor2_1 _0904_ (.A(_0000_),
    .B(_0345_),
    .Y(_0088_));
 sky130_fd_sc_hd__mux2i_1 _0905_ (.A0(\lfsr_reg[22] ),
    .A1(\lfsr_reg[21] ),
    .S(_0333_),
    .Y(_0346_));
 sky130_fd_sc_hd__nand2_1 _0906_ (.A(_0324_),
    .B(_0346_),
    .Y(_0089_));
 sky130_fd_sc_hd__mux2i_1 _0907_ (.A0(\lfsr_reg[23] ),
    .A1(\lfsr_reg[22] ),
    .S(_0333_),
    .Y(_0347_));
 sky130_fd_sc_hd__nand2_1 _0908_ (.A(_0324_),
    .B(_0347_),
    .Y(_0090_));
 sky130_fd_sc_hd__mux2i_1 _0909_ (.A0(\lfsr_reg[24] ),
    .A1(\lfsr_reg[23] ),
    .S(_0333_),
    .Y(_0348_));
 sky130_fd_sc_hd__nand2_1 _0910_ (.A(_0151_),
    .B(_0348_),
    .Y(_0091_));
 sky130_fd_sc_hd__mux2i_1 _0911_ (.A0(\lfsr_reg[25] ),
    .A1(\lfsr_reg[24] ),
    .S(_0333_),
    .Y(_0349_));
 sky130_fd_sc_hd__nand2_1 _0912_ (.A(_0151_),
    .B(_0349_),
    .Y(_0092_));
 sky130_fd_sc_hd__mux2i_1 _0913_ (.A0(\lfsr_reg[26] ),
    .A1(\lfsr_reg[25] ),
    .S(_0304_),
    .Y(_0350_));
 sky130_fd_sc_hd__nor2_1 _0914_ (.A(_0237_),
    .B(_0350_),
    .Y(_0093_));
 sky130_fd_sc_hd__xnor2_1 _0915_ (.A(_0325_),
    .B(\lfsr_reg[26] ),
    .Y(_0351_));
 sky130_fd_sc_hd__nand2_1 _0916_ (.A(_0326_),
    .B(_0351_),
    .Y(_0352_));
 sky130_fd_sc_hd__o21ai_0 _0917_ (.A1(_0326_),
    .A2(\lfsr_reg[27] ),
    .B1(_0352_),
    .Y(_0353_));
 sky130_fd_sc_hd__nand2_1 _0918_ (.A(_0151_),
    .B(_0353_),
    .Y(_0094_));
 sky130_fd_sc_hd__buf_4 _0919_ (.A(_0152_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2i_1 _0920_ (.A0(\lfsr_reg[28] ),
    .A1(\lfsr_reg[27] ),
    .S(_0354_),
    .Y(_0355_));
 sky130_fd_sc_hd__nor2_1 _0921_ (.A(_0237_),
    .B(_0355_),
    .Y(_0095_));
 sky130_fd_sc_hd__xor2_1 _0922_ (.A(_0325_),
    .B(\lfsr_reg[28] ),
    .X(_0356_));
 sky130_fd_sc_hd__a21oi_1 _0923_ (.A1(_0354_),
    .A2(_0356_),
    .B1(\lfsr_reg[29] ),
    .Y(_0357_));
 sky130_fd_sc_hd__and3_1 _0924_ (.A(_0354_),
    .B(\lfsr_reg[29] ),
    .C(_0356_),
    .X(_0358_));
 sky130_fd_sc_hd__buf_2 _0925_ (.A(_0145_),
    .X(_0359_));
 sky130_fd_sc_hd__o21ai_0 _0926_ (.A1(_0357_),
    .A2(_0358_),
    .B1(_0359_),
    .Y(_0096_));
 sky130_fd_sc_hd__mux2i_1 _0927_ (.A0(\lfsr_reg[2] ),
    .A1(\lfsr_reg[1] ),
    .S(_0354_),
    .Y(_0360_));
 sky130_fd_sc_hd__nor2_1 _0928_ (.A(_0237_),
    .B(_0360_),
    .Y(_0097_));
 sky130_fd_sc_hd__nand2_1 _0929_ (.A(_0354_),
    .B(\lfsr_reg[29] ),
    .Y(_0361_));
 sky130_fd_sc_hd__xor2_1 _0930_ (.A(\lfsr_reg[30] ),
    .B(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__nor2_1 _0931_ (.A(_0237_),
    .B(_0362_),
    .Y(_0098_));
 sky130_fd_sc_hd__a21oi_1 _0932_ (.A1(_0354_),
    .A2(\lfsr_reg[30] ),
    .B1(_0325_),
    .Y(_0363_));
 sky130_fd_sc_hd__and3_1 _0933_ (.A(_0354_),
    .B(\lfsr_reg[30] ),
    .C(_0325_),
    .X(_0364_));
 sky130_fd_sc_hd__o21ai_0 _0934_ (.A1(_0363_),
    .A2(_0364_),
    .B1(_0359_),
    .Y(_0099_));
 sky130_fd_sc_hd__mux2i_1 _0935_ (.A0(\lfsr_reg[3] ),
    .A1(\lfsr_reg[2] ),
    .S(_0354_),
    .Y(_0365_));
 sky130_fd_sc_hd__nor2_1 _0936_ (.A(_0237_),
    .B(_0365_),
    .Y(_0100_));
 sky130_fd_sc_hd__mux2i_1 _0937_ (.A0(\lfsr_reg[4] ),
    .A1(\lfsr_reg[3] ),
    .S(_0333_),
    .Y(_0366_));
 sky130_fd_sc_hd__nand2_1 _0938_ (.A(_0151_),
    .B(_0366_),
    .Y(_0101_));
 sky130_fd_sc_hd__xnor2_1 _0939_ (.A(\lfsr_reg[29] ),
    .B(\lfsr_reg[4] ),
    .Y(_0367_));
 sky130_fd_sc_hd__nand2_1 _0940_ (.A(_0326_),
    .B(_0367_),
    .Y(_0368_));
 sky130_fd_sc_hd__o21ai_0 _0941_ (.A1(_0326_),
    .A2(\lfsr_reg[5] ),
    .B1(_0368_),
    .Y(_0369_));
 sky130_fd_sc_hd__nand2_1 _0942_ (.A(_0151_),
    .B(_0369_),
    .Y(_0102_));
 sky130_fd_sc_hd__mux2i_1 _0943_ (.A0(\lfsr_reg[6] ),
    .A1(\lfsr_reg[5] ),
    .S(_0304_),
    .Y(_0370_));
 sky130_fd_sc_hd__nand2_1 _0944_ (.A(_0151_),
    .B(_0370_),
    .Y(_0103_));
 sky130_fd_sc_hd__mux2i_1 _0945_ (.A0(\lfsr_reg[7] ),
    .A1(\lfsr_reg[6] ),
    .S(_0354_),
    .Y(_0371_));
 sky130_fd_sc_hd__nor2_1 _0946_ (.A(_0237_),
    .B(_0371_),
    .Y(_0104_));
 sky130_fd_sc_hd__mux2i_1 _0947_ (.A0(\lfsr_reg[8] ),
    .A1(\lfsr_reg[7] ),
    .S(_0304_),
    .Y(_0372_));
 sky130_fd_sc_hd__nand2_1 _0948_ (.A(_0151_),
    .B(_0372_),
    .Y(_0105_));
 sky130_fd_sc_hd__mux2i_1 _0949_ (.A0(\lfsr_reg[9] ),
    .A1(\lfsr_reg[8] ),
    .S(_0354_),
    .Y(_0373_));
 sky130_fd_sc_hd__nor2_1 _0950_ (.A(_0237_),
    .B(_0373_),
    .Y(_0106_));
 sky130_fd_sc_hd__clkbuf_2 _0951_ (.A(_0148_),
    .X(_0374_));
 sky130_fd_sc_hd__xnor2_2 _0952_ (.A(\entropy_pool[0] ),
    .B(\entropy_pool[24] ),
    .Y(_0375_));
 sky130_fd_sc_hd__xnor2_2 _0953_ (.A(\lfsr_reg[0] ),
    .B(\lfsr_reg[16] ),
    .Y(_0376_));
 sky130_fd_sc_hd__xnor2_1 _0954_ (.A(\entropy_pool2[0] ),
    .B(_0376_),
    .Y(_0377_));
 sky130_fd_sc_hd__or3_1 _0955_ (.A(_0374_),
    .B(_0375_),
    .C(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__nand3_1 _0956_ (.A(_0001_),
    .B(_0375_),
    .C(_0377_),
    .Y(_0379_));
 sky130_fd_sc_hd__buf_2 _0957_ (.A(_0145_),
    .X(_0380_));
 sky130_fd_sc_hd__nand2b_2 _0958_ (.A_N(\state[0] ),
    .B(\state[1] ),
    .Y(_0381_));
 sky130_fd_sc_hd__buf_2 _0959_ (.A(_0381_),
    .X(_0382_));
 sky130_fd_sc_hd__nand3_1 _0960_ (.A(_0380_),
    .B(\mixed_output[0] ),
    .C(_0382_),
    .Y(_0383_));
 sky130_fd_sc_hd__nand3_1 _0961_ (.A(_0378_),
    .B(_0379_),
    .C(_0383_),
    .Y(_0107_));
 sky130_fd_sc_hd__xnor2_2 _0962_ (.A(\lfsr_reg[10] ),
    .B(\lfsr_reg[26] ),
    .Y(_0384_));
 sky130_fd_sc_hd__xnor2_2 _0963_ (.A(\entropy_pool[10] ),
    .B(\entropy_pool[18] ),
    .Y(_0385_));
 sky130_fd_sc_hd__xnor2_1 _0964_ (.A(\entropy_pool2[10] ),
    .B(_0385_),
    .Y(_0386_));
 sky130_fd_sc_hd__or3_1 _0965_ (.A(_0374_),
    .B(_0384_),
    .C(_0386_),
    .X(_0387_));
 sky130_fd_sc_hd__nand3_1 _0966_ (.A(_0001_),
    .B(_0384_),
    .C(_0386_),
    .Y(_0388_));
 sky130_fd_sc_hd__nand3_1 _0967_ (.A(_0380_),
    .B(\mixed_output[10] ),
    .C(_0382_),
    .Y(_0389_));
 sky130_fd_sc_hd__nand3_1 _0968_ (.A(_0387_),
    .B(_0388_),
    .C(_0389_),
    .Y(_0108_));
 sky130_fd_sc_hd__buf_2 _0969_ (.A(_0148_),
    .X(_0390_));
 sky130_fd_sc_hd__xnor2_2 _0970_ (.A(\entropy_pool[11] ),
    .B(\entropy_pool[19] ),
    .Y(_0391_));
 sky130_fd_sc_hd__nor2_1 _0971_ (.A(_0390_),
    .B(_0391_),
    .Y(_0392_));
 sky130_fd_sc_hd__buf_2 _0972_ (.A(_0148_),
    .X(_0393_));
 sky130_fd_sc_hd__nor2b_1 _0973_ (.A(_0393_),
    .B_N(_0391_),
    .Y(_0394_));
 sky130_fd_sc_hd__xor2_2 _0974_ (.A(\lfsr_reg[11] ),
    .B(\lfsr_reg[27] ),
    .X(_0395_));
 sky130_fd_sc_hd__xor2_1 _0975_ (.A(\entropy_pool2[11] ),
    .B(_0395_),
    .X(_0396_));
 sky130_fd_sc_hd__mux2i_1 _0976_ (.A0(_0392_),
    .A1(_0394_),
    .S(_0396_),
    .Y(_0397_));
 sky130_fd_sc_hd__buf_2 _0977_ (.A(_0381_),
    .X(_0398_));
 sky130_fd_sc_hd__nand3_1 _0978_ (.A(_0359_),
    .B(\mixed_output[11] ),
    .C(_0398_),
    .Y(_0399_));
 sky130_fd_sc_hd__nand2_1 _0979_ (.A(_0397_),
    .B(_0399_),
    .Y(_0109_));
 sky130_fd_sc_hd__xnor2_2 _0980_ (.A(\entropy_pool[12] ),
    .B(\entropy_pool[20] ),
    .Y(_0400_));
 sky130_fd_sc_hd__nor2_1 _0981_ (.A(_0390_),
    .B(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__nor2b_1 _0982_ (.A(_0393_),
    .B_N(_0400_),
    .Y(_0402_));
 sky130_fd_sc_hd__xor2_4 _0983_ (.A(\lfsr_reg[12] ),
    .B(\lfsr_reg[28] ),
    .X(_0403_));
 sky130_fd_sc_hd__xor2_1 _0984_ (.A(\entropy_pool2[12] ),
    .B(_0403_),
    .X(_0404_));
 sky130_fd_sc_hd__mux2i_1 _0985_ (.A0(_0401_),
    .A1(_0402_),
    .S(_0404_),
    .Y(_0405_));
 sky130_fd_sc_hd__nand3_1 _0986_ (.A(_0359_),
    .B(\mixed_output[12] ),
    .C(_0398_),
    .Y(_0406_));
 sky130_fd_sc_hd__nand2_1 _0987_ (.A(_0405_),
    .B(_0406_),
    .Y(_0110_));
 sky130_fd_sc_hd__xnor2_2 _0988_ (.A(\lfsr_reg[29] ),
    .B(\lfsr_reg[13] ),
    .Y(_0407_));
 sky130_fd_sc_hd__xnor2_2 _0989_ (.A(\entropy_pool[13] ),
    .B(\entropy_pool[21] ),
    .Y(_0408_));
 sky130_fd_sc_hd__xnor2_1 _0990_ (.A(\entropy_pool2[13] ),
    .B(_0408_),
    .Y(_0409_));
 sky130_fd_sc_hd__or3_1 _0991_ (.A(_0374_),
    .B(_0407_),
    .C(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__nand3_1 _0992_ (.A(_0001_),
    .B(_0407_),
    .C(_0409_),
    .Y(_0411_));
 sky130_fd_sc_hd__nand3_1 _0993_ (.A(_0380_),
    .B(\mixed_output[13] ),
    .C(_0382_),
    .Y(_0412_));
 sky130_fd_sc_hd__nand3_1 _0994_ (.A(_0410_),
    .B(_0411_),
    .C(_0412_),
    .Y(_0111_));
 sky130_fd_sc_hd__xnor2_2 _0995_ (.A(\lfsr_reg[30] ),
    .B(\lfsr_reg[14] ),
    .Y(_0413_));
 sky130_fd_sc_hd__xnor2_2 _0996_ (.A(\entropy_pool[14] ),
    .B(\entropy_pool[22] ),
    .Y(_0414_));
 sky130_fd_sc_hd__xnor2_1 _0997_ (.A(\entropy_pool2[14] ),
    .B(_0414_),
    .Y(_0415_));
 sky130_fd_sc_hd__or3_1 _0998_ (.A(_0374_),
    .B(_0413_),
    .C(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__nand3_1 _0999_ (.A(_0001_),
    .B(_0413_),
    .C(_0415_),
    .Y(_0417_));
 sky130_fd_sc_hd__nand3_1 _1000_ (.A(_0380_),
    .B(\mixed_output[14] ),
    .C(_0382_),
    .Y(_0418_));
 sky130_fd_sc_hd__nand3_1 _1001_ (.A(_0416_),
    .B(_0417_),
    .C(_0418_),
    .Y(_0112_));
 sky130_fd_sc_hd__xnor2_2 _1002_ (.A(_0325_),
    .B(\lfsr_reg[15] ),
    .Y(_0419_));
 sky130_fd_sc_hd__xnor2_2 _1003_ (.A(\entropy_pool[15] ),
    .B(\entropy_pool[23] ),
    .Y(_0420_));
 sky130_fd_sc_hd__xnor2_1 _1004_ (.A(\entropy_pool2[15] ),
    .B(_0420_),
    .Y(_0421_));
 sky130_fd_sc_hd__or3_1 _1005_ (.A(_0374_),
    .B(_0419_),
    .C(_0421_),
    .X(_0422_));
 sky130_fd_sc_hd__nand3_1 _1006_ (.A(_0001_),
    .B(_0419_),
    .C(_0421_),
    .Y(_0423_));
 sky130_fd_sc_hd__nand3_1 _1007_ (.A(_0380_),
    .B(\mixed_output[15] ),
    .C(_0382_),
    .Y(_0424_));
 sky130_fd_sc_hd__nand3_1 _1008_ (.A(_0422_),
    .B(_0423_),
    .C(_0424_),
    .Y(_0113_));
 sky130_fd_sc_hd__xnor2_2 _1009_ (.A(\entropy_pool[8] ),
    .B(\entropy_pool[16] ),
    .Y(_0425_));
 sky130_fd_sc_hd__xnor2_1 _1010_ (.A(\entropy_pool2[16] ),
    .B(_0425_),
    .Y(_0426_));
 sky130_fd_sc_hd__or3_1 _1011_ (.A(_0374_),
    .B(_0376_),
    .C(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__nand3_1 _1012_ (.A(_0001_),
    .B(_0376_),
    .C(_0426_),
    .Y(_0428_));
 sky130_fd_sc_hd__nand3_1 _1013_ (.A(_0380_),
    .B(\mixed_output[16] ),
    .C(_0382_),
    .Y(_0429_));
 sky130_fd_sc_hd__nand3_1 _1014_ (.A(_0427_),
    .B(_0428_),
    .C(_0429_),
    .Y(_0114_));
 sky130_fd_sc_hd__xnor2_2 _1015_ (.A(\lfsr_reg[1] ),
    .B(\lfsr_reg[17] ),
    .Y(_0430_));
 sky130_fd_sc_hd__xnor2_2 _1016_ (.A(\entropy_pool[9] ),
    .B(\entropy_pool[17] ),
    .Y(_0431_));
 sky130_fd_sc_hd__xnor2_1 _1017_ (.A(\entropy_pool2[17] ),
    .B(_0431_),
    .Y(_0432_));
 sky130_fd_sc_hd__or3_1 _1018_ (.A(_0374_),
    .B(_0430_),
    .C(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__nand3_1 _1019_ (.A(_0001_),
    .B(_0430_),
    .C(_0432_),
    .Y(_0434_));
 sky130_fd_sc_hd__nand3_1 _1020_ (.A(_0380_),
    .B(\mixed_output[17] ),
    .C(_0382_),
    .Y(_0435_));
 sky130_fd_sc_hd__nand3_1 _1021_ (.A(_0433_),
    .B(_0434_),
    .C(_0435_),
    .Y(_0115_));
 sky130_fd_sc_hd__xnor2_2 _1022_ (.A(\lfsr_reg[2] ),
    .B(\lfsr_reg[18] ),
    .Y(_0436_));
 sky130_fd_sc_hd__xnor2_1 _1023_ (.A(\entropy_pool2[18] ),
    .B(_0436_),
    .Y(_0437_));
 sky130_fd_sc_hd__or3_1 _1024_ (.A(_0374_),
    .B(_0385_),
    .C(_0437_),
    .X(_0438_));
 sky130_fd_sc_hd__nand3_1 _1025_ (.A(_0001_),
    .B(_0385_),
    .C(_0437_),
    .Y(_0439_));
 sky130_fd_sc_hd__nand3_1 _1026_ (.A(_0380_),
    .B(\mixed_output[18] ),
    .C(_0382_),
    .Y(_0440_));
 sky130_fd_sc_hd__nand3_1 _1027_ (.A(_0438_),
    .B(_0439_),
    .C(_0440_),
    .Y(_0116_));
 sky130_fd_sc_hd__xor2_4 _1028_ (.A(\lfsr_reg[3] ),
    .B(\lfsr_reg[19] ),
    .X(_0441_));
 sky130_fd_sc_hd__xor2_1 _1029_ (.A(\entropy_pool2[19] ),
    .B(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__mux2i_2 _1030_ (.A0(_0392_),
    .A1(_0394_),
    .S(_0442_),
    .Y(_0443_));
 sky130_fd_sc_hd__nand3_1 _1031_ (.A(_0359_),
    .B(\mixed_output[19] ),
    .C(_0398_),
    .Y(_0444_));
 sky130_fd_sc_hd__nand2_1 _1032_ (.A(_0443_),
    .B(_0444_),
    .Y(_0117_));
 sky130_fd_sc_hd__xnor2_2 _1033_ (.A(\entropy_pool[1] ),
    .B(\entropy_pool[25] ),
    .Y(_0445_));
 sky130_fd_sc_hd__xnor2_1 _1034_ (.A(\entropy_pool2[1] ),
    .B(_0430_),
    .Y(_0446_));
 sky130_fd_sc_hd__or3_1 _1035_ (.A(_0374_),
    .B(_0445_),
    .C(_0446_),
    .X(_0447_));
 sky130_fd_sc_hd__nand3_1 _1036_ (.A(_0001_),
    .B(_0445_),
    .C(_0446_),
    .Y(_0448_));
 sky130_fd_sc_hd__nand3_1 _1037_ (.A(_0150_),
    .B(\mixed_output[1] ),
    .C(_0382_),
    .Y(_0449_));
 sky130_fd_sc_hd__nand3_1 _1038_ (.A(_0447_),
    .B(_0448_),
    .C(_0449_),
    .Y(_0118_));
 sky130_fd_sc_hd__xor2_4 _1039_ (.A(\lfsr_reg[4] ),
    .B(\lfsr_reg[20] ),
    .X(_0450_));
 sky130_fd_sc_hd__xor2_1 _1040_ (.A(\entropy_pool2[20] ),
    .B(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__mux2i_2 _1041_ (.A0(_0401_),
    .A1(_0402_),
    .S(_0451_),
    .Y(_0452_));
 sky130_fd_sc_hd__nand3_1 _1042_ (.A(_0359_),
    .B(\mixed_output[20] ),
    .C(_0398_),
    .Y(_0453_));
 sky130_fd_sc_hd__nand2_1 _1043_ (.A(_0452_),
    .B(_0453_),
    .Y(_0119_));
 sky130_fd_sc_hd__xnor2_2 _1044_ (.A(\lfsr_reg[5] ),
    .B(\lfsr_reg[21] ),
    .Y(_0454_));
 sky130_fd_sc_hd__xnor2_1 _1045_ (.A(\entropy_pool2[21] ),
    .B(_0454_),
    .Y(_0455_));
 sky130_fd_sc_hd__or3_1 _1046_ (.A(_0374_),
    .B(_0408_),
    .C(_0455_),
    .X(_0456_));
 sky130_fd_sc_hd__nand3_1 _1047_ (.A(_0149_),
    .B(_0408_),
    .C(_0455_),
    .Y(_0457_));
 sky130_fd_sc_hd__nand3_1 _1048_ (.A(_0150_),
    .B(\mixed_output[21] ),
    .C(_0382_),
    .Y(_0458_));
 sky130_fd_sc_hd__nand3_1 _1049_ (.A(_0456_),
    .B(_0457_),
    .C(_0458_),
    .Y(_0120_));
 sky130_fd_sc_hd__xnor2_2 _1050_ (.A(\lfsr_reg[6] ),
    .B(\lfsr_reg[22] ),
    .Y(_0459_));
 sky130_fd_sc_hd__xnor2_1 _1051_ (.A(\entropy_pool2[22] ),
    .B(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__or3_1 _1052_ (.A(_0393_),
    .B(_0414_),
    .C(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__nand3_1 _1053_ (.A(_0149_),
    .B(_0414_),
    .C(_0460_),
    .Y(_0462_));
 sky130_fd_sc_hd__nand3_1 _1054_ (.A(_0150_),
    .B(\mixed_output[22] ),
    .C(_0381_),
    .Y(_0463_));
 sky130_fd_sc_hd__nand3_1 _1055_ (.A(_0461_),
    .B(_0462_),
    .C(_0463_),
    .Y(_0121_));
 sky130_fd_sc_hd__xnor2_2 _1056_ (.A(\lfsr_reg[7] ),
    .B(\lfsr_reg[23] ),
    .Y(_0464_));
 sky130_fd_sc_hd__xnor2_1 _1057_ (.A(\entropy_pool2[23] ),
    .B(_0420_),
    .Y(_0465_));
 sky130_fd_sc_hd__or3_1 _1058_ (.A(_0393_),
    .B(_0464_),
    .C(_0465_),
    .X(_0466_));
 sky130_fd_sc_hd__nand3_1 _1059_ (.A(_0149_),
    .B(_0464_),
    .C(_0465_),
    .Y(_0467_));
 sky130_fd_sc_hd__nand3_1 _1060_ (.A(_0150_),
    .B(\mixed_output[23] ),
    .C(_0381_),
    .Y(_0468_));
 sky130_fd_sc_hd__nand3_1 _1061_ (.A(_0466_),
    .B(_0467_),
    .C(_0468_),
    .Y(_0122_));
 sky130_fd_sc_hd__xnor2_1 _1062_ (.A(\lfsr_reg[8] ),
    .B(\lfsr_reg[24] ),
    .Y(_0469_));
 sky130_fd_sc_hd__nor2_1 _1063_ (.A(_0390_),
    .B(_0469_),
    .Y(_0470_));
 sky130_fd_sc_hd__nor2b_1 _1064_ (.A(_0393_),
    .B_N(_0469_),
    .Y(_0471_));
 sky130_fd_sc_hd__xnor2_1 _1065_ (.A(\entropy_pool2[24] ),
    .B(_0375_),
    .Y(_0472_));
 sky130_fd_sc_hd__mux2i_2 _1066_ (.A0(_0470_),
    .A1(_0471_),
    .S(_0472_),
    .Y(_0473_));
 sky130_fd_sc_hd__nand3_1 _1067_ (.A(_0359_),
    .B(\mixed_output[24] ),
    .C(_0398_),
    .Y(_0474_));
 sky130_fd_sc_hd__nand2_1 _1068_ (.A(_0473_),
    .B(_0474_),
    .Y(_0123_));
 sky130_fd_sc_hd__xnor2_1 _1069_ (.A(\lfsr_reg[9] ),
    .B(\lfsr_reg[25] ),
    .Y(_0475_));
 sky130_fd_sc_hd__nor2_1 _1070_ (.A(_0390_),
    .B(_0475_),
    .Y(_0476_));
 sky130_fd_sc_hd__nor2b_1 _1071_ (.A(_0393_),
    .B_N(_0475_),
    .Y(_0477_));
 sky130_fd_sc_hd__xnor2_1 _1072_ (.A(\entropy_pool2[25] ),
    .B(_0445_),
    .Y(_0478_));
 sky130_fd_sc_hd__mux2i_1 _1073_ (.A0(_0476_),
    .A1(_0477_),
    .S(_0478_),
    .Y(_0479_));
 sky130_fd_sc_hd__nand3_1 _1074_ (.A(_0359_),
    .B(\mixed_output[25] ),
    .C(_0398_),
    .Y(_0480_));
 sky130_fd_sc_hd__nand2_1 _1075_ (.A(_0479_),
    .B(_0480_),
    .Y(_0124_));
 sky130_fd_sc_hd__xnor2_1 _1076_ (.A(\entropy_pool[2] ),
    .B(\entropy_pool[26] ),
    .Y(_0481_));
 sky130_fd_sc_hd__nor2_1 _1077_ (.A(_0390_),
    .B(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__nor2b_1 _1078_ (.A(_0393_),
    .B_N(_0481_),
    .Y(_0483_));
 sky130_fd_sc_hd__xnor2_1 _1079_ (.A(\entropy_pool2[26] ),
    .B(_0384_),
    .Y(_0484_));
 sky130_fd_sc_hd__mux2i_1 _1080_ (.A0(_0482_),
    .A1(_0483_),
    .S(_0484_),
    .Y(_0485_));
 sky130_fd_sc_hd__nand3_1 _1081_ (.A(_0359_),
    .B(\mixed_output[26] ),
    .C(_0398_),
    .Y(_0486_));
 sky130_fd_sc_hd__nand2_1 _1082_ (.A(_0485_),
    .B(_0486_),
    .Y(_0125_));
 sky130_fd_sc_hd__xnor2_1 _1083_ (.A(\entropy_pool[3] ),
    .B(\entropy_pool[27] ),
    .Y(_0487_));
 sky130_fd_sc_hd__nor2_1 _1084_ (.A(_0390_),
    .B(_0487_),
    .Y(_0488_));
 sky130_fd_sc_hd__nor2b_1 _1085_ (.A(_0393_),
    .B_N(_0487_),
    .Y(_0489_));
 sky130_fd_sc_hd__xor2_1 _1086_ (.A(\entropy_pool2[27] ),
    .B(_0395_),
    .X(_0490_));
 sky130_fd_sc_hd__mux2i_2 _1087_ (.A0(_0488_),
    .A1(_0489_),
    .S(_0490_),
    .Y(_0491_));
 sky130_fd_sc_hd__nand3_1 _1088_ (.A(_0359_),
    .B(\mixed_output[27] ),
    .C(_0398_),
    .Y(_0492_));
 sky130_fd_sc_hd__nand2_1 _1089_ (.A(_0491_),
    .B(_0492_),
    .Y(_0126_));
 sky130_fd_sc_hd__xnor2_1 _1090_ (.A(\entropy_pool[4] ),
    .B(\entropy_pool[28] ),
    .Y(_0493_));
 sky130_fd_sc_hd__nor2_1 _1091_ (.A(_0390_),
    .B(_0493_),
    .Y(_0494_));
 sky130_fd_sc_hd__nor2b_1 _1092_ (.A(_0393_),
    .B_N(_0493_),
    .Y(_0495_));
 sky130_fd_sc_hd__xor2_1 _1093_ (.A(\entropy_pool2[28] ),
    .B(_0403_),
    .X(_0496_));
 sky130_fd_sc_hd__mux2i_2 _1094_ (.A0(_0494_),
    .A1(_0495_),
    .S(_0496_),
    .Y(_0497_));
 sky130_fd_sc_hd__buf_2 _1095_ (.A(_0145_),
    .X(_0498_));
 sky130_fd_sc_hd__nand3_1 _1096_ (.A(_0498_),
    .B(\mixed_output[28] ),
    .C(_0398_),
    .Y(_0499_));
 sky130_fd_sc_hd__nand2_1 _1097_ (.A(_0497_),
    .B(_0499_),
    .Y(_0127_));
 sky130_fd_sc_hd__xnor2_1 _1098_ (.A(\entropy_pool[5] ),
    .B(\entropy_pool[29] ),
    .Y(_0500_));
 sky130_fd_sc_hd__nor2_1 _1099_ (.A(_0390_),
    .B(_0500_),
    .Y(_0501_));
 sky130_fd_sc_hd__nor2b_1 _1100_ (.A(_0393_),
    .B_N(_0500_),
    .Y(_0502_));
 sky130_fd_sc_hd__xnor2_1 _1101_ (.A(\entropy_pool2[29] ),
    .B(_0407_),
    .Y(_0503_));
 sky130_fd_sc_hd__mux2i_1 _1102_ (.A0(_0501_),
    .A1(_0502_),
    .S(_0503_),
    .Y(_0504_));
 sky130_fd_sc_hd__nand3_1 _1103_ (.A(_0498_),
    .B(\mixed_output[29] ),
    .C(_0398_),
    .Y(_0505_));
 sky130_fd_sc_hd__nand2_1 _1104_ (.A(_0504_),
    .B(_0505_),
    .Y(_0128_));
 sky130_fd_sc_hd__xnor2_1 _1105_ (.A(\entropy_pool2[2] ),
    .B(_0436_),
    .Y(_0506_));
 sky130_fd_sc_hd__mux2i_1 _1106_ (.A0(_0482_),
    .A1(_0483_),
    .S(_0506_),
    .Y(_0507_));
 sky130_fd_sc_hd__buf_2 _1107_ (.A(_0381_),
    .X(_0508_));
 sky130_fd_sc_hd__nand3_1 _1108_ (.A(_0498_),
    .B(\mixed_output[2] ),
    .C(_0508_),
    .Y(_0509_));
 sky130_fd_sc_hd__nand2_1 _1109_ (.A(_0507_),
    .B(_0509_),
    .Y(_0129_));
 sky130_fd_sc_hd__xnor2_1 _1110_ (.A(\entropy_pool[6] ),
    .B(\entropy_pool[30] ),
    .Y(_0510_));
 sky130_fd_sc_hd__nor2_1 _1111_ (.A(_0390_),
    .B(_0510_),
    .Y(_0511_));
 sky130_fd_sc_hd__nor2b_1 _1112_ (.A(_0148_),
    .B_N(_0510_),
    .Y(_0512_));
 sky130_fd_sc_hd__xnor2_1 _1113_ (.A(\entropy_pool2[30] ),
    .B(_0413_),
    .Y(_0513_));
 sky130_fd_sc_hd__mux2i_1 _1114_ (.A0(_0511_),
    .A1(_0512_),
    .S(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__nand3_1 _1115_ (.A(_0498_),
    .B(\mixed_output[30] ),
    .C(_0508_),
    .Y(_0515_));
 sky130_fd_sc_hd__nand2_1 _1116_ (.A(_0514_),
    .B(_0515_),
    .Y(_0130_));
 sky130_fd_sc_hd__xnor2_1 _1117_ (.A(\entropy_pool[7] ),
    .B(\entropy_pool[31] ),
    .Y(_0516_));
 sky130_fd_sc_hd__nor2_1 _1118_ (.A(_0390_),
    .B(_0516_),
    .Y(_0517_));
 sky130_fd_sc_hd__nor2b_1 _1119_ (.A(_0148_),
    .B_N(_0516_),
    .Y(_0518_));
 sky130_fd_sc_hd__xnor2_1 _1120_ (.A(\entropy_pool2[31] ),
    .B(_0419_),
    .Y(_0519_));
 sky130_fd_sc_hd__mux2i_1 _1121_ (.A0(_0517_),
    .A1(_0518_),
    .S(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__nand3_1 _1122_ (.A(_0498_),
    .B(\mixed_output[31] ),
    .C(_0508_),
    .Y(_0521_));
 sky130_fd_sc_hd__nand2_1 _1123_ (.A(_0520_),
    .B(_0521_),
    .Y(_0131_));
 sky130_fd_sc_hd__xor2_1 _1124_ (.A(\entropy_pool2[3] ),
    .B(_0441_),
    .X(_0522_));
 sky130_fd_sc_hd__mux2i_1 _1125_ (.A0(_0488_),
    .A1(_0489_),
    .S(_0522_),
    .Y(_0523_));
 sky130_fd_sc_hd__nand3_1 _1126_ (.A(_0498_),
    .B(\mixed_output[3] ),
    .C(_0508_),
    .Y(_0524_));
 sky130_fd_sc_hd__nand2_1 _1127_ (.A(_0523_),
    .B(_0524_),
    .Y(_0132_));
 sky130_fd_sc_hd__xor2_1 _1128_ (.A(\entropy_pool2[4] ),
    .B(_0450_),
    .X(_0525_));
 sky130_fd_sc_hd__mux2i_1 _1129_ (.A0(_0494_),
    .A1(_0495_),
    .S(_0525_),
    .Y(_0526_));
 sky130_fd_sc_hd__nand3_1 _1130_ (.A(_0498_),
    .B(\mixed_output[4] ),
    .C(_0508_),
    .Y(_0527_));
 sky130_fd_sc_hd__nand2_1 _1131_ (.A(_0526_),
    .B(_0527_),
    .Y(_0133_));
 sky130_fd_sc_hd__xnor2_1 _1132_ (.A(\entropy_pool2[5] ),
    .B(_0454_),
    .Y(_0528_));
 sky130_fd_sc_hd__mux2i_1 _1133_ (.A0(_0501_),
    .A1(_0502_),
    .S(_0528_),
    .Y(_0529_));
 sky130_fd_sc_hd__nand3_1 _1134_ (.A(_0498_),
    .B(\mixed_output[5] ),
    .C(_0508_),
    .Y(_0530_));
 sky130_fd_sc_hd__nand2_1 _1135_ (.A(_0529_),
    .B(_0530_),
    .Y(_0134_));
 sky130_fd_sc_hd__xnor2_1 _1136_ (.A(\entropy_pool2[6] ),
    .B(_0459_),
    .Y(_0531_));
 sky130_fd_sc_hd__mux2i_1 _1137_ (.A0(_0511_),
    .A1(_0512_),
    .S(_0531_),
    .Y(_0532_));
 sky130_fd_sc_hd__nand3_1 _1138_ (.A(_0498_),
    .B(\mixed_output[6] ),
    .C(_0508_),
    .Y(_0533_));
 sky130_fd_sc_hd__nand2_1 _1139_ (.A(_0532_),
    .B(_0533_),
    .Y(_0135_));
 sky130_fd_sc_hd__xnor2_1 _1140_ (.A(\entropy_pool2[7] ),
    .B(_0464_),
    .Y(_0534_));
 sky130_fd_sc_hd__mux2i_1 _1141_ (.A0(_0517_),
    .A1(_0518_),
    .S(_0534_),
    .Y(_0535_));
 sky130_fd_sc_hd__nand3_1 _1142_ (.A(_0498_),
    .B(\mixed_output[7] ),
    .C(_0508_),
    .Y(_0536_));
 sky130_fd_sc_hd__nand2_1 _1143_ (.A(_0535_),
    .B(_0536_),
    .Y(_0136_));
 sky130_fd_sc_hd__xnor2_1 _1144_ (.A(\entropy_pool2[8] ),
    .B(_0425_),
    .Y(_0537_));
 sky130_fd_sc_hd__mux2i_1 _1145_ (.A0(_0470_),
    .A1(_0471_),
    .S(_0537_),
    .Y(_0538_));
 sky130_fd_sc_hd__nand3_1 _1146_ (.A(_0380_),
    .B(\mixed_output[8] ),
    .C(_0508_),
    .Y(_0539_));
 sky130_fd_sc_hd__nand2_1 _1147_ (.A(_0538_),
    .B(_0539_),
    .Y(_0137_));
 sky130_fd_sc_hd__xnor2_1 _1148_ (.A(\entropy_pool2[9] ),
    .B(_0431_),
    .Y(_0540_));
 sky130_fd_sc_hd__mux2i_1 _1149_ (.A0(_0476_),
    .A1(_0477_),
    .S(_0540_),
    .Y(_0541_));
 sky130_fd_sc_hd__nand3_1 _1150_ (.A(_0380_),
    .B(\mixed_output[9] ),
    .C(_0508_),
    .Y(_0542_));
 sky130_fd_sc_hd__nand2_1 _1151_ (.A(_0541_),
    .B(_0542_),
    .Y(_0138_));
 sky130_fd_sc_hd__nand2b_1 _1152_ (.A_N(\state[0] ),
    .B(net1),
    .Y(_0543_));
 sky130_fd_sc_hd__nand2_1 _1153_ (.A(_0326_),
    .B(_0150_),
    .Y(_0544_));
 sky130_fd_sc_hd__a21oi_1 _1154_ (.A1(_0306_),
    .A2(_0543_),
    .B1(_0544_),
    .Y(_0139_));
 sky130_fd_sc_hd__o31ai_1 _1155_ (.A1(_0306_),
    .A2(\health_counter[7] ),
    .A3(\health_counter[6] ),
    .B1(\state[0] ),
    .Y(_0545_));
 sky130_fd_sc_hd__nand2b_1 _1156_ (.A_N(net1),
    .B(_0306_),
    .Y(_0546_));
 sky130_fd_sc_hd__a21oi_1 _1157_ (.A1(_0545_),
    .A2(_0546_),
    .B1(_0544_),
    .Y(_0140_));
 sky130_fd_sc_hd__nor2_1 _1158_ (.A(\state[0] ),
    .B(_0306_),
    .Y(_0547_));
 sky130_fd_sc_hd__nor4_1 _1159_ (.A(\health_counter[7] ),
    .B(\health_counter[6] ),
    .C(\health_counter[5] ),
    .D(_0547_),
    .Y(net3));
 sky130_fd_sc_hd__nand4_1 _1160_ (.A(\mixed_output[13] ),
    .B(\mixed_output[14] ),
    .C(\mixed_output[15] ),
    .D(\mixed_output[16] ),
    .Y(_0548_));
 sky130_fd_sc_hd__nand4_1 _1161_ (.A(\mixed_output[0] ),
    .B(\mixed_output[10] ),
    .C(\mixed_output[11] ),
    .D(\mixed_output[12] ),
    .Y(_0549_));
 sky130_fd_sc_hd__nand4_1 _1162_ (.A(\mixed_output[3] ),
    .B(\mixed_output[7] ),
    .C(\mixed_output[8] ),
    .D(\mixed_output[9] ),
    .Y(_0550_));
 sky130_fd_sc_hd__nand4_1 _1163_ (.A(\mixed_output[24] ),
    .B(\mixed_output[4] ),
    .C(\mixed_output[5] ),
    .D(\mixed_output[6] ),
    .Y(_0551_));
 sky130_fd_sc_hd__or4_1 _1164_ (.A(_0548_),
    .B(_0549_),
    .C(_0550_),
    .D(_0551_),
    .X(_0552_));
 sky130_fd_sc_hd__nand4_1 _1165_ (.A(\mixed_output[17] ),
    .B(\mixed_output[20] ),
    .C(\mixed_output[21] ),
    .D(\mixed_output[22] ),
    .Y(_0553_));
 sky130_fd_sc_hd__nand4_1 _1166_ (.A(\mixed_output[18] ),
    .B(\mixed_output[19] ),
    .C(\mixed_output[1] ),
    .D(\mixed_output[23] ),
    .Y(_0554_));
 sky130_fd_sc_hd__nor3_1 _1167_ (.A(_0552_),
    .B(_0553_),
    .C(_0554_),
    .Y(_0555_));
 sky130_fd_sc_hd__nand3_1 _1168_ (.A(\mixed_output[25] ),
    .B(\mixed_output[26] ),
    .C(\mixed_output[27] ),
    .Y(_0556_));
 sky130_fd_sc_hd__nand4_1 _1169_ (.A(\mixed_output[28] ),
    .B(\mixed_output[29] ),
    .C(\mixed_output[30] ),
    .D(\mixed_output[31] ),
    .Y(_0557_));
 sky130_fd_sc_hd__nor2_1 _1170_ (.A(_0556_),
    .B(_0557_),
    .Y(_0558_));
 sky130_fd_sc_hd__nor4_1 _1171_ (.A(\mixed_output[24] ),
    .B(\mixed_output[29] ),
    .C(\mixed_output[2] ),
    .D(\mixed_output[30] ),
    .Y(_0559_));
 sky130_fd_sc_hd__nor4_1 _1172_ (.A(\mixed_output[25] ),
    .B(\mixed_output[26] ),
    .C(\mixed_output[27] ),
    .D(\mixed_output[28] ),
    .Y(_0560_));
 sky130_fd_sc_hd__nor4_1 _1173_ (.A(\mixed_output[31] ),
    .B(\mixed_output[7] ),
    .C(\mixed_output[8] ),
    .D(\mixed_output[9] ),
    .Y(_0561_));
 sky130_fd_sc_hd__nor4_1 _1174_ (.A(\mixed_output[3] ),
    .B(\mixed_output[4] ),
    .C(\mixed_output[5] ),
    .D(\mixed_output[6] ),
    .Y(_0562_));
 sky130_fd_sc_hd__nand4_1 _1175_ (.A(_0559_),
    .B(_0560_),
    .C(_0561_),
    .D(_0562_),
    .Y(_0563_));
 sky130_fd_sc_hd__nor4_1 _1176_ (.A(\mixed_output[13] ),
    .B(\mixed_output[14] ),
    .C(\mixed_output[15] ),
    .D(\mixed_output[23] ),
    .Y(_0564_));
 sky130_fd_sc_hd__nor4_1 _1177_ (.A(\mixed_output[0] ),
    .B(\mixed_output[10] ),
    .C(\mixed_output[11] ),
    .D(\mixed_output[12] ),
    .Y(_0565_));
 sky130_fd_sc_hd__nor4_1 _1178_ (.A(\mixed_output[16] ),
    .B(\mixed_output[20] ),
    .C(\mixed_output[21] ),
    .D(\mixed_output[22] ),
    .Y(_0566_));
 sky130_fd_sc_hd__nor4_1 _1179_ (.A(\mixed_output[17] ),
    .B(\mixed_output[18] ),
    .C(\mixed_output[19] ),
    .D(\mixed_output[1] ),
    .Y(_0567_));
 sky130_fd_sc_hd__nand4_1 _1180_ (.A(_0564_),
    .B(_0565_),
    .C(_0566_),
    .D(_0567_),
    .Y(_0568_));
 sky130_fd_sc_hd__o21ai_0 _1181_ (.A1(_0563_),
    .A2(_0568_),
    .B1(_0141_),
    .Y(_0569_));
 sky130_fd_sc_hd__a31o_1 _1182_ (.A1(net26),
    .A2(_0555_),
    .A3(_0558_),
    .B1(_0569_),
    .X(net36));
 sky130_fd_sc_hd__ha_1 _1183_ (.A(_0570_),
    .B(_0571_),
    .COUT(_0572_),
    .SUM(_0573_));
 sky130_fd_sc_hd__ha_1 _1184_ (.A(\health_counter[0] ),
    .B(\health_counter[1] ),
    .COUT(_0574_),
    .SUM(_0575_));
 sky130_fd_sc_hd__dfxtp_1 \data_valid_reg$_SDFF_PN0_  (.D(_0001_),
    .Q(net2),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[0]$_SDFFE_PN1P_  (.D(_0002_),
    .Q(\entropy_pool2[0] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[10]$_SDFFE_PN1P_  (.D(_0003_),
    .Q(\entropy_pool2[10] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[11]$_SDFFE_PN1P_  (.D(_0004_),
    .Q(\entropy_pool2[11] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[12]$_SDFFE_PN1P_  (.D(_0005_),
    .Q(\entropy_pool2[12] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[13]$_SDFFE_PN1P_  (.D(_0006_),
    .Q(\entropy_pool2[13] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[14]$_SDFFE_PN1P_  (.D(_0007_),
    .Q(\entropy_pool2[14] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[15]$_SDFFE_PN1P_  (.D(_0008_),
    .Q(\entropy_pool2[15] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[16]$_SDFFE_PN1P_  (.D(_0009_),
    .Q(\entropy_pool2[16] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[17]$_SDFFE_PN1P_  (.D(_0010_),
    .Q(\entropy_pool2[17] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[18]$_SDFFE_PN1P_  (.D(_0011_),
    .Q(\entropy_pool2[18] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[19]$_SDFFE_PN1P_  (.D(_0012_),
    .Q(\entropy_pool2[19] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[1]$_SDFFE_PN1P_  (.D(_0013_),
    .Q(\entropy_pool2[1] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[20]$_SDFFE_PN1P_  (.D(_0014_),
    .Q(\entropy_pool2[20] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[21]$_SDFFE_PN1P_  (.D(_0015_),
    .Q(\entropy_pool2[21] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[22]$_SDFFE_PN1P_  (.D(_0016_),
    .Q(\entropy_pool2[22] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[23]$_SDFFE_PN1P_  (.D(_0017_),
    .Q(\entropy_pool2[23] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[24]$_SDFFE_PN1P_  (.D(_0018_),
    .Q(\entropy_pool2[24] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[25]$_SDFFE_PN1P_  (.D(_0019_),
    .Q(\entropy_pool2[25] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[26]$_SDFFE_PN1P_  (.D(_0020_),
    .Q(\entropy_pool2[26] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[27]$_SDFFE_PN1P_  (.D(_0021_),
    .Q(\entropy_pool2[27] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[28]$_SDFFE_PN1P_  (.D(_0022_),
    .Q(\entropy_pool2[28] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[29]$_SDFFE_PN1P_  (.D(_0023_),
    .Q(\entropy_pool2[29] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[2]$_SDFFE_PN1P_  (.D(_0024_),
    .Q(\entropy_pool2[2] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[30]$_SDFFE_PN1P_  (.D(_0025_),
    .Q(\entropy_pool2[30] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[31]$_SDFFE_PN1P_  (.D(_0026_),
    .Q(\entropy_pool2[31] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[3]$_SDFFE_PN1P_  (.D(_0027_),
    .Q(\entropy_pool2[3] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[4]$_SDFFE_PN1P_  (.D(_0028_),
    .Q(\entropy_pool2[4] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[5]$_SDFFE_PN1P_  (.D(_0029_),
    .Q(\entropy_pool2[5] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[6]$_SDFFE_PN1P_  (.D(_0030_),
    .Q(\entropy_pool2[6] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[7]$_SDFFE_PN1P_  (.D(_0031_),
    .Q(\entropy_pool2[7] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[8]$_SDFFE_PN1P_  (.D(_0032_),
    .Q(\entropy_pool2[8] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool2[9]$_SDFFE_PN1P_  (.D(_0033_),
    .Q(\entropy_pool2[9] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[0]$_SDFFE_PN1P_  (.D(_0034_),
    .Q(\entropy_pool[0] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[10]$_SDFFE_PN0P_  (.D(_0035_),
    .Q(\entropy_pool[10] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[11]$_SDFFE_PN0P_  (.D(_0036_),
    .Q(\entropy_pool[11] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[12]$_SDFFE_PN0P_  (.D(_0037_),
    .Q(\entropy_pool[12] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[13]$_SDFFE_PN0P_  (.D(_0038_),
    .Q(\entropy_pool[13] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[14]$_SDFFE_PN0P_  (.D(_0039_),
    .Q(\entropy_pool[14] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[15]$_SDFFE_PN0P_  (.D(_0040_),
    .Q(\entropy_pool[15] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[16]$_SDFFE_PN0P_  (.D(_0041_),
    .Q(\entropy_pool[16] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[17]$_SDFFE_PN0P_  (.D(_0042_),
    .Q(\entropy_pool[17] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[18]$_SDFFE_PN0P_  (.D(_0043_),
    .Q(\entropy_pool[18] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[19]$_SDFFE_PN0P_  (.D(_0044_),
    .Q(\entropy_pool[19] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[1]$_SDFFE_PN0P_  (.D(_0045_),
    .Q(\entropy_pool[1] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[20]$_SDFFE_PN0P_  (.D(_0046_),
    .Q(\entropy_pool[20] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[21]$_SDFFE_PN0P_  (.D(_0047_),
    .Q(\entropy_pool[21] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[22]$_SDFFE_PN0P_  (.D(_0048_),
    .Q(\entropy_pool[22] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[23]$_SDFFE_PN0P_  (.D(_0049_),
    .Q(\entropy_pool[23] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[24]$_SDFFE_PN0P_  (.D(_0050_),
    .Q(\entropy_pool[24] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[25]$_SDFFE_PN0P_  (.D(_0051_),
    .Q(\entropy_pool[25] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[26]$_SDFFE_PN0P_  (.D(_0052_),
    .Q(\entropy_pool[26] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[27]$_SDFFE_PN0P_  (.D(_0053_),
    .Q(\entropy_pool[27] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[28]$_SDFFE_PN0P_  (.D(_0054_),
    .Q(\entropy_pool[28] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[29]$_SDFFE_PN0P_  (.D(_0055_),
    .Q(\entropy_pool[29] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[2]$_SDFFE_PN0P_  (.D(_0056_),
    .Q(\entropy_pool[2] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[30]$_SDFFE_PN0P_  (.D(_0057_),
    .Q(\entropy_pool[30] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[31]$_SDFFE_PN0P_  (.D(_0058_),
    .Q(\entropy_pool[31] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[3]$_SDFFE_PN0P_  (.D(_0059_),
    .Q(\entropy_pool[3] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[4]$_SDFFE_PN0P_  (.D(_0060_),
    .Q(\entropy_pool[4] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[5]$_SDFFE_PN0P_  (.D(_0061_),
    .Q(\entropy_pool[5] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[6]$_SDFFE_PN0P_  (.D(_0062_),
    .Q(\entropy_pool[6] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[7]$_SDFFE_PN0P_  (.D(_0063_),
    .Q(\entropy_pool[7] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[8]$_SDFFE_PN0P_  (.D(_0064_),
    .Q(\entropy_pool[8] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \entropy_pool[9]$_SDFFE_PN0P_  (.D(_0065_),
    .Q(\entropy_pool[9] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \gen_ring_osc.init_osc$_DFF_P_  (.D(_0000_),
    .Q(\gen_ring_osc.init_osc ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \gen_ring_osc.toggle_sampling$_SDFFE_PN0P_  (.D(_0066_),
    .Q(\gen_ring_osc.toggle_sampling ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \health_counter[0]$_SDFFE_PN0P_  (.D(_0067_),
    .Q(\health_counter[0] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \health_counter[1]$_SDFFE_PN0P_  (.D(_0068_),
    .Q(\health_counter[1] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \health_counter[2]$_SDFFE_PN0P_  (.D(_0069_),
    .Q(\health_counter[2] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \health_counter[3]$_SDFFE_PN0P_  (.D(_0070_),
    .Q(\health_counter[3] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \health_counter[4]$_SDFFE_PN0P_  (.D(_0071_),
    .Q(\health_counter[4] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \health_counter[5]$_SDFFE_PN0P_  (.D(_0072_),
    .Q(\health_counter[5] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \health_counter[6]$_SDFFE_PN0P_  (.D(_0073_),
    .Q(\health_counter[6] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \health_counter[7]$_SDFFE_PN0P_  (.D(_0074_),
    .Q(\health_counter[7] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \lfsr_reg[0]$_SDFFE_PN1P_  (.D(_0075_),
    .Q(\lfsr_reg[0] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \lfsr_reg[10]$_SDFFE_PN0P_  (.D(_0076_),
    .Q(\lfsr_reg[10] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \lfsr_reg[11]$_SDFFE_PN1P_  (.D(_0077_),
    .Q(\lfsr_reg[11] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfxtp_2 \lfsr_reg[12]$_SDFFE_PN0P_  (.D(_0078_),
    .Q(\lfsr_reg[12] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \lfsr_reg[13]$_SDFFE_PN1P_  (.D(_0079_),
    .Q(\lfsr_reg[13] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \lfsr_reg[14]$_SDFFE_PN1P_  (.D(_0080_),
    .Q(\lfsr_reg[14] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \lfsr_reg[15]$_SDFFE_PN1P_  (.D(_0081_),
    .Q(\lfsr_reg[15] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \lfsr_reg[16]$_SDFFE_PN1P_  (.D(_0082_),
    .Q(\lfsr_reg[16] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \lfsr_reg[17]$_SDFFE_PN0P_  (.D(_0083_),
    .Q(\lfsr_reg[17] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \lfsr_reg[18]$_SDFFE_PN1P_  (.D(_0084_),
    .Q(\lfsr_reg[18] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \lfsr_reg[19]$_SDFFE_PN1P_  (.D(_0085_),
    .Q(\lfsr_reg[19] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \lfsr_reg[1]$_SDFFE_PN0P_  (.D(_0086_),
    .Q(\lfsr_reg[1] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \lfsr_reg[20]$_SDFFE_PN0P_  (.D(_0087_),
    .Q(\lfsr_reg[20] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \lfsr_reg[21]$_SDFFE_PN0P_  (.D(_0088_),
    .Q(\lfsr_reg[21] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \lfsr_reg[22]$_SDFFE_PN1P_  (.D(_0089_),
    .Q(\lfsr_reg[22] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \lfsr_reg[23]$_SDFFE_PN1P_  (.D(_0090_),
    .Q(\lfsr_reg[23] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \lfsr_reg[24]$_SDFFE_PN1P_  (.D(_0091_),
    .Q(\lfsr_reg[24] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \lfsr_reg[25]$_SDFFE_PN1P_  (.D(_0092_),
    .Q(\lfsr_reg[25] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \lfsr_reg[26]$_SDFFE_PN0P_  (.D(_0093_),
    .Q(\lfsr_reg[26] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \lfsr_reg[27]$_SDFFE_PN1P_  (.D(_0094_),
    .Q(\lfsr_reg[27] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfxtp_2 \lfsr_reg[28]$_SDFFE_PN0P_  (.D(_0095_),
    .Q(\lfsr_reg[28] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfxtp_2 \lfsr_reg[29]$_SDFFE_PN1P_  (.D(_0096_),
    .Q(\lfsr_reg[29] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \lfsr_reg[2]$_SDFFE_PN0P_  (.D(_0097_),
    .Q(\lfsr_reg[2] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfxtp_2 \lfsr_reg[30]$_SDFFE_PN0P_  (.D(_0098_),
    .Q(\lfsr_reg[30] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \lfsr_reg[31]$_SDFFE_PN1P_  (.D(_0099_),
    .Q(\lfsr_reg[31] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfxtp_2 \lfsr_reg[3]$_SDFFE_PN0P_  (.D(_0100_),
    .Q(\lfsr_reg[3] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfxtp_2 \lfsr_reg[4]$_SDFFE_PN1P_  (.D(_0101_),
    .Q(\lfsr_reg[4] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \lfsr_reg[5]$_SDFFE_PN1P_  (.D(_0102_),
    .Q(\lfsr_reg[5] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \lfsr_reg[6]$_SDFFE_PN1P_  (.D(_0103_),
    .Q(\lfsr_reg[6] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \lfsr_reg[7]$_SDFFE_PN0P_  (.D(_0104_),
    .Q(\lfsr_reg[7] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \lfsr_reg[8]$_SDFFE_PN1P_  (.D(_0105_),
    .Q(\lfsr_reg[8] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \lfsr_reg[9]$_SDFFE_PN0P_  (.D(_0106_),
    .Q(\lfsr_reg[9] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[0]$_SDFFE_PN0N_  (.D(_0107_),
    .Q(\mixed_output[0] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[10]$_SDFFE_PN0N_  (.D(_0108_),
    .Q(\mixed_output[10] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[11]$_SDFFE_PN0N_  (.D(_0109_),
    .Q(\mixed_output[11] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[12]$_SDFFE_PN0N_  (.D(_0110_),
    .Q(\mixed_output[12] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[13]$_SDFFE_PN0N_  (.D(_0111_),
    .Q(\mixed_output[13] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[14]$_SDFFE_PN0N_  (.D(_0112_),
    .Q(\mixed_output[14] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[15]$_SDFFE_PN0N_  (.D(_0113_),
    .Q(\mixed_output[15] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[16]$_SDFFE_PN0N_  (.D(_0114_),
    .Q(\mixed_output[16] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[17]$_SDFFE_PN0N_  (.D(_0115_),
    .Q(\mixed_output[17] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[18]$_SDFFE_PN0N_  (.D(_0116_),
    .Q(\mixed_output[18] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[19]$_SDFFE_PN0N_  (.D(_0117_),
    .Q(\mixed_output[19] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[1]$_SDFFE_PN0N_  (.D(_0118_),
    .Q(\mixed_output[1] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[20]$_SDFFE_PN0N_  (.D(_0119_),
    .Q(\mixed_output[20] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[21]$_SDFFE_PN0N_  (.D(_0120_),
    .Q(\mixed_output[21] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[22]$_SDFFE_PN0N_  (.D(_0121_),
    .Q(\mixed_output[22] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[23]$_SDFFE_PN0N_  (.D(_0122_),
    .Q(\mixed_output[23] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[24]$_SDFFE_PN0N_  (.D(_0123_),
    .Q(\mixed_output[24] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[25]$_SDFFE_PN0N_  (.D(_0124_),
    .Q(\mixed_output[25] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[26]$_SDFFE_PN0N_  (.D(_0125_),
    .Q(\mixed_output[26] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[27]$_SDFFE_PN0N_  (.D(_0126_),
    .Q(\mixed_output[27] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[28]$_SDFFE_PN0N_  (.D(_0127_),
    .Q(\mixed_output[28] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[29]$_SDFFE_PN0N_  (.D(_0128_),
    .Q(\mixed_output[29] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[2]$_SDFFE_PN0N_  (.D(_0129_),
    .Q(\mixed_output[2] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[30]$_SDFFE_PN0N_  (.D(_0130_),
    .Q(\mixed_output[30] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[31]$_SDFFE_PN0N_  (.D(_0131_),
    .Q(\mixed_output[31] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[3]$_SDFFE_PN0N_  (.D(_0132_),
    .Q(\mixed_output[3] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[4]$_SDFFE_PN0N_  (.D(_0133_),
    .Q(\mixed_output[4] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[5]$_SDFFE_PN0N_  (.D(_0134_),
    .Q(\mixed_output[5] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[6]$_SDFFE_PN0N_  (.D(_0135_),
    .Q(\mixed_output[6] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[7]$_SDFFE_PN0N_  (.D(_0136_),
    .Q(\mixed_output[7] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[8]$_SDFFE_PN0N_  (.D(_0137_),
    .Q(\mixed_output[8] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \mixed_output[9]$_SDFFE_PN0N_  (.D(_0138_),
    .Q(\mixed_output[9] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfxtp_2 \state[0]$_SDFF_PN0_  (.D(_0139_),
    .Q(\state[0] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfxtp_2 \state[1]$_SDFF_PN0_  (.D(_0140_),
    .Q(\state[1] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_139 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(read_next),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 output2 (.A(net2),
    .X(data_valid));
 sky130_fd_sc_hd__clkbuf_1 output3 (.A(net3),
    .X(entropy_low));
 sky130_fd_sc_hd__clkbuf_1 output4 (.A(net4),
    .X(random_data[0]));
 sky130_fd_sc_hd__clkbuf_1 output5 (.A(net5),
    .X(random_data[10]));
 sky130_fd_sc_hd__clkbuf_1 output6 (.A(net6),
    .X(random_data[11]));
 sky130_fd_sc_hd__clkbuf_1 output7 (.A(net7),
    .X(random_data[12]));
 sky130_fd_sc_hd__clkbuf_1 output8 (.A(net8),
    .X(random_data[13]));
 sky130_fd_sc_hd__clkbuf_1 output9 (.A(net9),
    .X(random_data[14]));
 sky130_fd_sc_hd__clkbuf_1 output10 (.A(net10),
    .X(random_data[15]));
 sky130_fd_sc_hd__clkbuf_1 output11 (.A(net11),
    .X(random_data[16]));
 sky130_fd_sc_hd__clkbuf_1 output12 (.A(net12),
    .X(random_data[17]));
 sky130_fd_sc_hd__clkbuf_1 output13 (.A(net13),
    .X(random_data[18]));
 sky130_fd_sc_hd__clkbuf_1 output14 (.A(net14),
    .X(random_data[19]));
 sky130_fd_sc_hd__clkbuf_1 output15 (.A(net15),
    .X(random_data[1]));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net16),
    .X(random_data[20]));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net17),
    .X(random_data[21]));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net18),
    .X(random_data[22]));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net19),
    .X(random_data[23]));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net20),
    .X(random_data[24]));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net21),
    .X(random_data[25]));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net22),
    .X(random_data[26]));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net23),
    .X(random_data[27]));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net24),
    .X(random_data[28]));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net25),
    .X(random_data[29]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net26),
    .X(random_data[2]));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net27),
    .X(random_data[30]));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net28),
    .X(random_data[31]));
 sky130_fd_sc_hd__clkbuf_1 output29 (.A(net29),
    .X(random_data[3]));
 sky130_fd_sc_hd__clkbuf_1 output30 (.A(net30),
    .X(random_data[4]));
 sky130_fd_sc_hd__clkbuf_1 output31 (.A(net31),
    .X(random_data[5]));
 sky130_fd_sc_hd__clkbuf_1 output32 (.A(net32),
    .X(random_data[6]));
 sky130_fd_sc_hd__clkbuf_1 output33 (.A(net33),
    .X(random_data[7]));
 sky130_fd_sc_hd__clkbuf_1 output34 (.A(net34),
    .X(random_data[8]));
 sky130_fd_sc_hd__clkbuf_1 output35 (.A(net35),
    .X(random_data[9]));
 sky130_fd_sc_hd__clkbuf_1 output36 (.A(net36),
    .X(test_failed));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload0 (.A(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload1 (.A(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload2 (.A(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload3 (.A(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload4 (.A(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload5 (.A(clknet_4_8_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload6 (.A(clknet_4_9_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload7 (.A(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload8 (.A(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload9 (.A(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload10 (.A(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload11 (.A(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload12 (.A(clknet_4_15_0_clk));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_124 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_74 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_230 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_117 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_230 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_230 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_87 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_230 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_174 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_143 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_230 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_53 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_122 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_162 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_23 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_62 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_192 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_230 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_25 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_36 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_21 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_227 ();
endmodule
