module cordic_core (x_in,
    x_out,
    y_in,
    y_out,
    z_in);
 input [15:0] x_in;
 output [15:0] x_out;
 input [15:0] y_in;
 output [15:0] y_out;
 input [15:0] z_in;

 wire _0000_;
 wire net10;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire net4;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire net9;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire net17;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire net3;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire _4277_;
 wire _4278_;
 wire _4279_;
 wire _4280_;
 wire _4281_;
 wire _4282_;
 wire _4283_;
 wire _4284_;
 wire _4285_;
 wire _4286_;
 wire _4287_;
 wire _4288_;
 wire _4289_;
 wire _4290_;
 wire _4291_;
 wire _4292_;
 wire _4293_;
 wire _4294_;
 wire _4295_;
 wire _4296_;
 wire _4297_;
 wire _4298_;
 wire _4299_;
 wire _4300_;
 wire _4301_;
 wire _4302_;
 wire _4303_;
 wire _4304_;
 wire _4305_;
 wire _4306_;
 wire _4307_;
 wire _4308_;
 wire _4309_;
 wire _4310_;
 wire _4311_;
 wire _4312_;
 wire _4313_;
 wire _4314_;
 wire _4315_;
 wire _4316_;
 wire _4317_;
 wire _4318_;
 wire _4319_;
 wire _4320_;
 wire _4321_;
 wire _4322_;
 wire _4323_;
 wire _4324_;
 wire _4325_;
 wire _4326_;
 wire _4327_;
 wire _4328_;
 wire _4329_;
 wire _4330_;
 wire _4331_;
 wire _4332_;
 wire _4333_;
 wire _4334_;
 wire _4335_;
 wire _4336_;
 wire _4337_;
 wire _4338_;
 wire _4339_;
 wire _4340_;
 wire _4341_;
 wire _4342_;
 wire _4343_;
 wire _4344_;
 wire _4345_;
 wire _4346_;
 wire _4347_;
 wire _4348_;
 wire _4349_;
 wire _4350_;
 wire _4351_;
 wire _4352_;
 wire _4353_;
 wire _4354_;
 wire _4355_;
 wire _4356_;
 wire _4357_;
 wire _4358_;
 wire _4359_;
 wire _4360_;
 wire _4361_;
 wire _4362_;
 wire _4363_;
 wire _4364_;
 wire _4365_;
 wire _4366_;
 wire _4367_;
 wire _4368_;
 wire _4369_;
 wire _4370_;
 wire _4371_;
 wire _4372_;
 wire _4373_;
 wire _4374_;
 wire _4375_;
 wire _4376_;
 wire _4377_;
 wire _4378_;
 wire _4379_;
 wire _4380_;
 wire _4381_;
 wire _4382_;
 wire _4383_;
 wire _4384_;
 wire _4385_;
 wire _4386_;
 wire _4387_;
 wire _4388_;
 wire _4389_;
 wire _4390_;
 wire _4391_;
 wire _4392_;
 wire _4393_;
 wire _4394_;
 wire _4395_;
 wire _4396_;
 wire _4397_;
 wire _4398_;
 wire _4399_;
 wire _4400_;
 wire _4401_;
 wire _4402_;
 wire _4403_;
 wire _4404_;
 wire _4405_;
 wire _4406_;
 wire _4407_;
 wire _4408_;
 wire _4409_;
 wire _4410_;
 wire _4411_;
 wire _4412_;
 wire _4413_;
 wire _4414_;
 wire _4415_;
 wire _4416_;
 wire _4417_;
 wire _4418_;
 wire _4419_;
 wire _4420_;
 wire _4421_;
 wire _4422_;
 wire _4423_;
 wire _4424_;
 wire _4425_;
 wire _4426_;
 wire _4427_;
 wire _4428_;
 wire _4429_;
 wire _4430_;
 wire _4431_;
 wire _4432_;
 wire _4433_;
 wire _4434_;
 wire _4435_;
 wire _4436_;
 wire _4437_;
 wire _4438_;
 wire _4439_;
 wire _4440_;
 wire _4441_;
 wire _4442_;
 wire _4443_;
 wire _4444_;
 wire _4445_;
 wire _4446_;
 wire _4447_;
 wire _4448_;
 wire _4449_;
 wire _4450_;
 wire _4451_;
 wire _4452_;
 wire _4453_;
 wire _4454_;
 wire _4455_;
 wire _4456_;
 wire _4457_;
 wire _4458_;
 wire _4459_;
 wire _4460_;
 wire _4461_;
 wire _4462_;
 wire _4463_;
 wire _4464_;
 wire _4465_;
 wire _4466_;
 wire _4467_;
 wire _4468_;
 wire _4469_;
 wire _4470_;
 wire _4471_;
 wire _4472_;
 wire _4473_;
 wire _4474_;
 wire _4475_;
 wire _4476_;
 wire _4477_;
 wire _4478_;
 wire _4479_;
 wire _4480_;
 wire _4481_;
 wire _4482_;
 wire _4483_;
 wire _4484_;
 wire _4485_;
 wire _4486_;
 wire _4487_;
 wire _4488_;
 wire _4489_;
 wire _4490_;
 wire _4491_;
 wire _4492_;
 wire _4493_;
 wire _4494_;
 wire _4495_;
 wire _4496_;
 wire _4497_;
 wire _4498_;
 wire _4499_;
 wire _4500_;
 wire _4501_;
 wire _4502_;
 wire _4503_;
 wire _4504_;
 wire _4505_;
 wire _4506_;
 wire _4507_;
 wire _4508_;
 wire _4509_;
 wire _4510_;
 wire _4511_;
 wire _4512_;
 wire _4513_;
 wire _4514_;
 wire _4515_;
 wire _4516_;
 wire _4517_;
 wire _4518_;
 wire _4519_;
 wire _4520_;
 wire _4521_;
 wire _4522_;
 wire _4523_;
 wire _4524_;
 wire _4525_;
 wire _4526_;
 wire _4527_;
 wire _4528_;
 wire _4529_;
 wire _4530_;
 wire _4531_;
 wire _4532_;
 wire _4533_;
 wire _4534_;
 wire _4535_;
 wire _4536_;
 wire _4537_;
 wire _4538_;
 wire _4539_;
 wire _4540_;
 wire _4541_;
 wire _4542_;
 wire _4543_;
 wire _4544_;
 wire _4545_;
 wire _4546_;
 wire _4547_;
 wire _4548_;
 wire _4549_;
 wire _4550_;
 wire _4551_;
 wire _4552_;
 wire _4553_;
 wire _4554_;
 wire _4555_;
 wire _4556_;
 wire _4557_;
 wire _4558_;
 wire _4559_;
 wire _4560_;
 wire _4561_;
 wire _4562_;
 wire _4563_;
 wire _4564_;
 wire net1;
 wire net2;
 wire net18;
 wire net34;
 wire net67;
 wire net68;
 wire net69;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net173;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net209;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net303;
 wire net153;
 wire net154;
 wire net155;
 wire net168;
 wire net172;
 wire net178;
 wire net180;
 wire net202;
 wire net203;
 wire net204;
 wire net284;
 wire net285;
 wire net297;
 wire net314;
 wire net315;
 wire net316;

 BUF_X8 _4565_ (.A(net47),
    .Z(_0000_));
 INV_X8 _4566_ (.A(_0000_),
    .ZN(_4502_));
 NAND2_X2 clone10 (.A1(_0511_),
    .A2(_0516_),
    .ZN(net10));
 INV_X4 _4568_ (.A(_4503_),
    .ZN(_0002_));
 INV_X2 _4569_ (.A(net46),
    .ZN(_4501_));
 CLKBUF_X2 _4570_ (.A(_4505_),
    .Z(_0003_));
 OAI211_X4 _4571_ (.A(_4501_),
    .B(_0002_),
    .C1(_0003_),
    .C2(_4502_),
    .ZN(_0004_));
 BUF_X32 _4572_ (.A(z_in[0]),
    .Z(_0005_));
 NOR3_X2 _4573_ (.A1(net49),
    .A2(net48),
    .A3(_0005_),
    .ZN(_0006_));
 BUF_X4 _4574_ (.A(z_in[3]),
    .Z(_0007_));
 NOR4_X4 _4575_ (.A1(net52),
    .A2(net51),
    .A3(net50),
    .A4(_0007_),
    .ZN(_0008_));
 NOR4_X4 _4576_ (.A1(net42),
    .A2(net44),
    .A3(net43),
    .A4(net45),
    .ZN(_0009_));
 NOR3_X4 _4577_ (.A1(net55),
    .A2(net54),
    .A3(net53),
    .ZN(_0010_));
 NAND4_X2 _4578_ (.A1(_0006_),
    .A2(_0008_),
    .A3(_0009_),
    .A4(_0010_),
    .ZN(_0011_));
 OAI22_X4 _4579_ (.A1(_4502_),
    .A2(_0002_),
    .B1(_0011_),
    .B2(_0004_),
    .ZN(_0012_));
 INV_X4 _4580_ (.A(_0012_),
    .ZN(_0013_));
 BUF_X8 _4581_ (.A(_0013_),
    .Z(_0014_));
 BUF_X8 _4582_ (.A(_0014_),
    .Z(_0015_));
 BUF_X8 _4583_ (.A(_0015_),
    .Z(_2909_));
 CLKBUF_X2 _4584_ (.A(_2903_),
    .Z(_0016_));
 BUF_X8 _4585_ (.A(_0012_),
    .Z(_0017_));
 BUF_X8 _4586_ (.A(_0017_),
    .Z(_0018_));
 BUF_X8 _4587_ (.A(_0018_),
    .Z(_0019_));
 BUF_X4 _4588_ (.A(_0019_),
    .Z(_0020_));
 BUF_X4 _4589_ (.A(_0020_),
    .Z(_0021_));
 MUX2_X2 _4590_ (.A(_2899_),
    .B(_0016_),
    .S(_0021_),
    .Z(_3025_));
 INV_X2 _4591_ (.A(_3025_),
    .ZN(_2914_));
 BUF_X4 _4592_ (.A(_3029_),
    .Z(_0022_));
 BUF_X4 _4593_ (.A(_0022_),
    .Z(_0023_));
 BUF_X2 _4594_ (.A(_3036_),
    .Z(_0024_));
 INV_X1 _4595_ (.A(_3020_),
    .ZN(_0025_));
 BUF_X4 _4596_ (.A(_3019_),
    .Z(_0026_));
 INV_X2 _4597_ (.A(_0026_),
    .ZN(_0027_));
 OAI21_X1 _4598_ (.A(_0025_),
    .B1(_2904_),
    .B2(_0027_),
    .ZN(_0028_));
 BUF_X4 _4599_ (.A(_3037_),
    .Z(_0029_));
 AOI21_X2 _4600_ (.A(_0024_),
    .B1(_0028_),
    .B2(net130),
    .ZN(_0030_));
 XNOR2_X2 _4601_ (.A(_0023_),
    .B(_0030_),
    .ZN(_0031_));
 NAND2_X1 _4602_ (.A1(_0021_),
    .A2(_0031_),
    .ZN(_0032_));
 NOR2_X1 _4603_ (.A1(_3037_),
    .A2(_0026_),
    .ZN(_0033_));
 INV_X4 _4604_ (.A(_0029_),
    .ZN(_0034_));
 AOI221_X2 _4605_ (.A(_3041_),
    .B1(_0033_),
    .B2(_3017_),
    .C1(_0034_),
    .C2(_3023_),
    .ZN(_0035_));
 XNOR2_X2 _4606_ (.A(_0023_),
    .B(_0035_),
    .ZN(_0036_));
 OAI21_X2 _4607_ (.A(_0032_),
    .B1(_0036_),
    .B2(_0021_),
    .ZN(_3090_));
 BUF_X2 _4608_ (.A(_2905_),
    .Z(_0037_));
 NAND2_X1 _4609_ (.A1(_0037_),
    .A2(_0020_),
    .ZN(_0038_));
 BUF_X4 clone4 (.A(_1590_),
    .Z(net4));
 OAI21_X1 _4611_ (.A(_0038_),
    .B1(_0020_),
    .B2(_2902_),
    .ZN(_0040_));
 XNOR2_X2 _4612_ (.A(_0034_),
    .B(_0040_),
    .ZN(_3049_));
 INV_X1 _4613_ (.A(_3049_),
    .ZN(_3094_));
 MUX2_X2 _4614_ (.A(_0016_),
    .B(_2906_),
    .S(_0021_),
    .Z(_2919_));
 INV_X1 _4615_ (.A(_2919_),
    .ZN(_2923_));
 INV_X1 _4616_ (.A(_0003_),
    .ZN(_0041_));
 AOI21_X4 _4617_ (.A(_4503_),
    .B1(_0041_),
    .B2(_0000_),
    .ZN(_0042_));
 AND2_X1 _4618_ (.A1(_0006_),
    .A2(_0008_),
    .ZN(_0043_));
 NAND2_X1 _4619_ (.A1(_0043_),
    .A2(_0010_),
    .ZN(_0044_));
 OR2_X1 _4620_ (.A1(net43),
    .A2(net42),
    .ZN(_0045_));
 OR2_X1 _4621_ (.A1(net44),
    .A2(_0045_),
    .ZN(_0046_));
 OAI21_X1 _4622_ (.A(_0042_),
    .B1(_0044_),
    .B2(_0046_),
    .ZN(_0047_));
 XNOR2_X2 _4623_ (.A(net45),
    .B(_0047_),
    .ZN(_2907_));
 INV_X1 _4624_ (.A(_2907_),
    .ZN(_3102_));
 BUF_X4 _4625_ (.A(net130),
    .Z(_0048_));
 BUF_X2 _4626_ (.A(_2898_),
    .Z(_0049_));
 INV_X1 _4627_ (.A(_0049_),
    .ZN(_0050_));
 MUX2_X1 _4628_ (.A(_0050_),
    .B(_2902_),
    .S(_0020_),
    .Z(_0051_));
 XNOR2_X2 _4629_ (.A(_0048_),
    .B(_0051_),
    .ZN(_3097_));
 INV_X1 _4630_ (.A(_3097_),
    .ZN(_3045_));
 BUF_X8 _4631_ (.A(_2910_),
    .Z(_0052_));
 INV_X16 _4632_ (.A(_0052_),
    .ZN(_0053_));
 MUX2_X1 _4633_ (.A(_3051_),
    .B(_3094_),
    .S(_0053_),
    .Z(_3052_));
 INV_X1 _4634_ (.A(_3052_),
    .ZN(_2913_));
 BUF_X2 _4635_ (.A(_3048_),
    .Z(_0054_));
 XNOR2_X2 _4636_ (.A(_0054_),
    .B(_2915_),
    .ZN(_3055_));
 INV_X1 _4637_ (.A(_3055_),
    .ZN(_3246_));
 CLKBUF_X3 _4638_ (.A(_3033_),
    .Z(_0055_));
 INV_X1 _4639_ (.A(_0055_),
    .ZN(_0056_));
 BUF_X8 clone9 (.A(_0517_),
    .Z(net9));
 CLKBUF_X3 _4641_ (.A(_3059_),
    .Z(_0058_));
 BUF_X2 _4642_ (.A(_3071_),
    .Z(_0059_));
 INV_X1 _4643_ (.A(_0059_),
    .ZN(_0060_));
 NAND3_X1 _4644_ (.A1(_0056_),
    .A2(_0058_),
    .A3(_0060_),
    .ZN(_0061_));
 INV_X1 _4645_ (.A(_3041_),
    .ZN(_0062_));
 OR2_X1 _4646_ (.A1(_3037_),
    .A2(_0026_),
    .ZN(_0063_));
 INV_X1 _4647_ (.A(_3017_),
    .ZN(_2901_));
 INV_X1 _4648_ (.A(_3023_),
    .ZN(_0064_));
 OAI221_X2 _4649_ (.A(_0062_),
    .B1(_0063_),
    .B2(_2901_),
    .C1(_0029_),
    .C2(_0064_),
    .ZN(_0065_));
 INV_X4 _4650_ (.A(_0023_),
    .ZN(_0066_));
 AOI21_X1 _4651_ (.A(_0061_),
    .B1(_0065_),
    .B2(_0066_),
    .ZN(_0067_));
 BUF_X2 _4652_ (.A(_3067_),
    .Z(_0068_));
 BUF_X4 _4653_ (.A(_0068_),
    .Z(_0069_));
 NOR4_X2 _4654_ (.A1(_0023_),
    .A2(_0069_),
    .A3(_0058_),
    .A4(_0035_),
    .ZN(_0070_));
 INV_X4 _4655_ (.A(net117),
    .ZN(_0071_));
 NAND2_X1 _4656_ (.A1(_0071_),
    .A2(_0059_),
    .ZN(_0072_));
 NAND3_X1 _4657_ (.A1(_0069_),
    .A2(_0058_),
    .A3(_0060_),
    .ZN(_0073_));
 INV_X4 _4658_ (.A(_0068_),
    .ZN(_0074_));
 NAND3_X1 _4659_ (.A1(_0055_),
    .A2(_0074_),
    .A3(_0071_),
    .ZN(_0075_));
 NAND3_X1 _4660_ (.A1(_0072_),
    .A2(_0073_),
    .A3(_0075_),
    .ZN(_0076_));
 NOR3_X2 _4661_ (.A1(_0067_),
    .A2(_0070_),
    .A3(_0076_),
    .ZN(_0077_));
 BUF_X2 _4662_ (.A(_3028_),
    .Z(_0078_));
 INV_X1 _4663_ (.A(_0078_),
    .ZN(_0079_));
 CLKBUF_X3 _4664_ (.A(_3066_),
    .Z(_0080_));
 NOR2_X1 _4665_ (.A1(_0071_),
    .A2(_0080_),
    .ZN(_0081_));
 OAI21_X2 _4666_ (.A(_0022_),
    .B1(_0024_),
    .B2(_0029_),
    .ZN(_0082_));
 OR2_X1 _4667_ (.A1(_3020_),
    .A2(_0024_),
    .ZN(_0083_));
 INV_X1 _4668_ (.A(_2904_),
    .ZN(_0084_));
 AOI21_X2 _4669_ (.A(_0083_),
    .B1(_0084_),
    .B2(_0026_),
    .ZN(_0085_));
 OAI211_X2 _4670_ (.A(_0079_),
    .B(_0081_),
    .C1(_0082_),
    .C2(_0085_),
    .ZN(_0086_));
 NOR3_X1 _4671_ (.A1(_0069_),
    .A2(_0071_),
    .A3(_0080_),
    .ZN(_0087_));
 AOI21_X2 _4672_ (.A(_0087_),
    .B1(_0080_),
    .B2(_0071_),
    .ZN(_0088_));
 NOR2_X1 _4673_ (.A1(_3020_),
    .A2(_0024_),
    .ZN(_0089_));
 OAI21_X2 _4674_ (.A(_0089_),
    .B1(_2904_),
    .B2(_0027_),
    .ZN(_0090_));
 INV_X1 _4675_ (.A(_0082_),
    .ZN(_0091_));
 AOI21_X2 _4676_ (.A(_0078_),
    .B1(_0090_),
    .B2(_0091_),
    .ZN(_0092_));
 NOR2_X2 _4677_ (.A1(_0074_),
    .A2(_0058_),
    .ZN(_0093_));
 INV_X1 _4678_ (.A(_0093_),
    .ZN(_0094_));
 OAI211_X4 _4679_ (.A(_0086_),
    .B(_0088_),
    .C1(_0092_),
    .C2(_0094_),
    .ZN(_0095_));
 MUX2_X1 _4680_ (.A(_0077_),
    .B(_0095_),
    .S(_0021_),
    .Z(_3082_));
 BUF_X2 _4681_ (.A(_3075_),
    .Z(_0096_));
 INV_X2 _4682_ (.A(_0096_),
    .ZN(_0097_));
 NOR2_X1 _4683_ (.A1(_0058_),
    .A2(_0097_),
    .ZN(_0098_));
 BUF_X2 _4684_ (.A(_3063_),
    .Z(_0099_));
 OR2_X1 _4685_ (.A1(_0099_),
    .A2(_0096_),
    .ZN(_0100_));
 AOI211_X2 _4686_ (.A(_0059_),
    .B(_0100_),
    .C1(_0055_),
    .C2(_0074_),
    .ZN(_0101_));
 NOR2_X1 _4687_ (.A1(_0023_),
    .A2(_0069_),
    .ZN(_0102_));
 NOR2_X1 _4688_ (.A1(_0029_),
    .A2(_2902_),
    .ZN(_0103_));
 OAI21_X2 _4689_ (.A(_0102_),
    .B1(_0103_),
    .B2(_3041_),
    .ZN(_0104_));
 MUX2_X1 _4690_ (.A(_0098_),
    .B(_0101_),
    .S(_0104_),
    .Z(_0105_));
 INV_X1 _4691_ (.A(_0099_),
    .ZN(_0106_));
 NAND3_X1 _4692_ (.A1(_0058_),
    .A2(_0106_),
    .A3(_0097_),
    .ZN(_0107_));
 CLKBUF_X3 _4693_ (.A(_0096_),
    .Z(_0108_));
 NAND2_X1 _4694_ (.A1(_0071_),
    .A2(_0108_),
    .ZN(_0109_));
 AOI21_X2 _4695_ (.A(_0059_),
    .B1(_0074_),
    .B2(_0055_),
    .ZN(_0110_));
 OAI221_X2 _4696_ (.A(_0107_),
    .B1(_0109_),
    .B2(_0110_),
    .C1(_0106_),
    .C2(_0097_),
    .ZN(_0111_));
 OR3_X1 _4697_ (.A1(_0014_),
    .A2(_0105_),
    .A3(_0111_),
    .ZN(_0112_));
 BUF_X2 _4698_ (.A(_3069_),
    .Z(_0113_));
 OR2_X1 _4699_ (.A1(_0113_),
    .A2(_3061_),
    .ZN(_0114_));
 BUF_X2 _4700_ (.A(_3039_),
    .Z(_0115_));
 BUF_X2 _4701_ (.A(_3031_),
    .Z(_0116_));
 NOR2_X1 _4702_ (.A1(_0115_),
    .A2(_0116_),
    .ZN(_0117_));
 OAI21_X2 _4703_ (.A(_0117_),
    .B1(_0049_),
    .B2(_0034_),
    .ZN(_0118_));
 INV_X1 _4704_ (.A(_0116_),
    .ZN(_0119_));
 AOI21_X2 _4705_ (.A(_0074_),
    .B1(_0119_),
    .B2(_0066_),
    .ZN(_0120_));
 AOI21_X1 _4706_ (.A(_0114_),
    .B1(_0118_),
    .B2(_0120_),
    .ZN(_0121_));
 NOR2_X2 _4707_ (.A1(_3059_),
    .A2(_3061_),
    .ZN(_0122_));
 OR2_X1 _4708_ (.A1(_0121_),
    .A2(_0122_),
    .ZN(_0123_));
 XNOR2_X1 _4709_ (.A(_0108_),
    .B(_0123_),
    .ZN(_0124_));
 OAI21_X2 _4710_ (.A(_0112_),
    .B1(_0124_),
    .B2(_0020_),
    .ZN(_0125_));
 INV_X1 _4711_ (.A(_0125_),
    .ZN(_3210_));
 NOR3_X1 _4712_ (.A1(_0071_),
    .A2(_0113_),
    .A3(_0116_),
    .ZN(_0126_));
 OAI21_X2 _4713_ (.A(_0023_),
    .B1(_0115_),
    .B2(net130),
    .ZN(_0127_));
 OR2_X1 _4714_ (.A1(_0115_),
    .A2(_3021_),
    .ZN(_0128_));
 INV_X1 _4715_ (.A(_2897_),
    .ZN(_0129_));
 AOI21_X4 _4716_ (.A(_0128_),
    .B1(_0129_),
    .B2(_0026_),
    .ZN(_0130_));
 OAI21_X1 _4717_ (.A(_0126_),
    .B1(_0127_),
    .B2(_0130_),
    .ZN(_0131_));
 NOR2_X1 _4718_ (.A1(_0115_),
    .A2(_3021_),
    .ZN(_0132_));
 OAI21_X2 _4719_ (.A(_0132_),
    .B1(_2897_),
    .B2(_0027_),
    .ZN(_0133_));
 INV_X1 _4720_ (.A(_0127_),
    .ZN(_0134_));
 NAND3_X1 _4721_ (.A1(_0093_),
    .A2(_0133_),
    .A3(_0134_),
    .ZN(_0135_));
 NOR3_X1 _4722_ (.A1(_0069_),
    .A2(_0071_),
    .A3(_0113_),
    .ZN(_0136_));
 AOI221_X2 _4723_ (.A(_0136_),
    .B1(_0093_),
    .B2(_0116_),
    .C1(_0071_),
    .C2(_0113_),
    .ZN(_0137_));
 NAND4_X1 _4724_ (.A1(_0014_),
    .A2(_0131_),
    .A3(_0135_),
    .A4(_0137_),
    .ZN(_0138_));
 OR3_X1 _4725_ (.A1(_0067_),
    .A2(_0070_),
    .A3(_0076_),
    .ZN(_0139_));
 NAND2_X1 _4726_ (.A1(_0020_),
    .A2(_0139_),
    .ZN(_0140_));
 AND2_X1 _4727_ (.A1(_0138_),
    .A2(_0140_),
    .ZN(_3214_));
 OR2_X1 _4728_ (.A1(_0115_),
    .A2(_0116_),
    .ZN(_0141_));
 AOI21_X2 _4729_ (.A(_0141_),
    .B1(_0050_),
    .B2(_0048_),
    .ZN(_0142_));
 OAI21_X1 _4730_ (.A(_0069_),
    .B1(_0116_),
    .B2(_0023_),
    .ZN(_0143_));
 NOR2_X1 _4731_ (.A1(_0142_),
    .A2(_0143_),
    .ZN(_0144_));
 NAND2_X1 _4732_ (.A1(_0074_),
    .A2(_0119_),
    .ZN(_0145_));
 INV_X1 _4733_ (.A(_0115_),
    .ZN(_0146_));
 OAI21_X1 _4734_ (.A(_0146_),
    .B1(_0049_),
    .B2(_0034_),
    .ZN(_0147_));
 AOI21_X1 _4735_ (.A(_0145_),
    .B1(_0147_),
    .B2(_0023_),
    .ZN(_0148_));
 OAI21_X1 _4736_ (.A(_2909_),
    .B1(_0144_),
    .B2(_0148_),
    .ZN(_0149_));
 OR2_X1 _4737_ (.A1(net130),
    .A2(_2902_),
    .ZN(_0150_));
 AOI21_X2 _4738_ (.A(_0023_),
    .B1(_0062_),
    .B2(_0150_),
    .ZN(_0151_));
 OAI21_X2 _4739_ (.A(_0069_),
    .B1(_0151_),
    .B2(_0055_),
    .ZN(_0152_));
 OR3_X2 _4740_ (.A1(_0055_),
    .A2(_0069_),
    .A3(_0151_),
    .ZN(_0153_));
 NAND3_X1 _4741_ (.A1(_0021_),
    .A2(_0152_),
    .A3(_0153_),
    .ZN(_0154_));
 AND2_X1 _4742_ (.A1(_0149_),
    .A2(_0154_),
    .ZN(_3218_));
 NOR2_X2 _4743_ (.A1(_0130_),
    .A2(_0127_),
    .ZN(_0155_));
 INV_X1 _4744_ (.A(_3021_),
    .ZN(_0156_));
 OAI21_X1 _4745_ (.A(_0156_),
    .B1(_2897_),
    .B2(_0027_),
    .ZN(_0157_));
 AOI211_X2 _4746_ (.A(_0023_),
    .B(_0115_),
    .C1(_0157_),
    .C2(_0048_),
    .ZN(_0158_));
 OAI21_X1 _4747_ (.A(_2909_),
    .B1(_0155_),
    .B2(_0158_),
    .ZN(_0159_));
 NAND2_X1 _4748_ (.A1(_0021_),
    .A2(_0036_),
    .ZN(_0160_));
 AND2_X1 _4749_ (.A1(_0159_),
    .A2(_0160_),
    .ZN(_3135_));
 BUF_X32 _4750_ (.A(_0053_),
    .Z(_2929_));
 XNOR2_X1 _4751_ (.A(_0048_),
    .B(_0049_),
    .ZN(_0161_));
 OR2_X1 _4752_ (.A1(_2899_),
    .A2(_0161_),
    .ZN(_0162_));
 OAI22_X1 _4753_ (.A1(_0144_),
    .A2(_0148_),
    .B1(_0158_),
    .B2(_0155_),
    .ZN(_0163_));
 NAND2_X1 _4754_ (.A1(_0048_),
    .A2(_2902_),
    .ZN(_0164_));
 AOI21_X1 _4755_ (.A(_0016_),
    .B1(_0150_),
    .B2(_0164_),
    .ZN(_0165_));
 NAND4_X1 _4756_ (.A1(_0036_),
    .A2(_0152_),
    .A3(_0153_),
    .A4(_0165_),
    .ZN(_0166_));
 OAI33_X1 _4757_ (.A1(_0138_),
    .A2(_0162_),
    .A3(_0163_),
    .B1(_0166_),
    .B2(_0015_),
    .B3(_0077_),
    .ZN(_0167_));
 NOR2_X1 _4758_ (.A1(net227),
    .A2(_0167_),
    .ZN(_0168_));
 XOR2_X2 _4759_ (.A(_0125_),
    .B(_0168_),
    .Z(_3081_));
 NAND2_X1 _4760_ (.A1(_0152_),
    .A2(_0153_),
    .ZN(_0169_));
 INV_X1 _4761_ (.A(_0037_),
    .ZN(_0170_));
 AOI21_X1 _4762_ (.A(_0024_),
    .B1(_0170_),
    .B2(net130),
    .ZN(_0171_));
 OAI21_X1 _4763_ (.A(_0079_),
    .B1(_0171_),
    .B2(_0066_),
    .ZN(_0172_));
 XNOR2_X1 _4764_ (.A(_0074_),
    .B(_0172_),
    .ZN(_0173_));
 MUX2_X1 _4765_ (.A(_0169_),
    .B(_0173_),
    .S(_0021_),
    .Z(_3086_));
 INV_X1 _4766_ (.A(_3098_),
    .ZN(_0174_));
 NAND3_X1 _4767_ (.A1(_0036_),
    .A2(_0152_),
    .A3(_0153_),
    .ZN(_0175_));
 MUX2_X1 _4768_ (.A(_0163_),
    .B(_0175_),
    .S(_0020_),
    .Z(_0176_));
 NOR2_X2 _4769_ (.A1(_0174_),
    .A2(_0176_),
    .ZN(_0177_));
 NOR2_X1 _4770_ (.A1(net227),
    .A2(_0177_),
    .ZN(_0178_));
 XNOR2_X1 _4771_ (.A(_3214_),
    .B(_0178_),
    .ZN(_3085_));
 BUF_X8 _4772_ (.A(_0052_),
    .Z(_0179_));
 OR2_X1 _4773_ (.A1(_2899_),
    .A2(_0020_),
    .ZN(_0180_));
 NOR2_X1 _4774_ (.A1(_0050_),
    .A2(_0180_),
    .ZN(_0181_));
 NOR2_X1 _4775_ (.A1(_0016_),
    .A2(_2902_),
    .ZN(_0182_));
 AOI21_X1 _4776_ (.A(_0181_),
    .B1(_0182_),
    .B2(_0020_),
    .ZN(_0183_));
 NOR2_X1 _4777_ (.A1(_0048_),
    .A2(_0183_),
    .ZN(_0184_));
 INV_X1 _4778_ (.A(_0016_),
    .ZN(_0185_));
 NAND2_X1 _4779_ (.A1(_0185_),
    .A2(_2902_),
    .ZN(_0186_));
 OAI22_X1 _4780_ (.A1(_0049_),
    .A2(_0180_),
    .B1(_0186_),
    .B2(_2909_),
    .ZN(_0187_));
 AOI21_X1 _4781_ (.A(_0184_),
    .B1(_0187_),
    .B2(_0048_),
    .ZN(_0188_));
 OAI21_X1 _4782_ (.A(_0179_),
    .B1(_3135_),
    .B2(_0188_),
    .ZN(_0189_));
 XOR2_X2 _4783_ (.A(_3218_),
    .B(_0189_),
    .Z(_3089_));
 NOR2_X1 _4784_ (.A1(_2929_),
    .A2(_3098_),
    .ZN(_0190_));
 XNOR2_X1 _4785_ (.A(_3135_),
    .B(_0190_),
    .ZN(_3093_));
 BUF_X4 _4786_ (.A(_0179_),
    .Z(_0191_));
 NOR2_X1 _4787_ (.A1(_0191_),
    .A2(_3097_),
    .ZN(_0192_));
 AOI21_X2 _4788_ (.A(_0192_),
    .B1(_3099_),
    .B2(_0191_),
    .ZN(_2918_));
 INV_X1 _4789_ (.A(_2922_),
    .ZN(_2917_));
 INV_X1 _4790_ (.A(_3100_),
    .ZN(_0193_));
 INV_X1 _4791_ (.A(_3101_),
    .ZN(_0194_));
 OAI21_X1 _4792_ (.A(_0193_),
    .B1(_2922_),
    .B2(_0194_),
    .ZN(_0195_));
 BUF_X1 _4793_ (.A(_3096_),
    .Z(_0196_));
 AOI21_X1 _4794_ (.A(_3095_),
    .B1(_0195_),
    .B2(_0196_),
    .ZN(_0197_));
 XNOR2_X2 _4795_ (.A(_0197_),
    .B(_3092_),
    .ZN(_3238_));
 INV_X1 _4796_ (.A(_3238_),
    .ZN(_3146_));
 XNOR2_X2 _4797_ (.A(_0196_),
    .B(_2920_),
    .ZN(_3145_));
 INV_X1 _4798_ (.A(_3145_),
    .ZN(_3242_));
 INV_X1 _4799_ (.A(_3091_),
    .ZN(_0198_));
 OR2_X1 _4800_ (.A1(_3095_),
    .A2(_3100_),
    .ZN(_0199_));
 AOI21_X1 _4801_ (.A(_0199_),
    .B1(_2917_),
    .B2(_3101_),
    .ZN(_0200_));
 OAI21_X1 _4802_ (.A(_3092_),
    .B1(_3095_),
    .B2(_0196_),
    .ZN(_0201_));
 OAI21_X1 _4803_ (.A(_0198_),
    .B1(_0200_),
    .B2(_0201_),
    .ZN(_0202_));
 BUF_X2 _4804_ (.A(_3088_),
    .Z(_0203_));
 AOI21_X2 _4805_ (.A(_3087_),
    .B1(_0202_),
    .B2(_0203_),
    .ZN(_0204_));
 XNOR2_X2 _4806_ (.A(_3084_),
    .B(_0204_),
    .ZN(_3230_));
 INV_X16 _4807_ (.A(_0005_),
    .ZN(_2940_));
 INV_X1 _4808_ (.A(net49),
    .ZN(_0205_));
 AOI211_X2 _4809_ (.A(_3290_),
    .B(_4503_),
    .C1(_0041_),
    .C2(_0000_),
    .ZN(_0206_));
 XNOR2_X2 _4810_ (.A(_0205_),
    .B(_0206_),
    .ZN(_2924_));
 INV_X1 _4811_ (.A(_2924_),
    .ZN(_2928_));
 XNOR2_X2 _4812_ (.A(_0052_),
    .B(_2911_),
    .ZN(_0207_));
 BUF_X1 _4813_ (.A(_3107_),
    .Z(_0208_));
 OAI21_X1 _4814_ (.A(_3104_),
    .B1(_0208_),
    .B2(_3106_),
    .ZN(_0209_));
 NOR2_X1 _4815_ (.A1(_0207_),
    .A2(_0209_),
    .ZN(_0210_));
 NOR2_X1 _4816_ (.A1(_3043_),
    .A2(_0210_),
    .ZN(_0211_));
 OR3_X2 _4817_ (.A1(_3043_),
    .A2(_3106_),
    .A3(_3109_),
    .ZN(_0212_));
 INV_X1 _4818_ (.A(_3110_),
    .ZN(_0213_));
 CLKBUF_X2 _4819_ (.A(_3113_),
    .Z(_0214_));
 NOR2_X1 _4820_ (.A1(_0214_),
    .A2(_3112_),
    .ZN(_0215_));
 NOR2_X1 _4821_ (.A1(_0213_),
    .A2(_0215_),
    .ZN(_0216_));
 INV_X1 _4822_ (.A(_3115_),
    .ZN(_0217_));
 BUF_X4 _4823_ (.A(_3122_),
    .Z(_0218_));
 AOI21_X4 _4824_ (.A(_3121_),
    .B1(_3124_),
    .B2(_0218_),
    .ZN(_0219_));
 INV_X4 _4825_ (.A(_0219_),
    .ZN(_0220_));
 BUF_X2 _4826_ (.A(_3119_),
    .Z(_0221_));
 AOI21_X4 _4827_ (.A(_3118_),
    .B1(_0220_),
    .B2(_0221_),
    .ZN(_0222_));
 INV_X1 _4828_ (.A(_3116_),
    .ZN(_0223_));
 OAI21_X4 _4829_ (.A(_0217_),
    .B1(_0222_),
    .B2(_0223_),
    .ZN(_0224_));
 NOR2_X4 _4830_ (.A1(_0224_),
    .A2(_3112_),
    .ZN(_0225_));
 NAND4_X1 _4831_ (.A1(_3116_),
    .A2(_0218_),
    .A3(_3125_),
    .A4(_0221_),
    .ZN(_0226_));
 BUF_X1 _4832_ (.A(_3131_),
    .Z(_0227_));
 AOI21_X1 _4833_ (.A(_3130_),
    .B1(_3132_),
    .B2(_0227_),
    .ZN(_0228_));
 NAND2_X1 _4834_ (.A1(_0227_),
    .A2(_3133_),
    .ZN(_0229_));
 OAI21_X2 _4835_ (.A(_0228_),
    .B1(_0229_),
    .B2(_2928_),
    .ZN(_0230_));
 AOI21_X2 _4836_ (.A(_3127_),
    .B1(_0230_),
    .B2(_3128_),
    .ZN(_0231_));
 OAI21_X4 _4837_ (.A(_0225_),
    .B1(_0226_),
    .B2(_0231_),
    .ZN(_0232_));
 AOI21_X4 _4838_ (.A(_0212_),
    .B1(_0232_),
    .B2(_0216_),
    .ZN(_0233_));
 NOR2_X4 _4839_ (.A1(_0233_),
    .A2(_0211_),
    .ZN(_0234_));
 INV_X8 _4840_ (.A(_0234_),
    .ZN(_0235_));
 BUF_X16 _4841_ (.A(_0235_),
    .Z(_3261_));
 BUF_X2 _4842_ (.A(_3137_),
    .Z(_0236_));
 INV_X1 _4843_ (.A(_0236_),
    .ZN(_0237_));
 INV_X1 _4844_ (.A(_3047_),
    .ZN(_0238_));
 AOI21_X2 _4845_ (.A(_3053_),
    .B1(_3149_),
    .B2(_3054_),
    .ZN(_0239_));
 INV_X1 _4846_ (.A(_0054_),
    .ZN(_0240_));
 OAI21_X1 _4847_ (.A(_0238_),
    .B1(_0239_),
    .B2(_0240_),
    .ZN(_0241_));
 XNOR2_X2 _4848_ (.A(_0237_),
    .B(_0241_),
    .ZN(_3138_));
 INV_X1 _4849_ (.A(_3138_),
    .ZN(_3245_));
 CLKBUF_X2 _4850_ (.A(_3141_),
    .Z(_0242_));
 INV_X1 _4851_ (.A(_3143_),
    .ZN(_0243_));
 AOI21_X1 _4852_ (.A(_3150_),
    .B1(_3151_),
    .B2(_2930_),
    .ZN(_0244_));
 INV_X1 _4853_ (.A(_3144_),
    .ZN(_0245_));
 OAI21_X2 _4854_ (.A(_0243_),
    .B1(_0244_),
    .B2(_0245_),
    .ZN(_0246_));
 XNOR2_X2 _4855_ (.A(_0242_),
    .B(_0246_),
    .ZN(_3464_));
 BUF_X2 _4856_ (.A(_3159_),
    .Z(_0247_));
 BUF_X4 _4857_ (.A(_0247_),
    .Z(_0248_));
 INV_X2 _4858_ (.A(_0248_),
    .ZN(_0249_));
 BUF_X2 _4859_ (.A(_3074_),
    .Z(_0250_));
 BUF_X2 _4860_ (.A(_3058_),
    .Z(_0251_));
 AOI21_X1 _4861_ (.A(_0250_),
    .B1(_0251_),
    .B2(_0096_),
    .ZN(_0252_));
 NAND2_X1 _4862_ (.A1(net117),
    .A2(_0096_),
    .ZN(_0253_));
 NOR2_X1 _4863_ (.A1(_0068_),
    .A2(_0080_),
    .ZN(_0254_));
 OAI21_X2 _4864_ (.A(_0252_),
    .B1(_0253_),
    .B2(_0254_),
    .ZN(_0255_));
 NOR4_X1 _4865_ (.A1(_0078_),
    .A2(_0080_),
    .A3(_0251_),
    .A4(_0250_),
    .ZN(_0256_));
 OAI21_X2 _4866_ (.A(_0256_),
    .B1(_0082_),
    .B2(_0085_),
    .ZN(_0257_));
 AOI21_X2 _4867_ (.A(_0249_),
    .B1(_0255_),
    .B2(_0257_),
    .ZN(_0258_));
 OR4_X1 _4868_ (.A1(_0078_),
    .A2(_0080_),
    .A3(_0251_),
    .A4(_0250_),
    .ZN(_0259_));
 AOI21_X4 _4869_ (.A(_0259_),
    .B1(_0091_),
    .B2(_0090_),
    .ZN(_0260_));
 NAND2_X1 _4870_ (.A1(_0249_),
    .A2(_0255_),
    .ZN(_0261_));
 OAI21_X2 _4871_ (.A(_0017_),
    .B1(_0260_),
    .B2(_0261_),
    .ZN(_0262_));
 BUF_X2 _4872_ (.A(_3079_),
    .Z(_0263_));
 INV_X1 _4873_ (.A(_0263_),
    .ZN(_0264_));
 NOR2_X1 _4874_ (.A1(_0022_),
    .A2(_3059_),
    .ZN(_0265_));
 OAI211_X2 _4875_ (.A(_0097_),
    .B(_0265_),
    .C1(_0059_),
    .C2(_0074_),
    .ZN(_0266_));
 OR2_X1 _4876_ (.A1(_0099_),
    .A2(_0059_),
    .ZN(_0267_));
 AOI21_X2 _4877_ (.A(_0267_),
    .B1(_0074_),
    .B2(_0055_),
    .ZN(_0268_));
 OAI21_X2 _4878_ (.A(_0097_),
    .B1(_0099_),
    .B2(_0071_),
    .ZN(_0269_));
 OAI221_X2 _4879_ (.A(_0264_),
    .B1(_0035_),
    .B2(_0266_),
    .C1(_0268_),
    .C2(_0269_),
    .ZN(_0270_));
 XNOR2_X2 _4880_ (.A(_0248_),
    .B(_0270_),
    .ZN(_0271_));
 OAI22_X1 _4881_ (.A1(_0258_),
    .A2(_0262_),
    .B1(_0271_),
    .B2(_0021_),
    .ZN(_0272_));
 INV_X1 _4882_ (.A(_0272_),
    .ZN(_3174_));
 BUF_X2 _4883_ (.A(_3167_),
    .Z(_0273_));
 INV_X2 _4884_ (.A(_0273_),
    .ZN(_0274_));
 CLKBUF_X3 _4885_ (.A(_3077_),
    .Z(_0275_));
 AOI21_X4 _4886_ (.A(_3161_),
    .B1(_0275_),
    .B2(_0247_),
    .ZN(_0276_));
 NAND2_X1 _4887_ (.A1(_0096_),
    .A2(_0248_),
    .ZN(_0277_));
 OAI21_X2 _4888_ (.A(_0276_),
    .B1(_0277_),
    .B2(_0122_),
    .ZN(_0278_));
 NOR2_X1 _4889_ (.A1(_0113_),
    .A2(_3061_),
    .ZN(_0279_));
 AND2_X1 _4890_ (.A1(_0279_),
    .A2(_0276_),
    .ZN(_0280_));
 OAI21_X2 _4891_ (.A(_0280_),
    .B1(_0143_),
    .B2(_0142_),
    .ZN(_0281_));
 AOI21_X1 _4892_ (.A(_0019_),
    .B1(_0278_),
    .B2(_0281_),
    .ZN(_0282_));
 BUF_X2 _4893_ (.A(_3163_),
    .Z(_0283_));
 NOR3_X4 _4894_ (.A1(_0099_),
    .A2(_0263_),
    .A3(_0283_),
    .ZN(_0284_));
 AND3_X2 _4895_ (.A1(_0104_),
    .A2(_0110_),
    .A3(_0284_),
    .ZN(_0285_));
 AOI21_X2 _4896_ (.A(_0096_),
    .B1(_0106_),
    .B2(net117),
    .ZN(_0286_));
 OAI21_X1 _4897_ (.A(_0249_),
    .B1(_0286_),
    .B2(_0263_),
    .ZN(_0287_));
 INV_X2 _4898_ (.A(_0283_),
    .ZN(_0288_));
 AOI21_X2 _4899_ (.A(_0285_),
    .B1(_0287_),
    .B2(_0288_),
    .ZN(_0289_));
 AOI21_X2 _4900_ (.A(_0282_),
    .B1(_0289_),
    .B2(_0019_),
    .ZN(_0290_));
 XNOR2_X2 _4901_ (.A(_0274_),
    .B(_0290_),
    .ZN(_3202_));
 INV_X1 _4902_ (.A(_0275_),
    .ZN(_0291_));
 NAND2_X1 _4903_ (.A1(_0119_),
    .A2(_0279_),
    .ZN(_0292_));
 AOI21_X4 _4904_ (.A(_0292_),
    .B1(_0134_),
    .B2(_0133_),
    .ZN(_0293_));
 INV_X1 _4905_ (.A(_3061_),
    .ZN(_0294_));
 OAI21_X1 _4906_ (.A(_3059_),
    .B1(_0113_),
    .B2(_0069_),
    .ZN(_0295_));
 NAND2_X2 _4907_ (.A1(_0294_),
    .A2(_0295_),
    .ZN(_0296_));
 NAND2_X1 _4908_ (.A1(_0108_),
    .A2(_0296_),
    .ZN(_0297_));
 OAI21_X1 _4909_ (.A(_0291_),
    .B1(_0293_),
    .B2(_0297_),
    .ZN(_0298_));
 XNOR2_X1 _4910_ (.A(_0249_),
    .B(_0298_),
    .ZN(_0299_));
 MUX2_X2 _4911_ (.A(_0271_),
    .B(_0299_),
    .S(_0015_),
    .Z(_3206_));
 NAND2_X1 _4912_ (.A1(_0108_),
    .A2(_0014_),
    .ZN(_0300_));
 INV_X1 _4913_ (.A(_0296_),
    .ZN(_0301_));
 OAI211_X2 _4914_ (.A(_0249_),
    .B(_0291_),
    .C1(_0293_),
    .C2(_0301_),
    .ZN(_0302_));
 NAND3_X1 _4915_ (.A1(_0119_),
    .A2(_0291_),
    .A3(_0279_),
    .ZN(_0303_));
 OAI221_X2 _4916_ (.A(_0248_),
    .B1(_0275_),
    .B2(_0296_),
    .C1(_0303_),
    .C2(_0155_),
    .ZN(_0304_));
 AOI211_X2 _4917_ (.A(_0123_),
    .B(_0300_),
    .C1(_0302_),
    .C2(_0304_),
    .ZN(_0305_));
 XNOR2_X1 _4918_ (.A(_0248_),
    .B(_0275_),
    .ZN(_0306_));
 OAI211_X2 _4919_ (.A(_0015_),
    .B(_0306_),
    .C1(_0122_),
    .C2(_0121_),
    .ZN(_0307_));
 OAI22_X2 _4920_ (.A1(_0112_),
    .A2(_0271_),
    .B1(_0307_),
    .B2(_0108_),
    .ZN(_0308_));
 OAI21_X2 _4921_ (.A(_0167_),
    .B1(_0305_),
    .B2(_0308_),
    .ZN(_0309_));
 NAND2_X1 _4922_ (.A1(_0179_),
    .A2(_0309_),
    .ZN(_0310_));
 XOR2_X1 _4923_ (.A(_3202_),
    .B(_0310_),
    .Z(_3173_));
 INV_X1 _4924_ (.A(_0080_),
    .ZN(_0311_));
 NOR2_X1 _4925_ (.A1(_0097_),
    .A2(_0251_),
    .ZN(_0312_));
 OAI21_X2 _4926_ (.A(_0069_),
    .B1(_0078_),
    .B2(_0022_),
    .ZN(_0313_));
 OR2_X1 _4927_ (.A1(_0024_),
    .A2(_0078_),
    .ZN(_0314_));
 AOI21_X2 _4928_ (.A(_0314_),
    .B1(_0170_),
    .B2(_0029_),
    .ZN(_0315_));
 OAI211_X2 _4929_ (.A(_0311_),
    .B(_0312_),
    .C1(_0313_),
    .C2(_0315_),
    .ZN(_0316_));
 MUX2_X1 _4930_ (.A(_0109_),
    .B(_0108_),
    .S(_0251_),
    .Z(_0317_));
 NOR2_X1 _4931_ (.A1(_0024_),
    .A2(_0078_),
    .ZN(_0318_));
 OAI21_X2 _4932_ (.A(_0318_),
    .B1(_0037_),
    .B2(_0034_),
    .ZN(_0319_));
 INV_X1 _4933_ (.A(_0313_),
    .ZN(_0320_));
 AOI21_X2 _4934_ (.A(_0080_),
    .B1(_0319_),
    .B2(_0320_),
    .ZN(_0321_));
 NAND2_X1 _4935_ (.A1(_0058_),
    .A2(_0097_),
    .ZN(_0322_));
 OAI211_X4 _4936_ (.A(_0316_),
    .B(_0317_),
    .C1(_0321_),
    .C2(_0322_),
    .ZN(_0323_));
 NOR2_X1 _4937_ (.A1(_2909_),
    .A2(_0323_),
    .ZN(_0324_));
 NOR2_X1 _4938_ (.A1(_0105_),
    .A2(_0111_),
    .ZN(_0325_));
 AOI21_X2 _4939_ (.A(_0324_),
    .B1(_0325_),
    .B2(_2909_),
    .ZN(_3178_));
 INV_X1 _4940_ (.A(_3214_),
    .ZN(_0326_));
 NAND3_X1 _4941_ (.A1(_0125_),
    .A2(_0326_),
    .A3(_0177_),
    .ZN(_0327_));
 NAND2_X1 _4942_ (.A1(_0179_),
    .A2(_0327_),
    .ZN(_0328_));
 XOR2_X2 _4943_ (.A(_3206_),
    .B(_0328_),
    .Z(_3177_));
 BUF_X2 _4944_ (.A(_3176_),
    .Z(_0329_));
 BUF_X2 _4945_ (.A(_3179_),
    .Z(_0330_));
 INV_X1 _4946_ (.A(_0330_),
    .ZN(_0331_));
 CLKBUF_X2 _4947_ (.A(_3083_),
    .Z(_0332_));
 NOR2_X1 _4948_ (.A1(_3087_),
    .A2(_3091_),
    .ZN(_0333_));
 OAI21_X1 _4949_ (.A(_0333_),
    .B1(_0201_),
    .B2(_0200_),
    .ZN(_0334_));
 OAI21_X1 _4950_ (.A(_3084_),
    .B1(_0203_),
    .B2(_3087_),
    .ZN(_0335_));
 INV_X1 _4951_ (.A(_0335_),
    .ZN(_0336_));
 AOI21_X1 _4952_ (.A(_0332_),
    .B1(_0334_),
    .B2(_0336_),
    .ZN(_0337_));
 INV_X1 _4953_ (.A(_3180_),
    .ZN(_0338_));
 OAI21_X1 _4954_ (.A(_0331_),
    .B1(_0337_),
    .B2(_0338_),
    .ZN(_0339_));
 XNOR2_X2 _4955_ (.A(_0339_),
    .B(_0329_),
    .ZN(_0340_));
 INV_X1 _4956_ (.A(_0340_),
    .ZN(_3222_));
 BUF_X2 _4957_ (.A(_3183_),
    .Z(_0341_));
 CLKBUF_X3 _4958_ (.A(_0341_),
    .Z(_0342_));
 CLKBUF_X3 _4959_ (.A(_3195_),
    .Z(_0343_));
 INV_X2 _4960_ (.A(_3191_),
    .ZN(_0344_));
 AOI21_X4 _4961_ (.A(_0343_),
    .B1(_0344_),
    .B2(_3171_),
    .ZN(_0345_));
 CLKBUF_X3 _4962_ (.A(_0273_),
    .Z(_0346_));
 CLKBUF_X3 _4963_ (.A(_3191_),
    .Z(_0347_));
 OR2_X1 _4964_ (.A1(_0346_),
    .A2(_0347_),
    .ZN(_0348_));
 AOI21_X2 _4965_ (.A(_0348_),
    .B1(_0288_),
    .B2(_0248_),
    .ZN(_0349_));
 NAND3_X2 _4966_ (.A1(_0108_),
    .A2(_0264_),
    .A3(_0288_),
    .ZN(_0350_));
 NAND2_X1 _4967_ (.A1(_0058_),
    .A2(_0284_),
    .ZN(_0351_));
 NAND3_X1 _4968_ (.A1(_0349_),
    .A2(_0350_),
    .A3(_0351_),
    .ZN(_0352_));
 OAI211_X2 _4969_ (.A(_0014_),
    .B(_0345_),
    .C1(_0352_),
    .C2(_0285_),
    .ZN(_0353_));
 AOI21_X2 _4970_ (.A(_3190_),
    .B1(_3166_),
    .B2(_0347_),
    .ZN(_0354_));
 INV_X1 _4971_ (.A(_0354_),
    .ZN(_0355_));
 AND2_X1 _4972_ (.A1(_0346_),
    .A2(_0347_),
    .ZN(_0356_));
 AOI21_X1 _4973_ (.A(_3158_),
    .B1(_0250_),
    .B2(_0248_),
    .ZN(_0357_));
 NOR2_X1 _4974_ (.A1(_0058_),
    .A2(_0251_),
    .ZN(_0358_));
 OAI21_X2 _4975_ (.A(_0357_),
    .B1(_0358_),
    .B2(_0277_),
    .ZN(_0359_));
 AND2_X1 _4976_ (.A1(_0356_),
    .A2(_0359_),
    .ZN(_0360_));
 NOR3_X1 _4977_ (.A1(_0080_),
    .A2(_0251_),
    .A3(_3158_),
    .ZN(_0361_));
 INV_X1 _4978_ (.A(_0250_),
    .ZN(_0362_));
 OAI221_X2 _4979_ (.A(_0361_),
    .B1(_0313_),
    .B2(_0315_),
    .C1(_0249_),
    .C2(_0362_),
    .ZN(_0363_));
 AOI21_X2 _4980_ (.A(_0355_),
    .B1(_0360_),
    .B2(_0363_),
    .ZN(_0364_));
 OAI211_X2 _4981_ (.A(_0342_),
    .B(_0353_),
    .C1(_0364_),
    .C2(_0014_),
    .ZN(_0365_));
 INV_X2 _4982_ (.A(_0341_),
    .ZN(_0366_));
 NAND2_X1 _4983_ (.A1(_0356_),
    .A2(_0359_),
    .ZN(_0367_));
 OR3_X1 _4984_ (.A1(_0080_),
    .A2(_0251_),
    .A3(_3158_),
    .ZN(_0368_));
 AOI221_X2 _4985_ (.A(_0368_),
    .B1(_0319_),
    .B2(_0320_),
    .C1(_0248_),
    .C2(_0250_),
    .ZN(_0369_));
 OAI211_X2 _4986_ (.A(_0018_),
    .B(_0354_),
    .C1(_0367_),
    .C2(_0369_),
    .ZN(_0370_));
 INV_X1 _4987_ (.A(_0343_),
    .ZN(_0371_));
 INV_X2 _4988_ (.A(_3171_),
    .ZN(_0372_));
 OAI21_X1 _4989_ (.A(_0371_),
    .B1(_0347_),
    .B2(_0372_),
    .ZN(_0373_));
 AND3_X1 _4990_ (.A1(_0349_),
    .A2(_0350_),
    .A3(_0351_),
    .ZN(_0374_));
 NAND3_X2 _4991_ (.A1(_0104_),
    .A2(_0110_),
    .A3(_0284_),
    .ZN(_0375_));
 AOI21_X1 _4992_ (.A(_0373_),
    .B1(_0374_),
    .B2(_0375_),
    .ZN(_0376_));
 OAI211_X2 _4993_ (.A(_0366_),
    .B(_0370_),
    .C1(_0376_),
    .C2(_0018_),
    .ZN(_0377_));
 AND2_X1 _4994_ (.A1(_0365_),
    .A2(_0377_),
    .ZN(_0378_));
 INV_X1 _4995_ (.A(_0378_),
    .ZN(_3388_));
 OAI21_X2 _4996_ (.A(_0372_),
    .B1(_0346_),
    .B2(_0288_),
    .ZN(_0379_));
 NOR2_X2 _4997_ (.A1(_0247_),
    .A2(_0273_),
    .ZN(_0380_));
 NOR2_X1 _4998_ (.A1(_0379_),
    .A2(_0380_),
    .ZN(_0381_));
 OAI211_X2 _4999_ (.A(_0264_),
    .B(_0372_),
    .C1(_0346_),
    .C2(_0288_),
    .ZN(_0382_));
 NOR2_X1 _5000_ (.A1(_0099_),
    .A2(_0059_),
    .ZN(_0383_));
 OAI21_X2 _5001_ (.A(_0383_),
    .B1(_0068_),
    .B2(_0056_),
    .ZN(_0384_));
 OR2_X1 _5002_ (.A1(_0022_),
    .A2(_3059_),
    .ZN(_0385_));
 AOI211_X2 _5003_ (.A(_0096_),
    .B(_0385_),
    .C1(_0060_),
    .C2(_0068_),
    .ZN(_0386_));
 AOI221_X2 _5004_ (.A(_0382_),
    .B1(_0286_),
    .B2(_0384_),
    .C1(_0065_),
    .C2(_0386_),
    .ZN(_0387_));
 NOR3_X1 _5005_ (.A1(_0387_),
    .A2(_0381_),
    .A3(_0017_),
    .ZN(_0388_));
 AOI21_X2 _5006_ (.A(_3166_),
    .B1(_3158_),
    .B2(_0346_),
    .ZN(_0389_));
 INV_X1 _5007_ (.A(_0389_),
    .ZN(_0390_));
 AND3_X1 _5008_ (.A1(_0248_),
    .A2(_0346_),
    .A3(_0255_),
    .ZN(_0391_));
 AOI211_X2 _5009_ (.A(_0013_),
    .B(_0390_),
    .C1(_0391_),
    .C2(_0257_),
    .ZN(_0392_));
 OR3_X1 _5010_ (.A1(_0347_),
    .A2(_0388_),
    .A3(_0392_),
    .ZN(_0393_));
 OAI21_X1 _5011_ (.A(_0347_),
    .B1(_0388_),
    .B2(_0392_),
    .ZN(_0394_));
 AND2_X1 _5012_ (.A1(_0393_),
    .A2(_0394_),
    .ZN(_0395_));
 INV_X1 _5013_ (.A(_0395_),
    .ZN(_3320_));
 NAND3_X1 _5014_ (.A1(_0018_),
    .A2(_0363_),
    .A3(_0359_),
    .ZN(_0396_));
 OAI21_X1 _5015_ (.A(_0396_),
    .B1(_0289_),
    .B2(_0018_),
    .ZN(_0397_));
 XNOR2_X2 _5016_ (.A(_0274_),
    .B(_0397_),
    .ZN(_3324_));
 NOR3_X1 _5017_ (.A1(_0014_),
    .A2(_0381_),
    .A3(_0387_),
    .ZN(_0398_));
 NOR2_X1 _5018_ (.A1(_0116_),
    .A2(_0114_),
    .ZN(_0399_));
 OAI21_X2 _5019_ (.A(_0399_),
    .B1(_0127_),
    .B2(_0130_),
    .ZN(_0400_));
 AND4_X1 _5020_ (.A1(_0108_),
    .A2(_0248_),
    .A3(_0346_),
    .A4(_0296_),
    .ZN(_0401_));
 INV_X1 _5021_ (.A(_0276_),
    .ZN(_0402_));
 AOI221_X2 _5022_ (.A(_3169_),
    .B1(_0400_),
    .B2(_0401_),
    .C1(_0402_),
    .C2(_0346_),
    .ZN(_0403_));
 AOI21_X2 _5023_ (.A(_0398_),
    .B1(_0403_),
    .B2(_0014_),
    .ZN(_0404_));
 XNOR2_X2 _5024_ (.A(_0344_),
    .B(_0404_),
    .ZN(_3197_));
 INV_X1 _5025_ (.A(_3200_),
    .ZN(_0405_));
 BUF_X2 _5026_ (.A(_3204_),
    .Z(_0406_));
 AOI21_X2 _5027_ (.A(_3203_),
    .B1(_3207_),
    .B2(_0406_),
    .ZN(_0407_));
 AOI21_X2 _5028_ (.A(_3136_),
    .B1(_3047_),
    .B2(_0236_),
    .ZN(_0408_));
 NOR3_X1 _5029_ (.A1(_3211_),
    .A2(_3215_),
    .A3(_3219_),
    .ZN(_0409_));
 NAND2_X1 _5030_ (.A1(_0054_),
    .A2(_0236_),
    .ZN(_0410_));
 OAI211_X2 _5031_ (.A(_0408_),
    .B(_0409_),
    .C1(_0239_),
    .C2(_0410_),
    .ZN(_0411_));
 NOR2_X2 _5032_ (.A1(_3212_),
    .A2(_3211_),
    .ZN(_0412_));
 NOR2_X2 _5033_ (.A1(_3211_),
    .A2(_3215_),
    .ZN(_0413_));
 BUF_X2 _5034_ (.A(_3216_),
    .Z(_0414_));
 BUF_X4 _5035_ (.A(_3220_),
    .Z(_0415_));
 OAI21_X2 _5036_ (.A(_0414_),
    .B1(_0415_),
    .B2(_3219_),
    .ZN(_0416_));
 AOI21_X2 _5037_ (.A(_0412_),
    .B1(_0413_),
    .B2(_0416_),
    .ZN(_0417_));
 NAND2_X2 _5038_ (.A1(_0411_),
    .A2(_0417_),
    .ZN(_0418_));
 BUF_X2 _5039_ (.A(_3208_),
    .Z(_0419_));
 NAND2_X1 _5040_ (.A1(_0406_),
    .A2(_0419_),
    .ZN(_0420_));
 OAI21_X1 _5041_ (.A(_0407_),
    .B1(_0418_),
    .B2(_0420_),
    .ZN(_0421_));
 XNOR2_X2 _5042_ (.A(_0405_),
    .B(_0421_),
    .ZN(_3412_));
 INV_X1 _5043_ (.A(_2915_),
    .ZN(_0422_));
 AOI21_X2 _5044_ (.A(_3047_),
    .B1(_0422_),
    .B2(_0054_),
    .ZN(_0423_));
 NAND3_X2 _5045_ (.A1(_0236_),
    .A2(_0414_),
    .A3(_0415_),
    .ZN(_0424_));
 AOI21_X2 _5046_ (.A(_3219_),
    .B1(_3136_),
    .B2(_0415_),
    .ZN(_0425_));
 INV_X1 _5047_ (.A(_0414_),
    .ZN(_0426_));
 OAI221_X2 _5048_ (.A(_0413_),
    .B1(_0423_),
    .B2(_0424_),
    .C1(_0425_),
    .C2(_0426_),
    .ZN(_0427_));
 INV_X1 _5049_ (.A(_0419_),
    .ZN(_0428_));
 NOR2_X1 _5050_ (.A1(_0428_),
    .A2(_0412_),
    .ZN(_0429_));
 AOI21_X2 _5051_ (.A(_3207_),
    .B1(_0427_),
    .B2(_0429_),
    .ZN(_0430_));
 XNOR2_X2 _5052_ (.A(_0406_),
    .B(_0430_),
    .ZN(_3416_));
 XNOR2_X2 _5053_ (.A(_0419_),
    .B(_0418_),
    .ZN(_3420_));
 INV_X1 _5054_ (.A(_3215_),
    .ZN(_0431_));
 OAI221_X2 _5055_ (.A(_0431_),
    .B1(_0423_),
    .B2(_0424_),
    .C1(_0425_),
    .C2(_0426_),
    .ZN(_0432_));
 XOR2_X2 _5056_ (.A(_3212_),
    .B(_0432_),
    .Z(_3424_));
 OAI21_X1 _5057_ (.A(_0408_),
    .B1(_0410_),
    .B2(_0239_),
    .ZN(_0433_));
 AOI21_X2 _5058_ (.A(_3219_),
    .B1(_0433_),
    .B2(_0415_),
    .ZN(_0434_));
 XNOR2_X2 _5059_ (.A(_0414_),
    .B(_0434_),
    .ZN(_3428_));
 BUF_X8 _5060_ (.A(_0234_),
    .Z(_0435_));
 INV_X1 _5061_ (.A(_3136_),
    .ZN(_0436_));
 NAND3_X1 _5062_ (.A1(_0237_),
    .A2(_0415_),
    .A3(_0436_),
    .ZN(_0437_));
 AND3_X1 _5063_ (.A1(_0415_),
    .A2(_0238_),
    .A3(_0436_),
    .ZN(_0438_));
 OAI21_X2 _5064_ (.A(_0240_),
    .B1(_0422_),
    .B2(_0438_),
    .ZN(_0439_));
 NOR2_X1 _5065_ (.A1(_0415_),
    .A2(_0408_),
    .ZN(_0440_));
 OAI21_X1 _5066_ (.A(_0422_),
    .B1(_0415_),
    .B2(_0237_),
    .ZN(_0441_));
 AOI21_X2 _5067_ (.A(_0440_),
    .B1(_0441_),
    .B2(_0054_),
    .ZN(_0442_));
 NAND4_X4 _5068_ (.A1(_3245_),
    .A2(_0437_),
    .A3(_0439_),
    .A4(_0442_),
    .ZN(_0443_));
 NOR4_X4 _5069_ (.A1(_3420_),
    .A2(_3424_),
    .A3(_3428_),
    .A4(_0443_),
    .ZN(_0444_));
 INV_X1 _5070_ (.A(_0444_),
    .ZN(_0445_));
 OAI21_X1 _5071_ (.A(net18),
    .B1(_3416_),
    .B2(_0445_),
    .ZN(_0446_));
 XOR2_X2 _5072_ (.A(_3412_),
    .B(_0446_),
    .Z(_3221_));
 INV_X1 _5073_ (.A(_0332_),
    .ZN(_0447_));
 AOI21_X1 _5074_ (.A(_3095_),
    .B1(_2920_),
    .B2(_0196_),
    .ZN(_0448_));
 INV_X1 _5075_ (.A(_3092_),
    .ZN(_0449_));
 OAI21_X2 _5076_ (.A(_0198_),
    .B1(_0448_),
    .B2(_0449_),
    .ZN(_0450_));
 AOI21_X2 _5077_ (.A(_3087_),
    .B1(_0450_),
    .B2(_0203_),
    .ZN(_0451_));
 INV_X1 _5078_ (.A(_3084_),
    .ZN(_0452_));
 OAI21_X1 _5079_ (.A(_0447_),
    .B1(_0451_),
    .B2(_0452_),
    .ZN(_0453_));
 XNOR2_X2 _5080_ (.A(_0338_),
    .B(_0453_),
    .ZN(_3226_));
 OAI21_X2 _5081_ (.A(_0238_),
    .B1(_2915_),
    .B2(_0240_),
    .ZN(_0454_));
 AOI21_X2 _5082_ (.A(_3136_),
    .B1(_0454_),
    .B2(_0236_),
    .ZN(_0455_));
 XNOR2_X2 _5083_ (.A(_0415_),
    .B(_0455_),
    .ZN(_3296_));
 NOR2_X1 _5084_ (.A1(_3424_),
    .A2(_3428_),
    .ZN(_0456_));
 INV_X1 _5085_ (.A(_0456_),
    .ZN(_0457_));
 INV_X1 _5086_ (.A(_3296_),
    .ZN(_0458_));
 NAND2_X1 _5087_ (.A1(_3247_),
    .A2(_0458_),
    .ZN(_0459_));
 OR3_X1 _5088_ (.A1(_3420_),
    .A2(_0457_),
    .A3(_0459_),
    .ZN(_0460_));
 NAND2_X1 _5089_ (.A1(_0435_),
    .A2(_0460_),
    .ZN(_0461_));
 XOR2_X2 _5090_ (.A(_3416_),
    .B(_0461_),
    .Z(_3225_));
 OAI21_X1 _5091_ (.A(_0435_),
    .B1(_0443_),
    .B2(_0457_),
    .ZN(_0462_));
 XOR2_X2 _5092_ (.A(_3420_),
    .B(_0462_),
    .Z(_3229_));
 OAI21_X1 _5093_ (.A(_0435_),
    .B1(_3428_),
    .B2(_0459_),
    .ZN(_0463_));
 XOR2_X2 _5094_ (.A(_3424_),
    .B(_0463_),
    .Z(_3233_));
 NAND2_X1 _5095_ (.A1(_0435_),
    .A2(_0443_),
    .ZN(_0464_));
 XOR2_X2 _5096_ (.A(_3428_),
    .B(_0464_),
    .Z(_3237_));
 NOR2_X1 _5097_ (.A1(_3247_),
    .A2(_3261_),
    .ZN(_0465_));
 XNOR2_X1 _5098_ (.A(_3296_),
    .B(_0465_),
    .ZN(_3241_));
 MUX2_X1 _5099_ (.A(_3248_),
    .B(_3138_),
    .S(_0235_),
    .Z(_2935_));
 INV_X1 _5100_ (.A(_2935_),
    .ZN(_2939_));
 INV_X1 _5101_ (.A(_3239_),
    .ZN(_0466_));
 INV_X1 _5102_ (.A(_3249_),
    .ZN(_0467_));
 INV_X1 _5103_ (.A(_3250_),
    .ZN(_0468_));
 OAI21_X1 _5104_ (.A(_0467_),
    .B1(_0468_),
    .B2(_2934_),
    .ZN(_0469_));
 AOI21_X2 _5105_ (.A(_3243_),
    .B1(_0469_),
    .B2(_3244_),
    .ZN(_0470_));
 BUF_X2 _5106_ (.A(_3240_),
    .Z(_0471_));
 INV_X1 _5107_ (.A(_0471_),
    .ZN(_0472_));
 OAI21_X1 _5108_ (.A(_0466_),
    .B1(_0470_),
    .B2(_0472_),
    .ZN(_0473_));
 CLKBUF_X2 _5109_ (.A(_3236_),
    .Z(_0474_));
 AOI21_X2 _5110_ (.A(_3235_),
    .B1(_0473_),
    .B2(_0474_),
    .ZN(_0475_));
 XOR2_X2 _5111_ (.A(_3232_),
    .B(_0475_),
    .Z(_0476_));
 INV_X1 _5112_ (.A(_0476_),
    .ZN(_3448_));
 INV_X1 _5113_ (.A(_3243_),
    .ZN(_0477_));
 INV_X1 _5114_ (.A(_3244_),
    .ZN(_0478_));
 OAI21_X2 _5115_ (.A(_0477_),
    .B1(_0478_),
    .B2(_2937_),
    .ZN(_0479_));
 AOI21_X4 _5116_ (.A(_3239_),
    .B1(_0479_),
    .B2(_0471_),
    .ZN(_0480_));
 XNOR2_X2 _5117_ (.A(_0474_),
    .B(_0480_),
    .ZN(_3452_));
 INV_X1 _5118_ (.A(_3452_),
    .ZN(_3311_));
 XNOR2_X2 _5119_ (.A(_0471_),
    .B(_0470_),
    .ZN(_3456_));
 INV_X1 _5120_ (.A(_3456_),
    .ZN(_3310_));
 OR3_X1 _5121_ (.A1(_3227_),
    .A2(_3231_),
    .A3(_3235_),
    .ZN(_0481_));
 AOI21_X1 _5122_ (.A(_0481_),
    .B1(_0473_),
    .B2(_0474_),
    .ZN(_0482_));
 OAI21_X1 _5123_ (.A(_3228_),
    .B1(_3232_),
    .B2(_3231_),
    .ZN(_0483_));
 INV_X1 _5124_ (.A(_0483_),
    .ZN(_0484_));
 NOR2_X1 _5125_ (.A1(_3227_),
    .A2(_0484_),
    .ZN(_0485_));
 OAI21_X1 _5126_ (.A(_3224_),
    .B1(_0482_),
    .B2(_0485_),
    .ZN(_0486_));
 OR3_X1 _5127_ (.A1(_3224_),
    .A2(_0482_),
    .A3(_0485_),
    .ZN(_0487_));
 AND2_X1 _5128_ (.A1(_0486_),
    .A2(_0487_),
    .ZN(_0488_));
 INV_X1 _5129_ (.A(_0488_),
    .ZN(_3440_));
 INV_X4 _5130_ (.A(net48),
    .ZN(_3289_));
 MUX2_X1 _5131_ (.A(net48),
    .B(_3291_),
    .S(_0042_),
    .Z(_3292_));
 INV_X1 _5132_ (.A(_3292_),
    .ZN(_2941_));
 NOR3_X1 _5133_ (.A1(_3265_),
    .A2(_3268_),
    .A3(_3271_),
    .ZN(_0489_));
 INV_X1 _5134_ (.A(_0489_),
    .ZN(_0490_));
 OAI21_X1 _5135_ (.A(_3272_),
    .B1(_3275_),
    .B2(_3274_),
    .ZN(_0491_));
 INV_X1 _5136_ (.A(_0491_),
    .ZN(_0492_));
 NOR2_X1 _5137_ (.A1(_3274_),
    .A2(_3277_),
    .ZN(_0493_));
 INV_X1 _5138_ (.A(_3283_),
    .ZN(_0494_));
 INV_X1 _5139_ (.A(_3287_),
    .ZN(_0495_));
 AOI21_X2 _5140_ (.A(_3293_),
    .B1(_3294_),
    .B2(_0005_),
    .ZN(_0496_));
 INV_X2 _5141_ (.A(_3288_),
    .ZN(_0497_));
 OAI21_X4 _5142_ (.A(_0495_),
    .B1(_0496_),
    .B2(_0497_),
    .ZN(_0498_));
 AOI21_X4 _5143_ (.A(_3285_),
    .B1(_3286_),
    .B2(_0498_),
    .ZN(_0499_));
 INV_X1 _5144_ (.A(_3284_),
    .ZN(_0500_));
 OAI21_X4 _5145_ (.A(_0494_),
    .B1(_0499_),
    .B2(_0500_),
    .ZN(_0501_));
 AOI21_X4 _5146_ (.A(_3280_),
    .B1(_0501_),
    .B2(_3281_),
    .ZN(_0502_));
 INV_X1 _5147_ (.A(_3278_),
    .ZN(_0503_));
 OAI21_X4 _5148_ (.A(_0493_),
    .B1(_0502_),
    .B2(_0503_),
    .ZN(_0504_));
 AOI21_X4 _5149_ (.A(_0490_),
    .B1(_0504_),
    .B2(_0492_),
    .ZN(_0505_));
 OR3_X1 _5150_ (.A1(_3269_),
    .A2(_3265_),
    .A3(_3268_),
    .ZN(_0506_));
 OAI21_X1 _5151_ (.A(_0506_),
    .B1(_3265_),
    .B2(_3266_),
    .ZN(_0507_));
 BUF_X1 _5152_ (.A(_3263_),
    .Z(_0508_));
 BUF_X1 _5153_ (.A(_3259_),
    .Z(_0509_));
 NAND4_X1 _5154_ (.A1(_3253_),
    .A2(_0508_),
    .A3(_3256_),
    .A4(_0509_),
    .ZN(_0510_));
 OR3_X4 _5155_ (.A1(_0510_),
    .A2(_0507_),
    .A3(_0505_),
    .ZN(_0511_));
 INV_X1 _5156_ (.A(_3255_),
    .ZN(_0512_));
 AOI21_X1 _5157_ (.A(_3258_),
    .B1(_3262_),
    .B2(_0509_),
    .ZN(_0513_));
 INV_X1 _5158_ (.A(_3256_),
    .ZN(_0514_));
 OAI21_X2 _5159_ (.A(_0512_),
    .B1(_0513_),
    .B2(_0514_),
    .ZN(_0515_));
 AOI21_X4 _5160_ (.A(_3252_),
    .B1(_0515_),
    .B2(_3253_),
    .ZN(_0516_));
 NAND2_X4 _5161_ (.A1(_0511_),
    .A2(_0516_),
    .ZN(_0517_));
 INV_X1 _5162_ (.A(_0517_),
    .ZN(_0518_));
 BUF_X4 _5163_ (.A(_0518_),
    .Z(_0519_));
 BUF_X4 _5164_ (.A(_0519_),
    .Z(_3483_));
 INV_X1 _5165_ (.A(_3140_),
    .ZN(_0520_));
 AOI21_X1 _5166_ (.A(_3143_),
    .B1(_2932_),
    .B2(_3144_),
    .ZN(_0521_));
 INV_X1 _5167_ (.A(_0242_),
    .ZN(_0522_));
 OAI21_X2 _5168_ (.A(_0520_),
    .B1(_0521_),
    .B2(_0522_),
    .ZN(_0523_));
 XNOR2_X2 _5169_ (.A(_3298_),
    .B(_0523_),
    .ZN(_3463_));
 INV_X1 _5170_ (.A(_3304_),
    .ZN(_0524_));
 AOI21_X1 _5171_ (.A(_3308_),
    .B1(_3309_),
    .B2(_2947_),
    .ZN(_0525_));
 INV_X1 _5172_ (.A(_3305_),
    .ZN(_0526_));
 OAI21_X2 _5173_ (.A(_0524_),
    .B1(_0525_),
    .B2(_0526_),
    .ZN(_0527_));
 XNOR2_X2 _5174_ (.A(_3302_),
    .B(_0527_),
    .ZN(_3660_));
 OR3_X1 _5175_ (.A1(_0342_),
    .A2(_0373_),
    .A3(_0351_),
    .ZN(_0528_));
 NAND2_X1 _5176_ (.A1(_0366_),
    .A2(_0345_),
    .ZN(_0529_));
 AND2_X1 _5177_ (.A1(_0349_),
    .A2(_0350_),
    .ZN(_0530_));
 NAND4_X1 _5178_ (.A1(_0342_),
    .A2(_0349_),
    .A3(_0350_),
    .A4(_0351_),
    .ZN(_0531_));
 OAI221_X2 _5179_ (.A(_0528_),
    .B1(_0529_),
    .B2(_0530_),
    .C1(_0285_),
    .C2(_0531_),
    .ZN(_0532_));
 NAND2_X1 _5180_ (.A1(_0342_),
    .A2(_0373_),
    .ZN(_0533_));
 OAI21_X2 _5181_ (.A(_0533_),
    .B1(_0529_),
    .B2(_0375_),
    .ZN(_0534_));
 OR2_X1 _5182_ (.A1(_0532_),
    .A2(_0534_),
    .ZN(_0535_));
 NAND2_X1 _5183_ (.A1(_0279_),
    .A2(_0276_),
    .ZN(_0536_));
 AOI21_X2 _5184_ (.A(_3193_),
    .B1(_3169_),
    .B2(_3191_),
    .ZN(_0537_));
 NAND2_X1 _5185_ (.A1(_0366_),
    .A2(_0537_),
    .ZN(_0538_));
 AOI211_X2 _5186_ (.A(_0536_),
    .B(_0538_),
    .C1(_0118_),
    .C2(_0120_),
    .ZN(_0539_));
 OR2_X1 _5187_ (.A1(_0366_),
    .A2(_0537_),
    .ZN(_0540_));
 OR2_X1 _5188_ (.A1(_0342_),
    .A2(_0356_),
    .ZN(_0541_));
 INV_X1 _5189_ (.A(_0537_),
    .ZN(_0542_));
 OAI221_X2 _5190_ (.A(_0540_),
    .B1(_0541_),
    .B2(_0542_),
    .C1(_0538_),
    .C2(_0278_),
    .ZN(_0543_));
 AND3_X1 _5191_ (.A1(_0342_),
    .A2(_0278_),
    .A3(_0356_),
    .ZN(_0544_));
 AOI211_X2 _5192_ (.A(_0539_),
    .B(_0543_),
    .C1(_0544_),
    .C2(_0281_),
    .ZN(_0545_));
 MUX2_X2 _5193_ (.A(_0535_),
    .B(_0545_),
    .S(_0015_),
    .Z(_3348_));
 NOR3_X1 _5194_ (.A1(_3202_),
    .A2(_0309_),
    .A3(_3197_),
    .ZN(_0546_));
 OR2_X1 _5195_ (.A1(_0053_),
    .A2(_0546_),
    .ZN(_0547_));
 XOR2_X2 _5196_ (.A(_3348_),
    .B(_0547_),
    .Z(_3319_));
 OR3_X1 _5197_ (.A1(_3202_),
    .A2(_3206_),
    .A3(_0327_),
    .ZN(_0548_));
 NAND2_X1 _5198_ (.A1(_0179_),
    .A2(_0548_),
    .ZN(_0549_));
 XOR2_X1 _5199_ (.A(_3197_),
    .B(_0549_),
    .Z(_3323_));
 INV_X1 _5200_ (.A(_3322_),
    .ZN(_0550_));
 NAND2_X2 _5201_ (.A1(_0329_),
    .A2(_3326_),
    .ZN(_0551_));
 NOR3_X4 _5202_ (.A1(_0551_),
    .A2(_0550_),
    .A3(_0338_),
    .ZN(_0552_));
 NAND3_X2 _5203_ (.A1(_0334_),
    .A2(_0336_),
    .A3(_0552_),
    .ZN(_0553_));
 INV_X1 _5204_ (.A(_3325_),
    .ZN(_0554_));
 CLKBUF_X2 _5205_ (.A(_3175_),
    .Z(_0555_));
 AOI21_X1 _5206_ (.A(_0555_),
    .B1(_0330_),
    .B2(_0329_),
    .ZN(_0556_));
 INV_X1 _5207_ (.A(_3326_),
    .ZN(_0557_));
 OAI21_X1 _5208_ (.A(_0554_),
    .B1(_0556_),
    .B2(_0557_),
    .ZN(_0558_));
 AOI22_X2 _5209_ (.A1(_3322_),
    .A2(_0558_),
    .B1(_0552_),
    .B2(_0332_),
    .ZN(_0559_));
 AND2_X1 _5210_ (.A1(_0553_),
    .A2(_0559_),
    .ZN(_0560_));
 OR2_X1 _5211_ (.A1(_3322_),
    .A2(_0558_),
    .ZN(_0561_));
 NOR3_X1 _5212_ (.A1(_0338_),
    .A2(_0337_),
    .A3(_0551_),
    .ZN(_0562_));
 OAI21_X2 _5213_ (.A(_0560_),
    .B1(_0561_),
    .B2(_0562_),
    .ZN(_0563_));
 INV_X2 _5214_ (.A(_0563_),
    .ZN(_3352_));
 BUF_X4 _5215_ (.A(_3329_),
    .Z(_0564_));
 INV_X2 _5216_ (.A(_0564_),
    .ZN(_0565_));
 CLKBUF_X2 _5217_ (.A(_3337_),
    .Z(_0566_));
 INV_X2 _5218_ (.A(_0566_),
    .ZN(_0567_));
 BUF_X2 _5219_ (.A(_3187_),
    .Z(_0568_));
 AOI21_X2 _5220_ (.A(_3341_),
    .B1(_0567_),
    .B2(_0568_),
    .ZN(_0569_));
 INV_X1 _5221_ (.A(_0569_),
    .ZN(_0570_));
 BUF_X4 _5222_ (.A(_0566_),
    .Z(_0571_));
 NOR2_X1 _5223_ (.A1(_0342_),
    .A2(_0571_),
    .ZN(_0572_));
 OAI21_X1 _5224_ (.A(_0345_),
    .B1(_0352_),
    .B2(_0285_),
    .ZN(_0573_));
 AOI21_X2 _5225_ (.A(_0570_),
    .B1(_0572_),
    .B2(_0573_),
    .ZN(_0574_));
 AOI21_X1 _5226_ (.A(_3336_),
    .B1(_3182_),
    .B2(_0571_),
    .ZN(_0575_));
 NAND2_X1 _5227_ (.A1(_0342_),
    .A2(_0571_),
    .ZN(_0576_));
 OAI21_X1 _5228_ (.A(_0575_),
    .B1(_0576_),
    .B2(_0364_),
    .ZN(_0577_));
 MUX2_X1 _5229_ (.A(_0574_),
    .B(_0577_),
    .S(_0019_),
    .Z(_0578_));
 XNOR2_X2 _5230_ (.A(_0565_),
    .B(_0578_),
    .ZN(_3384_));
 OR3_X1 _5231_ (.A1(_0263_),
    .A2(_0568_),
    .A3(_0343_),
    .ZN(_0579_));
 AOI211_X2 _5232_ (.A(_3171_),
    .B(_0579_),
    .C1(_0283_),
    .C2(_0274_),
    .ZN(_0580_));
 OAI221_X2 _5233_ (.A(_0580_),
    .B1(_0269_),
    .B2(_0268_),
    .C1(_0266_),
    .C2(_0035_),
    .ZN(_0581_));
 INV_X1 _5234_ (.A(_0568_),
    .ZN(_0582_));
 OAI21_X2 _5235_ (.A(_0366_),
    .B1(_0343_),
    .B2(_0344_),
    .ZN(_0583_));
 NOR3_X2 _5236_ (.A1(_0568_),
    .A2(_0343_),
    .A3(_0380_),
    .ZN(_0584_));
 AOI21_X2 _5237_ (.A(_3171_),
    .B1(_0274_),
    .B2(_0283_),
    .ZN(_0585_));
 AOI22_X4 _5238_ (.A1(_0582_),
    .A2(_0583_),
    .B1(_0584_),
    .B2(_0585_),
    .ZN(_0586_));
 NAND2_X1 _5239_ (.A1(_0586_),
    .A2(_0581_),
    .ZN(_0587_));
 AOI21_X1 _5240_ (.A(_3182_),
    .B1(_3190_),
    .B2(_0341_),
    .ZN(_0588_));
 NAND2_X1 _5241_ (.A1(_0347_),
    .A2(_0341_),
    .ZN(_0589_));
 OAI21_X2 _5242_ (.A(_0588_),
    .B1(_0589_),
    .B2(_0389_),
    .ZN(_0590_));
 INV_X1 _5243_ (.A(_0590_),
    .ZN(_0591_));
 AND4_X1 _5244_ (.A1(_0247_),
    .A2(_0346_),
    .A3(_0347_),
    .A4(_0341_),
    .ZN(_0592_));
 NAND2_X1 _5245_ (.A1(_0255_),
    .A2(_0592_),
    .ZN(_0593_));
 OAI21_X1 _5246_ (.A(_0591_),
    .B1(_0593_),
    .B2(_0260_),
    .ZN(_0594_));
 MUX2_X1 _5247_ (.A(_0587_),
    .B(_0594_),
    .S(_0017_),
    .Z(_0595_));
 XNOR2_X2 _5248_ (.A(_0595_),
    .B(_0567_),
    .ZN(_3392_));
 AND2_X1 _5249_ (.A1(_3161_),
    .A2(_0346_),
    .ZN(_0596_));
 OR2_X1 _5250_ (.A1(_3169_),
    .A2(_3193_),
    .ZN(_0597_));
 OAI221_X2 _5251_ (.A(_0342_),
    .B1(_0596_),
    .B2(_0597_),
    .C1(_3193_),
    .C2(_0347_),
    .ZN(_0598_));
 AOI21_X1 _5252_ (.A(_3185_),
    .B1(_0592_),
    .B2(_0275_),
    .ZN(_0599_));
 AND2_X1 _5253_ (.A1(_0598_),
    .A2(_0599_),
    .ZN(_0600_));
 NAND3_X2 _5254_ (.A1(_0108_),
    .A2(_0296_),
    .A3(_0592_),
    .ZN(_0601_));
 OAI21_X4 _5255_ (.A(_0600_),
    .B1(_0601_),
    .B2(_0293_),
    .ZN(_0602_));
 MUX2_X1 _5256_ (.A(_0587_),
    .B(_0602_),
    .S(_2909_),
    .Z(_0603_));
 XNOR2_X1 _5257_ (.A(_0571_),
    .B(_0603_),
    .ZN(_0604_));
 INV_X1 _5258_ (.A(_0604_),
    .ZN(_3343_));
 BUF_X2 _5259_ (.A(_3349_),
    .Z(_0605_));
 INV_X1 _5260_ (.A(_3199_),
    .ZN(_0606_));
 OAI21_X2 _5261_ (.A(_0606_),
    .B1(_0407_),
    .B2(_0405_),
    .ZN(_0607_));
 CLKBUF_X2 _5262_ (.A(_3350_),
    .Z(_0608_));
 AOI21_X1 _5263_ (.A(_0605_),
    .B1(_0607_),
    .B2(_0608_),
    .ZN(_0609_));
 NAND4_X1 _5264_ (.A1(_0406_),
    .A2(_3200_),
    .A3(_0419_),
    .A4(_0608_),
    .ZN(_0610_));
 OAI21_X1 _5265_ (.A(_0609_),
    .B1(_0610_),
    .B2(_0418_),
    .ZN(_0611_));
 XOR2_X2 _5266_ (.A(_3346_),
    .B(_0611_),
    .Z(_3404_));
 NAND3_X1 _5267_ (.A1(_0406_),
    .A2(_3200_),
    .A3(_0419_),
    .ZN(_0612_));
 NOR2_X1 _5268_ (.A1(_0412_),
    .A2(_0612_),
    .ZN(_0613_));
 AOI21_X2 _5269_ (.A(_0607_),
    .B1(_0613_),
    .B2(_0427_),
    .ZN(_0614_));
 XNOR2_X2 _5270_ (.A(_0608_),
    .B(_0614_),
    .ZN(_3408_));
 NOR3_X1 _5271_ (.A1(_3412_),
    .A2(_3416_),
    .A3(_3408_),
    .ZN(_0615_));
 AOI21_X1 _5272_ (.A(_0235_),
    .B1(_0444_),
    .B2(_0615_),
    .ZN(_0616_));
 XNOR2_X1 _5273_ (.A(_3404_),
    .B(_0616_),
    .ZN(_3351_));
 NOR3_X1 _5274_ (.A1(_0332_),
    .A2(_0555_),
    .A3(_0330_),
    .ZN(_0617_));
 OAI21_X1 _5275_ (.A(_0617_),
    .B1(_0451_),
    .B2(_0452_),
    .ZN(_0618_));
 OR2_X1 _5276_ (.A1(_3180_),
    .A2(_0555_),
    .ZN(_0619_));
 OAI221_X2 _5277_ (.A(_0618_),
    .B1(_0619_),
    .B2(_0330_),
    .C1(_0555_),
    .C2(_0329_),
    .ZN(_0620_));
 XNOR2_X2 _5278_ (.A(_0557_),
    .B(_0620_),
    .ZN(_0621_));
 INV_X1 _5279_ (.A(_0621_),
    .ZN(_3356_));
 NOR3_X1 _5280_ (.A1(_3412_),
    .A2(_3416_),
    .A3(_0460_),
    .ZN(_0622_));
 NOR2_X1 _5281_ (.A1(net17),
    .A2(_0622_),
    .ZN(_0623_));
 XNOR2_X1 _5282_ (.A(_3408_),
    .B(_0623_),
    .ZN(_3355_));
 CLKBUF_X2 _5283_ (.A(_3354_),
    .Z(_0624_));
 NOR3_X1 _5284_ (.A1(_3227_),
    .A2(_3231_),
    .A3(_3235_),
    .ZN(_0625_));
 NOR2_X2 _5285_ (.A1(_3223_),
    .A2(_3357_),
    .ZN(_0626_));
 AND2_X1 _5286_ (.A1(_0625_),
    .A2(_0626_),
    .ZN(_0627_));
 INV_X1 _5287_ (.A(_2934_),
    .ZN(_0628_));
 AOI21_X1 _5288_ (.A(_3249_),
    .B1(_3250_),
    .B2(_0628_),
    .ZN(_0629_));
 OAI21_X1 _5289_ (.A(_0477_),
    .B1(_0629_),
    .B2(_0478_),
    .ZN(_0630_));
 AOI21_X1 _5290_ (.A(_3239_),
    .B1(_0630_),
    .B2(_0471_),
    .ZN(_0631_));
 INV_X1 _5291_ (.A(_0474_),
    .ZN(_0632_));
 OAI21_X2 _5292_ (.A(_0627_),
    .B1(_0631_),
    .B2(_0632_),
    .ZN(_0633_));
 NOR2_X1 _5293_ (.A1(_3358_),
    .A2(_3357_),
    .ZN(_0634_));
 OAI21_X2 _5294_ (.A(_3224_),
    .B1(_3227_),
    .B2(_0484_),
    .ZN(_0635_));
 AOI21_X4 _5295_ (.A(_0634_),
    .B1(_0626_),
    .B2(_0635_),
    .ZN(_0636_));
 AND3_X1 _5296_ (.A1(_0624_),
    .A2(_0633_),
    .A3(_0636_),
    .ZN(_0637_));
 AOI21_X2 _5297_ (.A(_0624_),
    .B1(_0633_),
    .B2(_0636_),
    .ZN(_0638_));
 NOR2_X2 _5298_ (.A1(_0637_),
    .A2(_0638_),
    .ZN(_3432_));
 BUF_X2 _5299_ (.A(_3361_),
    .Z(_0639_));
 CLKBUF_X2 _5300_ (.A(_3369_),
    .Z(_0640_));
 CLKBUF_X3 _5301_ (.A(_0640_),
    .Z(_0641_));
 AOI21_X1 _5302_ (.A(_3368_),
    .B1(_3328_),
    .B2(_0641_),
    .ZN(_0642_));
 NAND4_X2 _5303_ (.A1(_0341_),
    .A2(_0566_),
    .A3(_0564_),
    .A4(_0640_),
    .ZN(_0643_));
 NAND2_X1 _5304_ (.A1(_0564_),
    .A2(_0641_),
    .ZN(_0644_));
 OAI221_X1 _5305_ (.A(_0642_),
    .B1(_0643_),
    .B2(_0354_),
    .C1(_0575_),
    .C2(_0644_),
    .ZN(_0645_));
 INV_X1 _5306_ (.A(_0645_),
    .ZN(_0646_));
 NOR3_X1 _5307_ (.A1(_0274_),
    .A2(_0344_),
    .A3(_0643_),
    .ZN(_0647_));
 NAND2_X1 _5308_ (.A1(_0359_),
    .A2(_0647_),
    .ZN(_0648_));
 OAI211_X2 _5309_ (.A(_0017_),
    .B(_0646_),
    .C1(_0648_),
    .C2(_0369_),
    .ZN(_0649_));
 INV_X2 _5310_ (.A(_0640_),
    .ZN(_0650_));
 AOI21_X1 _5311_ (.A(_3373_),
    .B1(_0650_),
    .B2(_3333_),
    .ZN(_0651_));
 OR4_X1 _5312_ (.A1(_0341_),
    .A2(_0566_),
    .A3(_0564_),
    .A4(_0640_),
    .ZN(_0652_));
 NAND2_X1 _5313_ (.A1(_0565_),
    .A2(_0650_),
    .ZN(_0653_));
 OAI221_X1 _5314_ (.A(_0651_),
    .B1(_0652_),
    .B2(_0345_),
    .C1(_0569_),
    .C2(_0653_),
    .ZN(_0654_));
 AOI21_X1 _5315_ (.A(_0652_),
    .B1(_0284_),
    .B2(_0058_),
    .ZN(_0655_));
 AND3_X1 _5316_ (.A1(_0349_),
    .A2(_0350_),
    .A3(_0655_),
    .ZN(_0656_));
 AOI21_X1 _5317_ (.A(_0654_),
    .B1(_0656_),
    .B2(_0375_),
    .ZN(_0657_));
 OAI21_X1 _5318_ (.A(_0649_),
    .B1(_0657_),
    .B2(_0018_),
    .ZN(_0658_));
 XNOR2_X2 _5319_ (.A(_0639_),
    .B(_0658_),
    .ZN(_3376_));
 INV_X2 _5320_ (.A(_0639_),
    .ZN(_0659_));
 INV_X1 _5321_ (.A(_3371_),
    .ZN(_0660_));
 OAI21_X1 _5322_ (.A(_0660_),
    .B1(_0537_),
    .B2(_0643_),
    .ZN(_0661_));
 AOI21_X2 _5323_ (.A(_3331_),
    .B1(_3339_),
    .B2(_0564_),
    .ZN(_0662_));
 NAND2_X2 _5324_ (.A1(_0571_),
    .A2(_0564_),
    .ZN(_0663_));
 INV_X1 _5325_ (.A(_3185_),
    .ZN(_0664_));
 OAI21_X1 _5326_ (.A(_0662_),
    .B1(_0663_),
    .B2(_0664_),
    .ZN(_0665_));
 AOI21_X1 _5327_ (.A(_0661_),
    .B1(_0665_),
    .B2(_0641_),
    .ZN(_0666_));
 NAND2_X1 _5328_ (.A1(_0278_),
    .A2(_0647_),
    .ZN(_0667_));
 AOI21_X1 _5329_ (.A(_0536_),
    .B1(_0120_),
    .B2(_0118_),
    .ZN(_0668_));
 OAI21_X1 _5330_ (.A(_0666_),
    .B1(_0667_),
    .B2(_0668_),
    .ZN(_0669_));
 MUX2_X1 _5331_ (.A(_0657_),
    .B(_0669_),
    .S(_0015_),
    .Z(_0670_));
 XNOR2_X2 _5332_ (.A(_0659_),
    .B(_0670_),
    .ZN(_3554_));
 NAND2_X1 _5333_ (.A1(_0650_),
    .A2(_0017_),
    .ZN(_0671_));
 NAND2_X1 _5334_ (.A1(_0641_),
    .A2(_0019_),
    .ZN(_0672_));
 AOI21_X2 _5335_ (.A(_3333_),
    .B1(_3341_),
    .B2(_0565_),
    .ZN(_0673_));
 NOR2_X1 _5336_ (.A1(_0571_),
    .A2(_0564_),
    .ZN(_0674_));
 OR3_X1 _5337_ (.A1(_0568_),
    .A2(_0343_),
    .A3(_0380_),
    .ZN(_0675_));
 AOI21_X1 _5338_ (.A(_0341_),
    .B1(_0371_),
    .B2(_0347_),
    .ZN(_0676_));
 OAI221_X1 _5339_ (.A(_0674_),
    .B1(_0675_),
    .B2(_0379_),
    .C1(_0568_),
    .C2(_0676_),
    .ZN(_0677_));
 NOR3_X1 _5340_ (.A1(_0263_),
    .A2(_0568_),
    .A3(_0343_),
    .ZN(_0678_));
 OAI211_X2 _5341_ (.A(_0372_),
    .B(_0678_),
    .C1(_0288_),
    .C2(_0273_),
    .ZN(_0679_));
 AOI221_X2 _5342_ (.A(_0679_),
    .B1(_0286_),
    .B2(_0384_),
    .C1(_0065_),
    .C2(_0386_),
    .ZN(_0680_));
 OAI21_X1 _5343_ (.A(_0673_),
    .B1(_0677_),
    .B2(_0680_),
    .ZN(_0681_));
 MUX2_X1 _5344_ (.A(_0671_),
    .B(_0672_),
    .S(_0681_),
    .Z(_0682_));
 AND2_X1 _5345_ (.A1(_0663_),
    .A2(_0662_),
    .ZN(_0683_));
 NAND3_X1 _5346_ (.A1(_0598_),
    .A2(_0599_),
    .A3(_0662_),
    .ZN(_0684_));
 AND3_X1 _5347_ (.A1(_0108_),
    .A2(_0296_),
    .A3(_0592_),
    .ZN(_0685_));
 AOI21_X2 _5348_ (.A(_0684_),
    .B1(_0685_),
    .B2(_0400_),
    .ZN(_0686_));
 OR4_X2 _5349_ (.A1(_0641_),
    .A2(_0019_),
    .A3(_0683_),
    .A4(_0686_),
    .ZN(_0687_));
 NOR2_X1 _5350_ (.A1(_0650_),
    .A2(_0017_),
    .ZN(_0688_));
 OAI21_X2 _5351_ (.A(_0688_),
    .B1(_0686_),
    .B2(_0683_),
    .ZN(_0689_));
 NAND3_X4 _5352_ (.A1(_0682_),
    .A2(_0687_),
    .A3(_0689_),
    .ZN(_3542_));
 NOR3_X1 _5353_ (.A1(_3185_),
    .A2(_3339_),
    .A3(_0542_),
    .ZN(_0690_));
 NAND2_X1 _5354_ (.A1(_0278_),
    .A2(_0356_),
    .ZN(_0691_));
 OAI21_X1 _5355_ (.A(_0690_),
    .B1(_0691_),
    .B2(_0668_),
    .ZN(_0692_));
 INV_X1 _5356_ (.A(_3339_),
    .ZN(_0693_));
 NOR2_X1 _5357_ (.A1(_0342_),
    .A2(_3185_),
    .ZN(_0694_));
 OAI21_X1 _5358_ (.A(_0693_),
    .B1(_0694_),
    .B2(_0567_),
    .ZN(_0695_));
 AND3_X1 _5359_ (.A1(_0015_),
    .A2(_0692_),
    .A3(_0695_),
    .ZN(_0696_));
 AOI21_X2 _5360_ (.A(_0696_),
    .B1(_0574_),
    .B2(_0019_),
    .ZN(_0697_));
 XNOR2_X2 _5361_ (.A(_0565_),
    .B(_0697_),
    .ZN(_0698_));
 INV_X2 _5362_ (.A(_0698_),
    .ZN(_3396_));
 XNOR2_X2 _5363_ (.A(net13),
    .B(net31),
    .ZN(_0699_));
 OAI21_X1 _5364_ (.A(_0660_),
    .B1(_0662_),
    .B2(_0650_),
    .ZN(_0700_));
 AND2_X1 _5365_ (.A1(_0639_),
    .A2(_0700_),
    .ZN(_0701_));
 OR3_X1 _5366_ (.A1(_3363_),
    .A2(_0017_),
    .A3(_0701_),
    .ZN(_0702_));
 NOR3_X2 _5367_ (.A1(_0650_),
    .A2(_0659_),
    .A3(_0663_),
    .ZN(_0703_));
 AOI21_X4 _5368_ (.A(_0702_),
    .B1(_0703_),
    .B2(_0602_),
    .ZN(_0704_));
 OAI21_X2 _5369_ (.A(_0018_),
    .B1(_3365_),
    .B2(_0659_),
    .ZN(_0705_));
 NOR2_X1 _5370_ (.A1(_3365_),
    .A2(_3373_),
    .ZN(_0706_));
 OAI21_X2 _5371_ (.A(_0706_),
    .B1(_0673_),
    .B2(_0641_),
    .ZN(_0707_));
 INV_X1 _5372_ (.A(_0707_),
    .ZN(_0708_));
 NOR3_X2 _5373_ (.A1(_0571_),
    .A2(_0564_),
    .A3(_0641_),
    .ZN(_0709_));
 NAND3_X2 _5374_ (.A1(_0581_),
    .A2(_0586_),
    .A3(_0709_),
    .ZN(_0710_));
 AOI21_X4 _5375_ (.A(_0705_),
    .B1(_0708_),
    .B2(_0710_),
    .ZN(_0711_));
 NOR2_X2 _5376_ (.A1(_0704_),
    .A2(_0711_),
    .ZN(_0712_));
 XNOR2_X1 _5377_ (.A(_0699_),
    .B(_0712_),
    .ZN(_0713_));
 OR2_X1 _5378_ (.A1(_3554_),
    .A2(_3542_),
    .ZN(_0714_));
 NOR3_X1 _5379_ (.A1(_3197_),
    .A2(_3348_),
    .A3(_0548_),
    .ZN(_0715_));
 NAND3_X1 _5380_ (.A1(_0604_),
    .A2(_0698_),
    .A3(_0715_),
    .ZN(_0716_));
 OAI21_X1 _5381_ (.A(_0191_),
    .B1(_0714_),
    .B2(_0716_),
    .ZN(_0717_));
 XNOR2_X1 _5382_ (.A(_0713_),
    .B(_0717_),
    .ZN(_3375_));
 AOI21_X2 _5383_ (.A(_3328_),
    .B1(_3336_),
    .B2(_0564_),
    .ZN(_0718_));
 NAND2_X1 _5384_ (.A1(_0663_),
    .A2(_0718_),
    .ZN(_0719_));
 INV_X1 _5385_ (.A(_0718_),
    .ZN(_0720_));
 NOR2_X1 _5386_ (.A1(_0590_),
    .A2(_0720_),
    .ZN(_0721_));
 OAI21_X1 _5387_ (.A(_0721_),
    .B1(_0593_),
    .B2(_0260_),
    .ZN(_0722_));
 AND4_X1 _5388_ (.A1(_0641_),
    .A2(_0018_),
    .A3(_0719_),
    .A4(_0722_),
    .ZN(_0723_));
 AOI21_X2 _5389_ (.A(_0671_),
    .B1(_0719_),
    .B2(_0722_),
    .ZN(_0724_));
 NOR2_X1 _5390_ (.A1(_0641_),
    .A2(_0017_),
    .ZN(_0725_));
 MUX2_X1 _5391_ (.A(_0688_),
    .B(_0725_),
    .S(_0681_),
    .Z(_0726_));
 NOR3_X4 _5392_ (.A1(_0723_),
    .A2(_0724_),
    .A3(_0726_),
    .ZN(_3380_));
 NAND2_X1 _5393_ (.A1(_0598_),
    .A2(_0599_),
    .ZN(_0727_));
 AOI21_X2 _5394_ (.A(_0727_),
    .B1(_0685_),
    .B2(_0400_),
    .ZN(_0728_));
 NOR4_X2 _5395_ (.A1(_0567_),
    .A2(_0019_),
    .A3(_0545_),
    .A4(_0728_),
    .ZN(_0729_));
 NOR4_X2 _5396_ (.A1(_0571_),
    .A2(_0019_),
    .A3(_0545_),
    .A4(_0602_),
    .ZN(_0730_));
 OAI22_X1 _5397_ (.A1(_0568_),
    .A2(_0676_),
    .B1(_0675_),
    .B2(_0379_),
    .ZN(_0731_));
 OAI21_X1 _5398_ (.A(_0571_),
    .B1(_0680_),
    .B2(_0731_),
    .ZN(_0732_));
 NOR4_X2 _5399_ (.A1(_0015_),
    .A2(_0532_),
    .A3(_0534_),
    .A4(_0732_),
    .ZN(_0733_));
 NAND3_X1 _5400_ (.A1(_0567_),
    .A2(_0581_),
    .A3(_0586_),
    .ZN(_0734_));
 NOR4_X2 _5401_ (.A1(_0015_),
    .A2(_0532_),
    .A3(_0534_),
    .A4(_0734_),
    .ZN(_0735_));
 NOR4_X2 _5402_ (.A1(_0729_),
    .A2(_0730_),
    .A3(_0733_),
    .A4(_0735_),
    .ZN(_0736_));
 OR4_X2 _5403_ (.A1(_3202_),
    .A2(_0309_),
    .A3(_3197_),
    .A4(_0736_),
    .ZN(_0737_));
 NOR3_X1 _5404_ (.A1(_3542_),
    .A2(_3396_),
    .A3(_0737_),
    .ZN(_0738_));
 NOR2_X1 _5405_ (.A1(net227),
    .A2(_0738_),
    .ZN(_0739_));
 XNOR2_X1 _5406_ (.A(_3554_),
    .B(_0739_),
    .ZN(_3379_));
 NAND2_X1 _5407_ (.A1(_0179_),
    .A2(_0716_),
    .ZN(_0740_));
 XOR2_X1 _5408_ (.A(_3542_),
    .B(_0740_),
    .Z(_3383_));
 NOR4_X2 _5409_ (.A1(_3202_),
    .A2(_0309_),
    .A3(_3197_),
    .A4(_0736_),
    .ZN(_0741_));
 NOR2_X1 _5410_ (.A1(net227),
    .A2(_0741_),
    .ZN(_0742_));
 XNOR2_X1 _5411_ (.A(_3396_),
    .B(_0742_),
    .ZN(_3391_));
 NOR2_X1 _5412_ (.A1(net227),
    .A2(_0715_),
    .ZN(_0743_));
 XNOR2_X1 _5413_ (.A(_3343_),
    .B(_0743_),
    .ZN(_3387_));
 INV_X1 _5414_ (.A(_3385_),
    .ZN(_0744_));
 CLKBUF_X2 _5415_ (.A(_3394_),
    .Z(_0745_));
 CLKBUF_X2 _5416_ (.A(_3386_),
    .Z(_0746_));
 AND3_X1 _5417_ (.A1(_0745_),
    .A2(_0746_),
    .A3(_3389_),
    .ZN(_0747_));
 BUF_X2 _5418_ (.A(_3393_),
    .Z(_0748_));
 AOI21_X2 _5419_ (.A(_0747_),
    .B1(_0748_),
    .B2(_0746_),
    .ZN(_0749_));
 BUF_X2 _5420_ (.A(_3390_),
    .Z(_0750_));
 NAND3_X1 _5421_ (.A1(_0745_),
    .A2(_0746_),
    .A3(_0750_),
    .ZN(_0751_));
 INV_X1 _5422_ (.A(_3321_),
    .ZN(_0752_));
 AOI21_X2 _5423_ (.A(_3325_),
    .B1(_0555_),
    .B2(_3326_),
    .ZN(_0753_));
 OAI21_X1 _5424_ (.A(_0752_),
    .B1(_0753_),
    .B2(_0550_),
    .ZN(_0754_));
 NOR3_X1 _5425_ (.A1(_0332_),
    .A2(_0330_),
    .A3(_0754_),
    .ZN(_0755_));
 OAI21_X1 _5426_ (.A(_0755_),
    .B1(_0451_),
    .B2(_0452_),
    .ZN(_0756_));
 NAND3_X1 _5427_ (.A1(_0329_),
    .A2(_3322_),
    .A3(_3326_),
    .ZN(_0757_));
 NOR2_X1 _5428_ (.A1(_3180_),
    .A2(_0330_),
    .ZN(_0758_));
 OAI221_X2 _5429_ (.A(_0752_),
    .B1(_0757_),
    .B2(_0758_),
    .C1(_0753_),
    .C2(_0550_),
    .ZN(_0759_));
 NAND2_X2 _5430_ (.A1(_0756_),
    .A2(_0759_),
    .ZN(_0760_));
 OAI211_X2 _5431_ (.A(_0744_),
    .B(_0749_),
    .C1(_0751_),
    .C2(_0760_),
    .ZN(_0761_));
 AOI21_X1 _5432_ (.A(_3381_),
    .B1(_0761_),
    .B2(_3382_),
    .ZN(_0762_));
 XOR2_X2 _5433_ (.A(_3378_),
    .B(_0762_),
    .Z(_0763_));
 INV_X1 _5434_ (.A(_0763_),
    .ZN(_3574_));
 NOR4_X2 _5435_ (.A1(_0750_),
    .A2(_3385_),
    .A3(_3389_),
    .A4(_0748_),
    .ZN(_0764_));
 OAI21_X1 _5436_ (.A(_0746_),
    .B1(_0748_),
    .B2(_0745_),
    .ZN(_0765_));
 AOI21_X2 _5437_ (.A(_0764_),
    .B1(_0765_),
    .B2(_0744_),
    .ZN(_0766_));
 OR4_X1 _5438_ (.A1(_3321_),
    .A2(_3385_),
    .A3(_3389_),
    .A4(_0748_),
    .ZN(_0767_));
 NAND2_X1 _5439_ (.A1(_0553_),
    .A2(_0559_),
    .ZN(_0768_));
 OAI21_X1 _5440_ (.A(_0766_),
    .B1(_0767_),
    .B2(_0768_),
    .ZN(_0769_));
 XNOR2_X2 _5441_ (.A(_3382_),
    .B(_0769_),
    .ZN(_3582_));
 OR3_X1 _5442_ (.A1(_0746_),
    .A2(_3389_),
    .A3(_0748_),
    .ZN(_0770_));
 AND3_X1 _5443_ (.A1(_0750_),
    .A2(_0756_),
    .A3(_0759_),
    .ZN(_0771_));
 OAI221_X1 _5444_ (.A(_0749_),
    .B1(_0770_),
    .B2(_0771_),
    .C1(_0751_),
    .C2(_0760_),
    .ZN(_0772_));
 NOR3_X1 _5445_ (.A1(_0745_),
    .A2(_0746_),
    .A3(_0748_),
    .ZN(_0773_));
 OR2_X1 _5446_ (.A1(_0772_),
    .A2(_0773_),
    .ZN(_0774_));
 INV_X1 _5447_ (.A(_0774_),
    .ZN(_3578_));
 NAND3_X1 _5448_ (.A1(_0752_),
    .A2(_0553_),
    .A3(_0559_),
    .ZN(_0775_));
 AOI21_X2 _5449_ (.A(_3389_),
    .B1(_0775_),
    .B2(_0750_),
    .ZN(_0776_));
 XNOR2_X2 _5450_ (.A(_0745_),
    .B(_0776_),
    .ZN(_3546_));
 XNOR2_X2 _5451_ (.A(_0750_),
    .B(_0760_),
    .ZN(_3550_));
 BUF_X2 _5452_ (.A(_3398_),
    .Z(_0777_));
 INV_X1 _5453_ (.A(_3345_),
    .ZN(_0778_));
 OAI21_X2 _5454_ (.A(_3346_),
    .B1(_0608_),
    .B2(_0605_),
    .ZN(_0779_));
 AOI211_X2 _5455_ (.A(_0605_),
    .B(_0607_),
    .C1(_0613_),
    .C2(_0427_),
    .ZN(_0780_));
 OAI21_X1 _5456_ (.A(_0778_),
    .B1(_0779_),
    .B2(_0780_),
    .ZN(_0781_));
 XNOR2_X2 _5457_ (.A(_0777_),
    .B(_0781_),
    .ZN(_0782_));
 INV_X1 _5458_ (.A(_0782_),
    .ZN(_3399_));
 INV_X1 _5459_ (.A(_3409_),
    .ZN(_0783_));
 CLKBUF_X2 _5460_ (.A(_3410_),
    .Z(_0784_));
 BUF_X1 _5461_ (.A(_3414_),
    .Z(_0785_));
 BUF_X1 _5462_ (.A(_3417_),
    .Z(_0786_));
 AND3_X1 _5463_ (.A1(_0784_),
    .A2(_0785_),
    .A3(_0786_),
    .ZN(_0787_));
 CLKBUF_X2 _5464_ (.A(_3418_),
    .Z(_0788_));
 AND3_X1 _5465_ (.A1(_0784_),
    .A2(_0785_),
    .A3(_0788_),
    .ZN(_0789_));
 BUF_X2 _5466_ (.A(_3422_),
    .Z(_0790_));
 AOI21_X2 _5467_ (.A(_3421_),
    .B1(_3425_),
    .B2(_0790_),
    .ZN(_0791_));
 BUF_X2 _5468_ (.A(_3426_),
    .Z(_0792_));
 NAND3_X1 _5469_ (.A1(_0790_),
    .A2(_0792_),
    .A3(_3430_),
    .ZN(_0793_));
 AOI21_X2 _5470_ (.A(_3297_),
    .B1(_0523_),
    .B2(_3298_),
    .ZN(_0794_));
 INV_X1 _5471_ (.A(_3429_),
    .ZN(_0795_));
 NAND2_X2 _5472_ (.A1(_0790_),
    .A2(_0792_),
    .ZN(_0796_));
 OAI221_X2 _5473_ (.A(_0791_),
    .B1(_0793_),
    .B2(_0794_),
    .C1(_0795_),
    .C2(_0796_),
    .ZN(_0797_));
 AOI221_X2 _5474_ (.A(_0787_),
    .B1(_0789_),
    .B2(_0797_),
    .C1(_0784_),
    .C2(_3413_),
    .ZN(_0798_));
 NAND2_X1 _5475_ (.A1(_0783_),
    .A2(_0798_),
    .ZN(_0799_));
 AOI21_X2 _5476_ (.A(_3405_),
    .B1(_0799_),
    .B2(_3406_),
    .ZN(_0800_));
 XOR2_X2 _5477_ (.A(_3402_),
    .B(_0800_),
    .Z(_0801_));
 INV_X1 _5478_ (.A(_0801_),
    .ZN(_3590_));
 INV_X1 _5479_ (.A(_3297_),
    .ZN(_0802_));
 NAND3_X1 _5480_ (.A1(_0520_),
    .A2(_0802_),
    .A3(_0795_),
    .ZN(_0803_));
 AOI21_X2 _5481_ (.A(_0803_),
    .B1(_0246_),
    .B2(_0242_),
    .ZN(_0804_));
 INV_X1 _5482_ (.A(_3298_),
    .ZN(_0805_));
 NAND2_X1 _5483_ (.A1(_0805_),
    .A2(_0802_),
    .ZN(_0806_));
 AOI21_X2 _5484_ (.A(_3429_),
    .B1(_0806_),
    .B2(_3430_),
    .ZN(_0807_));
 NOR3_X4 _5485_ (.A1(_0796_),
    .A2(_0804_),
    .A3(_0807_),
    .ZN(_0808_));
 INV_X1 _5486_ (.A(_0791_),
    .ZN(_0809_));
 OR3_X1 _5487_ (.A1(_3413_),
    .A2(_0786_),
    .A3(_0809_),
    .ZN(_0810_));
 OAI21_X1 _5488_ (.A(_0785_),
    .B1(_0788_),
    .B2(_0786_),
    .ZN(_0811_));
 INV_X1 _5489_ (.A(_0811_),
    .ZN(_0812_));
 OAI221_X2 _5490_ (.A(_0784_),
    .B1(_0808_),
    .B2(_0810_),
    .C1(_0812_),
    .C2(_3413_),
    .ZN(_0813_));
 NAND2_X1 _5491_ (.A1(_0783_),
    .A2(_0813_),
    .ZN(_0814_));
 XNOR2_X1 _5492_ (.A(_3406_),
    .B(_0814_),
    .ZN(_0815_));
 INV_X1 _5493_ (.A(_0815_),
    .ZN(_3620_));
 NOR2_X1 _5494_ (.A1(_0784_),
    .A2(_3413_),
    .ZN(_0816_));
 AOI21_X1 _5495_ (.A(_0786_),
    .B1(_0797_),
    .B2(_0788_),
    .ZN(_0817_));
 INV_X1 _5496_ (.A(_0785_),
    .ZN(_0818_));
 OAI21_X1 _5497_ (.A(_0816_),
    .B1(_0817_),
    .B2(_0818_),
    .ZN(_0819_));
 NAND2_X1 _5498_ (.A1(_0798_),
    .A2(_0819_),
    .ZN(_0820_));
 INV_X1 _5499_ (.A(_0820_),
    .ZN(_3596_));
 OR3_X2 _5500_ (.A1(_0786_),
    .A2(_0809_),
    .A3(_0808_),
    .ZN(_0821_));
 NOR2_X1 _5501_ (.A1(_0785_),
    .A2(_0786_),
    .ZN(_0822_));
 OAI21_X2 _5502_ (.A(_0788_),
    .B1(_0809_),
    .B2(_0808_),
    .ZN(_0823_));
 AOI22_X4 _5503_ (.A1(_0812_),
    .A2(_0821_),
    .B1(_0822_),
    .B2(_0823_),
    .ZN(_3600_));
 XNOR2_X1 _5504_ (.A(_0788_),
    .B(_0797_),
    .ZN(_0824_));
 INV_X2 _5505_ (.A(_0824_),
    .ZN(_3604_));
 INV_X1 _5506_ (.A(_3464_),
    .ZN(_3154_));
 INV_X1 _5507_ (.A(_3463_),
    .ZN(_3299_));
 NOR2_X2 _5508_ (.A1(_3154_),
    .A2(_3299_),
    .ZN(_0825_));
 NOR2_X1 _5509_ (.A1(_0804_),
    .A2(_0807_),
    .ZN(_0826_));
 AOI21_X2 _5510_ (.A(_3425_),
    .B1(_0826_),
    .B2(_0792_),
    .ZN(_0827_));
 XNOR2_X2 _5511_ (.A(_0790_),
    .B(_0827_),
    .ZN(_3608_));
 INV_X1 _5512_ (.A(_3430_),
    .ZN(_0828_));
 OAI21_X1 _5513_ (.A(_0795_),
    .B1(_0794_),
    .B2(_0828_),
    .ZN(_0829_));
 XOR2_X2 _5514_ (.A(_0792_),
    .B(_0829_),
    .Z(_3612_));
 AOI21_X1 _5515_ (.A(_3140_),
    .B1(_0246_),
    .B2(_0242_),
    .ZN(_0830_));
 OAI21_X1 _5516_ (.A(_0802_),
    .B1(_0830_),
    .B2(_0805_),
    .ZN(_0831_));
 XNOR2_X2 _5517_ (.A(_0828_),
    .B(_0831_),
    .ZN(_3514_));
 OR2_X1 _5518_ (.A1(_3612_),
    .A2(_3514_),
    .ZN(_0832_));
 NOR4_X2 _5519_ (.A1(_3600_),
    .A2(_3604_),
    .A3(_3608_),
    .A4(_0832_),
    .ZN(_0833_));
 AND3_X1 _5520_ (.A1(_0815_),
    .A2(_0820_),
    .A3(_0833_),
    .ZN(_0834_));
 AOI21_X1 _5521_ (.A(_3483_),
    .B1(_0825_),
    .B2(_0834_),
    .ZN(_0835_));
 XNOR2_X1 _5522_ (.A(_3590_),
    .B(_0835_),
    .ZN(_3431_));
 BUF_X16 _5523_ (.A(_0517_),
    .Z(_3470_));
 BUF_X2 _5524_ (.A(_3465_),
    .Z(_0836_));
 NAND3_X1 _5525_ (.A1(_0836_),
    .A2(_0820_),
    .A3(_0833_),
    .ZN(_0837_));
 AND2_X1 _5526_ (.A1(net9),
    .A2(_0837_),
    .ZN(_0838_));
 XNOR2_X1 _5527_ (.A(_3620_),
    .B(_0838_),
    .ZN(_3435_));
 AOI21_X1 _5528_ (.A(_3483_),
    .B1(_0825_),
    .B2(_0833_),
    .ZN(_0839_));
 XNOR2_X1 _5529_ (.A(_3596_),
    .B(_0839_),
    .ZN(_3439_));
 NOR3_X1 _5530_ (.A1(_3604_),
    .A2(_3608_),
    .A3(_0832_),
    .ZN(_0840_));
 AOI21_X1 _5531_ (.A(_3483_),
    .B1(_0840_),
    .B2(_0836_),
    .ZN(_0841_));
 XNOR2_X1 _5532_ (.A(_3600_),
    .B(_0841_),
    .ZN(_3443_));
 NOR2_X1 _5533_ (.A1(_3608_),
    .A2(_0832_),
    .ZN(_0842_));
 AOI21_X1 _5534_ (.A(_0519_),
    .B1(_0825_),
    .B2(_0842_),
    .ZN(_0843_));
 XNOR2_X1 _5535_ (.A(_3604_),
    .B(_0843_),
    .ZN(_3447_));
 NOR2_X1 _5536_ (.A1(_3612_),
    .A2(_3514_),
    .ZN(_0844_));
 AOI21_X1 _5537_ (.A(_0519_),
    .B1(_0844_),
    .B2(_0836_),
    .ZN(_0845_));
 XNOR2_X1 _5538_ (.A(_3608_),
    .B(_0845_),
    .ZN(_3451_));
 INV_X1 _5539_ (.A(_3514_),
    .ZN(_0846_));
 AOI21_X1 _5540_ (.A(_0519_),
    .B1(_0825_),
    .B2(_0846_),
    .ZN(_0847_));
 XNOR2_X1 _5541_ (.A(_3612_),
    .B(_0847_),
    .ZN(_3455_));
 NOR2_X1 _5542_ (.A1(_0836_),
    .A2(_3483_),
    .ZN(_0848_));
 XNOR2_X1 _5543_ (.A(_3514_),
    .B(_0848_),
    .ZN(_3459_));
 NOR2_X1 _5544_ (.A1(net218),
    .A2(_3463_),
    .ZN(_0849_));
 AOI21_X2 _5545_ (.A(_0849_),
    .B1(net9),
    .B2(_3466_),
    .ZN(_2950_));
 INV_X1 _5546_ (.A(_3441_),
    .ZN(_0850_));
 INV_X1 _5547_ (.A(_3449_),
    .ZN(_0851_));
 INV_X1 _5548_ (.A(_3457_),
    .ZN(_0852_));
 INV_X1 _5549_ (.A(_3467_),
    .ZN(_0853_));
 INV_X1 _5550_ (.A(_3468_),
    .ZN(_0854_));
 OAI21_X1 _5551_ (.A(_0853_),
    .B1(_0854_),
    .B2(_3155_),
    .ZN(_0855_));
 BUF_X1 _5552_ (.A(_3462_),
    .Z(_0856_));
 AOI21_X1 _5553_ (.A(_3461_),
    .B1(_0855_),
    .B2(_0856_),
    .ZN(_0857_));
 INV_X1 _5554_ (.A(_3458_),
    .ZN(_0858_));
 OAI21_X1 _5555_ (.A(_0852_),
    .B1(_0857_),
    .B2(_0858_),
    .ZN(_0859_));
 AOI21_X2 _5556_ (.A(_3453_),
    .B1(_0859_),
    .B2(_3454_),
    .ZN(_0860_));
 INV_X1 _5557_ (.A(_3450_),
    .ZN(_0861_));
 OAI21_X1 _5558_ (.A(_0851_),
    .B1(_0860_),
    .B2(_0861_),
    .ZN(_0862_));
 CLKBUF_X2 _5559_ (.A(_3446_),
    .Z(_0863_));
 AOI21_X2 _5560_ (.A(_3445_),
    .B1(_0862_),
    .B2(_0863_),
    .ZN(_0864_));
 INV_X1 _5561_ (.A(_3442_),
    .ZN(_0865_));
 OAI21_X1 _5562_ (.A(_0850_),
    .B1(_0864_),
    .B2(_0865_),
    .ZN(_0866_));
 BUF_X2 _5563_ (.A(_3438_),
    .Z(_0867_));
 AOI21_X2 _5564_ (.A(_3437_),
    .B1(_0866_),
    .B2(_0867_),
    .ZN(_0868_));
 XNOR2_X2 _5565_ (.A(_3434_),
    .B(_0868_),
    .ZN(_3666_));
 XNOR2_X2 _5566_ (.A(_3450_),
    .B(_0860_),
    .ZN(_3644_));
 INV_X1 _5567_ (.A(_3644_),
    .ZN(_3533_));
 INV_X1 _5568_ (.A(_3454_),
    .ZN(_0869_));
 AOI21_X1 _5569_ (.A(_3461_),
    .B1(_0856_),
    .B2(_2952_),
    .ZN(_0870_));
 OAI21_X2 _5570_ (.A(_0852_),
    .B1(_0870_),
    .B2(_0858_),
    .ZN(_0871_));
 XNOR2_X2 _5571_ (.A(_0869_),
    .B(_0871_),
    .ZN(_3648_));
 INV_X1 _5572_ (.A(_3648_),
    .ZN(_3532_));
 INV_X1 _5573_ (.A(_3471_),
    .ZN(_0872_));
 AND3_X1 _5574_ (.A1(_3472_),
    .A2(_3475_),
    .A3(_3477_),
    .ZN(_0873_));
 AOI21_X2 _5575_ (.A(_0873_),
    .B1(_3474_),
    .B2(_3472_),
    .ZN(_0874_));
 NAND3_X2 _5576_ (.A1(_3472_),
    .A2(_3475_),
    .A3(_3478_),
    .ZN(_0875_));
 INV_X1 _5577_ (.A(_3484_),
    .ZN(_0876_));
 BUF_X1 _5578_ (.A(_3491_),
    .Z(_0877_));
 AOI21_X1 _5579_ (.A(_3490_),
    .B1(_3493_),
    .B2(_0877_),
    .ZN(_0878_));
 NAND2_X1 _5580_ (.A1(_0877_),
    .A2(_3494_),
    .ZN(_0879_));
 INV_X1 _5581_ (.A(_3499_),
    .ZN(_0880_));
 INV_X1 _5582_ (.A(_3505_),
    .ZN(_0881_));
 INV_X1 _5583_ (.A(_3511_),
    .ZN(_0882_));
 INV_X2 _5584_ (.A(_3512_),
    .ZN(_0883_));
 OAI21_X4 _5585_ (.A(_0882_),
    .B1(_0883_),
    .B2(_0005_),
    .ZN(_0884_));
 AOI21_X4 _5586_ (.A(_3508_),
    .B1(_0884_),
    .B2(_3509_),
    .ZN(_0885_));
 BUF_X1 _5587_ (.A(_3506_),
    .Z(_0886_));
 INV_X1 _5588_ (.A(_0886_),
    .ZN(_0887_));
 OAI21_X4 _5589_ (.A(_0881_),
    .B1(_0885_),
    .B2(_0887_),
    .ZN(_0888_));
 AOI21_X4 _5590_ (.A(_3502_),
    .B1(_3503_),
    .B2(_0888_),
    .ZN(_0889_));
 BUF_X1 _5591_ (.A(_3500_),
    .Z(_0890_));
 INV_X1 _5592_ (.A(_0890_),
    .ZN(_0891_));
 OAI21_X4 _5593_ (.A(_0880_),
    .B1(_0889_),
    .B2(_0891_),
    .ZN(_0892_));
 AOI21_X4 _5594_ (.A(_3496_),
    .B1(_0892_),
    .B2(_3497_),
    .ZN(_0893_));
 OAI21_X4 _5595_ (.A(_0878_),
    .B1(_0893_),
    .B2(_0879_),
    .ZN(_0894_));
 AOI21_X4 _5596_ (.A(_3487_),
    .B1(_0894_),
    .B2(_3488_),
    .ZN(_0895_));
 INV_X1 _5597_ (.A(_3485_),
    .ZN(_0896_));
 OAI21_X4 _5598_ (.A(_0876_),
    .B1(_0895_),
    .B2(_0896_),
    .ZN(_0897_));
 AOI21_X4 _5599_ (.A(_3480_),
    .B1(_0897_),
    .B2(_3481_),
    .ZN(_0898_));
 OAI211_X4 _5600_ (.A(_0872_),
    .B(_0874_),
    .C1(_0898_),
    .C2(_0875_),
    .ZN(_0899_));
 INV_X8 _5601_ (.A(_0899_),
    .ZN(_0900_));
 BUF_X16 _5602_ (.A(_0900_),
    .Z(_0901_));
 BUF_X32 _5603_ (.A(_0901_),
    .Z(_3686_));
 INV_X1 _5604_ (.A(_0635_),
    .ZN(_0902_));
 OAI21_X2 _5605_ (.A(_0625_),
    .B1(_0480_),
    .B2(_0632_),
    .ZN(_0903_));
 AOI21_X4 _5606_ (.A(_3223_),
    .B1(_0902_),
    .B2(_0903_),
    .ZN(_0904_));
 XOR2_X2 _5607_ (.A(_3358_),
    .B(_0904_),
    .Z(_0905_));
 INV_X1 _5608_ (.A(_0905_),
    .ZN(_3436_));
 INV_X1 _5609_ (.A(_3301_),
    .ZN(_0906_));
 INV_X1 _5610_ (.A(_3308_),
    .ZN(_0907_));
 AOI21_X1 _5611_ (.A(_3314_),
    .B1(_3315_),
    .B2(_2945_),
    .ZN(_0908_));
 INV_X1 _5612_ (.A(_3309_),
    .ZN(_0909_));
 OAI21_X1 _5613_ (.A(_0907_),
    .B1(_0908_),
    .B2(_0909_),
    .ZN(_0910_));
 AOI21_X1 _5614_ (.A(_3304_),
    .B1(_0910_),
    .B2(_3305_),
    .ZN(_0911_));
 INV_X1 _5615_ (.A(_3302_),
    .ZN(_0912_));
 OAI21_X2 _5616_ (.A(_0906_),
    .B1(_0911_),
    .B2(_0912_),
    .ZN(_0913_));
 XNOR2_X2 _5617_ (.A(_3516_),
    .B(_0913_),
    .ZN(_3659_));
 AOI21_X1 _5618_ (.A(_3453_),
    .B1(_0871_),
    .B2(_3454_),
    .ZN(_0914_));
 OAI21_X2 _5619_ (.A(_0851_),
    .B1(_0914_),
    .B2(_0861_),
    .ZN(_0915_));
 XNOR2_X2 _5620_ (.A(_0863_),
    .B(_0915_),
    .ZN(_0916_));
 INV_X1 _5621_ (.A(_0916_),
    .ZN(_3640_));
 XNOR2_X2 _5622_ (.A(_0865_),
    .B(_0864_),
    .ZN(_0917_));
 INV_X1 _5623_ (.A(_0917_),
    .ZN(_3636_));
 INV_X1 _5624_ (.A(_3522_),
    .ZN(_0918_));
 INV_X1 _5625_ (.A(_3530_),
    .ZN(_0919_));
 AOI21_X1 _5626_ (.A(_3536_),
    .B1(_3537_),
    .B2(_2954_),
    .ZN(_0920_));
 INV_X1 _5627_ (.A(_3531_),
    .ZN(_0921_));
 OAI21_X1 _5628_ (.A(_0919_),
    .B1(_0920_),
    .B2(_0921_),
    .ZN(_0922_));
 AOI21_X1 _5629_ (.A(_3526_),
    .B1(_0922_),
    .B2(_3527_),
    .ZN(_0923_));
 INV_X1 _5630_ (.A(_3523_),
    .ZN(_0924_));
 OAI21_X2 _5631_ (.A(_0918_),
    .B1(_0923_),
    .B2(_0924_),
    .ZN(_0925_));
 XNOR2_X2 _5632_ (.A(_3520_),
    .B(_0925_),
    .ZN(_3842_));
 BUF_X4 _5633_ (.A(_3544_),
    .Z(_0926_));
 INV_X1 _5634_ (.A(_3397_),
    .ZN(_0927_));
 NOR3_X1 _5635_ (.A1(_3200_),
    .A2(_3199_),
    .A3(_0605_),
    .ZN(_0928_));
 AOI211_X2 _5636_ (.A(_3199_),
    .B(_3203_),
    .C1(_3207_),
    .C2(_0406_),
    .ZN(_0929_));
 INV_X1 _5637_ (.A(_0605_),
    .ZN(_0930_));
 AOI211_X2 _5638_ (.A(_0779_),
    .B(_0928_),
    .C1(_0929_),
    .C2(_0930_),
    .ZN(_0931_));
 OAI21_X1 _5639_ (.A(_0777_),
    .B1(_3345_),
    .B2(_0931_),
    .ZN(_0932_));
 NOR2_X1 _5640_ (.A1(_0612_),
    .A2(_0779_),
    .ZN(_0933_));
 NAND4_X1 _5641_ (.A1(_0777_),
    .A2(_0411_),
    .A3(_0417_),
    .A4(_0933_),
    .ZN(_0934_));
 AND3_X1 _5642_ (.A1(_0927_),
    .A2(_0932_),
    .A3(_0934_),
    .ZN(_0935_));
 XNOR2_X2 _5643_ (.A(_0926_),
    .B(_0935_),
    .ZN(_3562_));
 INV_X1 _5644_ (.A(_3562_),
    .ZN(_0936_));
 BUF_X16 _5645_ (.A(_0435_),
    .Z(_2942_));
 NOR4_X4 _5646_ (.A1(_3412_),
    .A2(_3416_),
    .A3(_3404_),
    .A4(_3408_),
    .ZN(_0937_));
 NAND3_X1 _5647_ (.A1(_0444_),
    .A2(_0782_),
    .A3(_0937_),
    .ZN(_0938_));
 NAND2_X1 _5648_ (.A1(net224),
    .A2(_0938_),
    .ZN(_0939_));
 XNOR2_X1 _5649_ (.A(_0936_),
    .B(_0939_),
    .ZN(_3545_));
 INV_X1 _5650_ (.A(_0937_),
    .ZN(_0940_));
 NOR2_X1 _5651_ (.A1(_0460_),
    .A2(_0940_),
    .ZN(_0941_));
 NOR2_X1 _5652_ (.A1(net17),
    .A2(_0941_),
    .ZN(_0942_));
 XNOR2_X1 _5653_ (.A(_3399_),
    .B(_0942_),
    .ZN(_3549_));
 BUF_X2 _5654_ (.A(_3552_),
    .Z(_0943_));
 NAND4_X2 _5655_ (.A1(_0624_),
    .A2(_0943_),
    .A3(_0633_),
    .A4(_0636_),
    .ZN(_0944_));
 AOI21_X2 _5656_ (.A(_3551_),
    .B1(_3353_),
    .B2(_0943_),
    .ZN(_0945_));
 NAND2_X1 _5657_ (.A1(_0944_),
    .A2(_0945_),
    .ZN(_0946_));
 XNOR2_X2 _5658_ (.A(_3548_),
    .B(_0946_),
    .ZN(_0947_));
 INV_X1 _5659_ (.A(_0947_),
    .ZN(_3566_));
 OR3_X1 _5660_ (.A1(_3345_),
    .A2(_3397_),
    .A3(_3543_),
    .ZN(_0948_));
 NOR2_X1 _5661_ (.A1(_0931_),
    .A2(_0948_),
    .ZN(_0949_));
 NOR3_X1 _5662_ (.A1(_0777_),
    .A2(_3397_),
    .A3(_3543_),
    .ZN(_0950_));
 NOR2_X1 _5663_ (.A1(_0926_),
    .A2(_3543_),
    .ZN(_0951_));
 NAND3_X1 _5664_ (.A1(_0777_),
    .A2(_0926_),
    .A3(_0933_),
    .ZN(_0952_));
 INV_X1 _5665_ (.A(_0413_),
    .ZN(_0953_));
 INV_X1 _5666_ (.A(_0424_),
    .ZN(_0954_));
 INV_X1 _5667_ (.A(_0425_),
    .ZN(_0955_));
 AOI221_X2 _5668_ (.A(_0953_),
    .B1(_0454_),
    .B2(_0954_),
    .C1(_0955_),
    .C2(_0414_),
    .ZN(_0956_));
 OAI33_X1 _5669_ (.A1(_0949_),
    .A2(_0950_),
    .A3(_0951_),
    .B1(_0952_),
    .B2(_0412_),
    .B3(_0956_),
    .ZN(_0957_));
 XOR2_X2 _5670_ (.A(_3556_),
    .B(_0957_),
    .Z(_3557_));
 INV_X1 _5671_ (.A(_3560_),
    .ZN(_0958_));
 INV_X1 _5672_ (.A(_3563_),
    .ZN(_0959_));
 OAI21_X2 _5673_ (.A(_3402_),
    .B1(_3406_),
    .B2(_3405_),
    .ZN(_0960_));
 NOR2_X1 _5674_ (.A1(_3405_),
    .A2(_3409_),
    .ZN(_0961_));
 AOI21_X1 _5675_ (.A(_0960_),
    .B1(_0961_),
    .B2(_0798_),
    .ZN(_0962_));
 OAI21_X1 _5676_ (.A(_3564_),
    .B1(_3401_),
    .B2(_0962_),
    .ZN(_0963_));
 AND2_X1 _5677_ (.A1(_0959_),
    .A2(_0963_),
    .ZN(_0964_));
 XNOR2_X2 _5678_ (.A(_0958_),
    .B(_0964_),
    .ZN(_0965_));
 INV_X1 _5679_ (.A(_0965_),
    .ZN(_3586_));
 AOI21_X2 _5680_ (.A(_0960_),
    .B1(_0813_),
    .B2(_0961_),
    .ZN(_0966_));
 NOR2_X1 _5681_ (.A1(_3401_),
    .A2(_0966_),
    .ZN(_0967_));
 XOR2_X2 _5682_ (.A(_3564_),
    .B(_0967_),
    .Z(_0968_));
 INV_X1 _5683_ (.A(_0968_),
    .ZN(_3616_));
 AND4_X2 _5684_ (.A1(_0801_),
    .A2(_0825_),
    .A3(_0834_),
    .A4(_0968_),
    .ZN(_0969_));
 NOR2_X1 _5685_ (.A1(_3483_),
    .A2(_0969_),
    .ZN(_0970_));
 XNOR2_X1 _5686_ (.A(_3586_),
    .B(_0970_),
    .ZN(_3565_));
 INV_X1 _5687_ (.A(_3353_),
    .ZN(_0971_));
 NAND2_X1 _5688_ (.A1(_0624_),
    .A2(_3358_),
    .ZN(_0972_));
 INV_X1 _5689_ (.A(_3357_),
    .ZN(_0973_));
 INV_X1 _5690_ (.A(_0624_),
    .ZN(_0974_));
 OAI221_X2 _5691_ (.A(_0971_),
    .B1(_0904_),
    .B2(_0972_),
    .C1(_0973_),
    .C2(_0974_),
    .ZN(_0975_));
 XOR2_X2 _5692_ (.A(_0943_),
    .B(_0975_),
    .Z(_3570_));
 AND2_X1 _5693_ (.A1(_0801_),
    .A2(_0834_),
    .ZN(_0976_));
 AOI21_X1 _5694_ (.A(_0519_),
    .B1(_0976_),
    .B2(_0836_),
    .ZN(_0977_));
 XNOR2_X1 _5695_ (.A(_3616_),
    .B(_0977_),
    .ZN(_3569_));
 BUF_X1 _5696_ (.A(_3571_),
    .Z(_0978_));
 INV_X1 _5697_ (.A(_3572_),
    .ZN(_0979_));
 NAND3_X1 _5698_ (.A1(_0867_),
    .A2(_3434_),
    .A3(_3441_),
    .ZN(_0980_));
 INV_X1 _5699_ (.A(_3437_),
    .ZN(_0981_));
 INV_X1 _5700_ (.A(_3434_),
    .ZN(_0982_));
 OAI21_X2 _5701_ (.A(_0980_),
    .B1(_0981_),
    .B2(_0982_),
    .ZN(_0983_));
 AND3_X1 _5702_ (.A1(_3442_),
    .A2(_0867_),
    .A3(_3434_),
    .ZN(_0984_));
 INV_X1 _5703_ (.A(_3445_),
    .ZN(_0985_));
 INV_X1 _5704_ (.A(_3453_),
    .ZN(_0986_));
 INV_X1 _5705_ (.A(_3461_),
    .ZN(_0987_));
 INV_X1 _5706_ (.A(_3155_),
    .ZN(_2949_));
 AOI21_X1 _5707_ (.A(_3467_),
    .B1(_3468_),
    .B2(_2949_),
    .ZN(_0988_));
 INV_X1 _5708_ (.A(_0856_),
    .ZN(_0989_));
 OAI21_X1 _5709_ (.A(_0987_),
    .B1(_0988_),
    .B2(_0989_),
    .ZN(_0990_));
 AOI21_X1 _5710_ (.A(_3457_),
    .B1(_0990_),
    .B2(_3458_),
    .ZN(_0991_));
 OAI21_X1 _5711_ (.A(_0986_),
    .B1(_0991_),
    .B2(_0869_),
    .ZN(_0992_));
 AOI21_X1 _5712_ (.A(_3449_),
    .B1(_0992_),
    .B2(_3450_),
    .ZN(_0993_));
 INV_X1 _5713_ (.A(_0863_),
    .ZN(_0994_));
 OAI21_X2 _5714_ (.A(_0985_),
    .B1(_0993_),
    .B2(_0994_),
    .ZN(_0995_));
 AOI211_X2 _5715_ (.A(_3433_),
    .B(_0983_),
    .C1(_0984_),
    .C2(_0995_),
    .ZN(_0996_));
 NOR2_X1 _5716_ (.A1(_0979_),
    .A2(_0996_),
    .ZN(_0997_));
 NOR2_X1 _5717_ (.A1(_0978_),
    .A2(_0997_),
    .ZN(_0998_));
 XNOR2_X2 _5718_ (.A(_3568_),
    .B(_0998_),
    .ZN(_3624_));
 NAND3_X1 _5719_ (.A1(_0782_),
    .A2(_0936_),
    .A3(_0941_),
    .ZN(_0999_));
 OAI21_X1 _5720_ (.A(net224),
    .B1(_3557_),
    .B2(_0999_),
    .ZN(_1000_));
 INV_X1 _5721_ (.A(_3555_),
    .ZN(_1001_));
 NOR2_X1 _5722_ (.A1(_0950_),
    .A2(_0951_),
    .ZN(_1002_));
 OAI211_X2 _5723_ (.A(_3556_),
    .B(_1002_),
    .C1(_0948_),
    .C2(_0931_),
    .ZN(_1003_));
 NAND2_X1 _5724_ (.A1(_0413_),
    .A2(_0416_),
    .ZN(_1004_));
 NAND2_X1 _5725_ (.A1(_0777_),
    .A2(_0926_),
    .ZN(_1005_));
 OAI21_X2 _5726_ (.A(_3556_),
    .B1(_3211_),
    .B2(_3212_),
    .ZN(_1006_));
 NOR4_X4 _5727_ (.A1(_1006_),
    .A2(_0779_),
    .A3(_0612_),
    .A4(_1005_),
    .ZN(_1007_));
 NAND3_X2 _5728_ (.A1(_0411_),
    .A2(_1007_),
    .A3(_1004_),
    .ZN(_1008_));
 AND3_X4 _5729_ (.A1(_1008_),
    .A2(_1003_),
    .A3(_1001_),
    .ZN(_1009_));
 NOR4_X4 _5730_ (.A1(_1009_),
    .A2(_0704_),
    .A3(_0711_),
    .A4(_0699_),
    .ZN(_1010_));
 NAND3_X4 _5731_ (.A1(_1008_),
    .A2(_1003_),
    .A3(_1001_),
    .ZN(_1011_));
 NAND2_X1 _5732_ (.A1(_0699_),
    .A2(_1011_),
    .ZN(_1012_));
 AND3_X1 _5733_ (.A1(_0581_),
    .A2(_0586_),
    .A3(_0709_),
    .ZN(_1013_));
 OAI221_X2 _5734_ (.A(_0019_),
    .B1(_1013_),
    .B2(_0707_),
    .C1(_3365_),
    .C2(_0659_),
    .ZN(_1014_));
 NOR3_X1 _5735_ (.A1(_3363_),
    .A2(_0018_),
    .A3(_0701_),
    .ZN(_1015_));
 NAND4_X1 _5736_ (.A1(_0571_),
    .A2(_0564_),
    .A3(_0641_),
    .A4(_0639_),
    .ZN(_1016_));
 OAI21_X1 _5737_ (.A(_1015_),
    .B1(_1016_),
    .B2(_0728_),
    .ZN(_1017_));
 AOI21_X2 _5738_ (.A(_1012_),
    .B1(_1014_),
    .B2(_1017_),
    .ZN(_1018_));
 XOR2_X2 _5739_ (.A(net13),
    .B(net31),
    .Z(_1019_));
 NAND2_X1 _5740_ (.A1(_1019_),
    .A2(_1009_),
    .ZN(_1020_));
 AOI21_X1 _5741_ (.A(_1020_),
    .B1(_1014_),
    .B2(_1017_),
    .ZN(_1021_));
 NOR4_X2 _5742_ (.A1(_1019_),
    .A2(_0704_),
    .A3(_0711_),
    .A4(_1011_),
    .ZN(_1022_));
 NOR4_X2 _5743_ (.A1(_1021_),
    .A2(_1018_),
    .A3(_1010_),
    .A4(_1022_),
    .ZN(_1023_));
 NOR2_X1 _5744_ (.A1(_0639_),
    .A2(_0652_),
    .ZN(_1024_));
 AND3_X1 _5745_ (.A1(_0344_),
    .A2(_0379_),
    .A3(_1024_),
    .ZN(_1025_));
 AND3_X1 _5746_ (.A1(_0344_),
    .A2(_0380_),
    .A3(_1024_),
    .ZN(_1026_));
 AOI221_X2 _5747_ (.A(_1025_),
    .B1(_1026_),
    .B2(_0270_),
    .C1(_0343_),
    .C2(_1024_),
    .ZN(_1027_));
 OAI21_X1 _5748_ (.A(_0651_),
    .B1(_0653_),
    .B2(_0569_),
    .ZN(_1028_));
 AOI211_X2 _5749_ (.A(_3365_),
    .B(_0017_),
    .C1(_1028_),
    .C2(_0659_),
    .ZN(_1029_));
 NOR2_X1 _5750_ (.A1(_0650_),
    .A2(_0718_),
    .ZN(_1030_));
 NOR4_X2 _5751_ (.A1(_3368_),
    .A2(_3360_),
    .A3(_0590_),
    .A4(_1030_),
    .ZN(_1031_));
 OAI21_X2 _5752_ (.A(_1031_),
    .B1(_0593_),
    .B2(_0260_),
    .ZN(_1032_));
 AOI21_X1 _5753_ (.A(_0650_),
    .B1(_0663_),
    .B2(_0718_),
    .ZN(_1033_));
 OAI21_X1 _5754_ (.A(_0639_),
    .B1(_3368_),
    .B2(_1033_),
    .ZN(_1034_));
 INV_X1 _5755_ (.A(_3360_),
    .ZN(_1035_));
 AOI21_X2 _5756_ (.A(_0014_),
    .B1(_1034_),
    .B2(_1035_),
    .ZN(_1036_));
 AOI22_X4 _5757_ (.A1(_1027_),
    .A2(_1029_),
    .B1(_1032_),
    .B2(_1036_),
    .ZN(_1037_));
 XNOR2_X2 _5758_ (.A(_0699_),
    .B(_1037_),
    .ZN(_1038_));
 NOR2_X1 _5759_ (.A1(_0179_),
    .A2(_1038_),
    .ZN(_1039_));
 XNOR2_X2 _5760_ (.A(_1019_),
    .B(_1037_),
    .ZN(_1040_));
 NOR2_X1 _5761_ (.A1(_0053_),
    .A2(_1040_),
    .ZN(_1041_));
 OAI21_X1 _5762_ (.A(_1023_),
    .B1(_1039_),
    .B2(_1041_),
    .ZN(_1042_));
 OR3_X2 _5763_ (.A1(_1023_),
    .A2(_1039_),
    .A3(_1041_),
    .ZN(_1043_));
 NOR4_X2 _5764_ (.A1(_0323_),
    .A2(_0258_),
    .A3(_0262_),
    .A4(_0095_),
    .ZN(_1044_));
 AND3_X1 _5765_ (.A1(_0014_),
    .A2(_0139_),
    .A3(_0325_),
    .ZN(_1045_));
 INV_X1 _5766_ (.A(_0271_),
    .ZN(_1046_));
 AOI21_X2 _5767_ (.A(_1044_),
    .B1(_1045_),
    .B2(_1046_),
    .ZN(_1047_));
 NAND4_X1 _5768_ (.A1(_0365_),
    .A2(_0377_),
    .A3(_0393_),
    .A4(_0394_),
    .ZN(_1048_));
 OR4_X4 _5769_ (.A1(_3324_),
    .A2(_3392_),
    .A3(_1047_),
    .A4(_1048_),
    .ZN(_1049_));
 XNOR2_X1 _5770_ (.A(_0048_),
    .B(_0037_),
    .ZN(_1050_));
 OR4_X1 _5771_ (.A1(_2906_),
    .A2(_0031_),
    .A3(_0173_),
    .A4(_1050_),
    .ZN(_1051_));
 MUX2_X2 _5772_ (.A(_0166_),
    .B(_1051_),
    .S(_0018_),
    .Z(_1052_));
 OR4_X1 _5773_ (.A1(net213),
    .A2(_3376_),
    .A3(_3380_),
    .A4(_1052_),
    .ZN(_1053_));
 NOR3_X1 _5774_ (.A1(_3384_),
    .A2(_1049_),
    .A3(_1053_),
    .ZN(_1054_));
 OR2_X4 _5775_ (.A1(_3384_),
    .A2(_1049_),
    .ZN(_1055_));
 NOR4_X1 _5776_ (.A1(net213),
    .A2(_3376_),
    .A3(_3380_),
    .A4(_1052_),
    .ZN(_1056_));
 NAND2_X1 _5777_ (.A1(_1023_),
    .A2(_1056_),
    .ZN(_1057_));
 OAI221_X2 _5778_ (.A(_1042_),
    .B1(_1054_),
    .B2(_1043_),
    .C1(_1055_),
    .C2(_1057_),
    .ZN(_1058_));
 BUF_X4 _5779_ (.A(_1058_),
    .Z(_1059_));
 MUX2_X1 _5780_ (.A(_1000_),
    .B(net224),
    .S(_1059_),
    .Z(_3573_));
 NOR2_X1 _5781_ (.A1(_3562_),
    .A2(_3557_),
    .ZN(_1060_));
 NAND4_X4 _5782_ (.A1(_0444_),
    .A2(_0782_),
    .A3(_0937_),
    .A4(_1060_),
    .ZN(_1061_));
 AND2_X1 _5783_ (.A1(_0232_),
    .A2(_0216_),
    .ZN(_1062_));
 OAI221_X2 _5784_ (.A(_1061_),
    .B1(_0212_),
    .B2(_1062_),
    .C1(_3043_),
    .C2(_0210_),
    .ZN(_1063_));
 XOR2_X2 _5785_ (.A(_1059_),
    .B(_1063_),
    .Z(_3581_));
 NAND2_X1 _5786_ (.A1(net18),
    .A2(_0999_),
    .ZN(_1064_));
 XOR2_X2 _5787_ (.A(_3557_),
    .B(_1064_),
    .Z(_3577_));
 BUF_X2 _5788_ (.A(_3580_),
    .Z(_1065_));
 INV_X1 _5789_ (.A(_3584_),
    .ZN(_1066_));
 NOR2_X1 _5790_ (.A1(_3576_),
    .A2(_1066_),
    .ZN(_1067_));
 NAND2_X1 _5791_ (.A1(_1065_),
    .A2(_1067_),
    .ZN(_1068_));
 INV_X2 _5792_ (.A(_3576_),
    .ZN(_1069_));
 CLKBUF_X2 _5793_ (.A(_3579_),
    .Z(_1070_));
 BUF_X1 _5794_ (.A(_3583_),
    .Z(_1071_));
 OR3_X1 _5795_ (.A1(_1069_),
    .A2(_1070_),
    .A3(_1071_),
    .ZN(_1072_));
 NOR3_X1 _5796_ (.A1(_3353_),
    .A2(_3547_),
    .A3(_3551_),
    .ZN(_1073_));
 OAI221_X2 _5797_ (.A(_1073_),
    .B1(_0972_),
    .B2(_0904_),
    .C1(_0974_),
    .C2(_0973_),
    .ZN(_1074_));
 OR2_X1 _5798_ (.A1(_0943_),
    .A2(_3547_),
    .ZN(_1075_));
 OAI221_X2 _5799_ (.A(_1074_),
    .B1(_1075_),
    .B2(_3551_),
    .C1(_3547_),
    .C2(_3548_),
    .ZN(_1076_));
 MUX2_X1 _5800_ (.A(_1068_),
    .B(_1072_),
    .S(_1076_),
    .Z(_1077_));
 NOR4_X1 _5801_ (.A1(_1069_),
    .A2(_1065_),
    .A3(_1070_),
    .A4(_1071_),
    .ZN(_1078_));
 NOR3_X1 _5802_ (.A1(_1069_),
    .A2(_3584_),
    .A3(_1071_),
    .ZN(_1079_));
 OR2_X2 _5803_ (.A1(_1078_),
    .A2(_1079_),
    .ZN(_1080_));
 AOI221_X2 _5804_ (.A(_1080_),
    .B1(_1067_),
    .B2(_1070_),
    .C1(_1069_),
    .C2(_1071_),
    .ZN(_1081_));
 NAND2_X2 _5805_ (.A1(_1077_),
    .A2(_1081_),
    .ZN(_3762_));
 AND2_X1 _5806_ (.A1(_3548_),
    .A2(_1065_),
    .ZN(_1082_));
 INV_X1 _5807_ (.A(_0945_),
    .ZN(_1083_));
 AND4_X1 _5808_ (.A1(_0624_),
    .A2(_0943_),
    .A3(_0633_),
    .A4(_0636_),
    .ZN(_1084_));
 OAI21_X2 _5809_ (.A(_1082_),
    .B1(_1083_),
    .B2(_1084_),
    .ZN(_1085_));
 AND2_X1 _5810_ (.A1(_1065_),
    .A2(_3547_),
    .ZN(_1086_));
 NOR2_X2 _5811_ (.A1(_1070_),
    .A2(_1086_),
    .ZN(_1087_));
 AOI21_X2 _5812_ (.A(_1066_),
    .B1(_1085_),
    .B2(_1087_),
    .ZN(_1088_));
 NAND2_X1 _5813_ (.A1(_3548_),
    .A2(_1065_),
    .ZN(_1089_));
 AOI21_X2 _5814_ (.A(_1089_),
    .B1(_0945_),
    .B2(_0944_),
    .ZN(_1090_));
 OR2_X1 _5815_ (.A1(_1070_),
    .A2(_1086_),
    .ZN(_1091_));
 NOR3_X2 _5816_ (.A1(_3584_),
    .A2(_1090_),
    .A3(_1091_),
    .ZN(_1092_));
 NOR2_X2 _5817_ (.A1(_1088_),
    .A2(_1092_),
    .ZN(_3746_));
 XOR2_X2 _5818_ (.A(_1065_),
    .B(_1076_),
    .Z(_1093_));
 INV_X1 _5819_ (.A(_1093_),
    .ZN(_3750_));
 INV_X1 _5820_ (.A(_3591_),
    .ZN(_1094_));
 INV_X1 _5821_ (.A(_3601_),
    .ZN(_1095_));
 INV_X1 _5822_ (.A(_3609_),
    .ZN(_1096_));
 INV_X1 _5823_ (.A(_3515_),
    .ZN(_1097_));
 AOI21_X1 _5824_ (.A(_3301_),
    .B1(_0527_),
    .B2(_3302_),
    .ZN(_1098_));
 INV_X1 _5825_ (.A(_3516_),
    .ZN(_1099_));
 OAI21_X2 _5826_ (.A(_1097_),
    .B1(_1098_),
    .B2(_1099_),
    .ZN(_1100_));
 AOI21_X1 _5827_ (.A(_3613_),
    .B1(_1100_),
    .B2(_3614_),
    .ZN(_1101_));
 INV_X1 _5828_ (.A(_3610_),
    .ZN(_1102_));
 OAI21_X1 _5829_ (.A(_1096_),
    .B1(_1101_),
    .B2(_1102_),
    .ZN(_1103_));
 AOI21_X1 _5830_ (.A(_3605_),
    .B1(_1103_),
    .B2(_3606_),
    .ZN(_1104_));
 INV_X1 _5831_ (.A(_3602_),
    .ZN(_1105_));
 OAI21_X2 _5832_ (.A(_1095_),
    .B1(_1104_),
    .B2(_1105_),
    .ZN(_1106_));
 CLKBUF_X2 _5833_ (.A(_3598_),
    .Z(_1107_));
 AND2_X1 _5834_ (.A1(_3622_),
    .A2(_1107_),
    .ZN(_1108_));
 AOI221_X2 _5835_ (.A(_3621_),
    .B1(_1106_),
    .B2(_1108_),
    .C1(_3597_),
    .C2(_3622_),
    .ZN(_1109_));
 INV_X1 _5836_ (.A(_3594_),
    .ZN(_1110_));
 OAI21_X1 _5837_ (.A(_1094_),
    .B1(_1109_),
    .B2(_1110_),
    .ZN(_1111_));
 AOI21_X1 _5838_ (.A(_3617_),
    .B1(_1111_),
    .B2(_3618_),
    .ZN(_1112_));
 XOR2_X2 _5839_ (.A(_3588_),
    .B(_1112_),
    .Z(_1113_));
 INV_X1 _5840_ (.A(_1113_),
    .ZN(_3766_));
 AND2_X2 _5841_ (.A1(_3622_),
    .A2(_3594_),
    .ZN(_1114_));
 AND2_X1 _5842_ (.A1(_1107_),
    .A2(_3601_),
    .ZN(_1115_));
 OAI21_X4 _5843_ (.A(_1114_),
    .B1(_1115_),
    .B2(_3597_),
    .ZN(_1116_));
 NAND3_X4 _5844_ (.A1(_1107_),
    .A2(_3602_),
    .A3(_1114_),
    .ZN(_1117_));
 NOR2_X1 _5845_ (.A1(_3609_),
    .A2(_3613_),
    .ZN(_1118_));
 AOI21_X2 _5846_ (.A(_3515_),
    .B1(_0913_),
    .B2(_3516_),
    .ZN(_1119_));
 INV_X1 _5847_ (.A(_3614_),
    .ZN(_1120_));
 OAI21_X2 _5848_ (.A(_1118_),
    .B1(_1119_),
    .B2(_1120_),
    .ZN(_1121_));
 OAI21_X1 _5849_ (.A(_3606_),
    .B1(_3609_),
    .B2(_3610_),
    .ZN(_1122_));
 INV_X1 _5850_ (.A(_1122_),
    .ZN(_1123_));
 AOI21_X4 _5851_ (.A(_3605_),
    .B1(_1121_),
    .B2(_1123_),
    .ZN(_1124_));
 OAI21_X4 _5852_ (.A(_1116_),
    .B1(_1124_),
    .B2(_1117_),
    .ZN(_1125_));
 NAND2_X1 _5853_ (.A1(_3592_),
    .A2(_3621_),
    .ZN(_1126_));
 NAND2_X1 _5854_ (.A1(_1094_),
    .A2(_1126_),
    .ZN(_1127_));
 NOR2_X1 _5855_ (.A1(_1125_),
    .A2(_1127_),
    .ZN(_1128_));
 XOR2_X2 _5856_ (.A(_3618_),
    .B(_1128_),
    .Z(_1129_));
 INV_X1 _5857_ (.A(_1129_),
    .ZN(_3792_));
 XNOR2_X2 _5858_ (.A(_3594_),
    .B(_1109_),
    .ZN(_3770_));
 OAI21_X1 _5859_ (.A(_1095_),
    .B1(_1124_),
    .B2(_1105_),
    .ZN(_1130_));
 AOI21_X2 _5860_ (.A(_3597_),
    .B1(_1130_),
    .B2(_1107_),
    .ZN(_1131_));
 XNOR2_X2 _5861_ (.A(_3622_),
    .B(_1131_),
    .ZN(_3796_));
 XNOR2_X2 _5862_ (.A(_1107_),
    .B(_1106_),
    .ZN(_1132_));
 INV_X1 _5863_ (.A(_1132_),
    .ZN(_3776_));
 XNOR2_X2 _5864_ (.A(_3602_),
    .B(_1124_),
    .ZN(_3780_));
 BUF_X8 _5865_ (.A(_0899_),
    .Z(_3670_));
 INV_X1 _5866_ (.A(_3613_),
    .ZN(_1133_));
 OAI21_X1 _5867_ (.A(_1133_),
    .B1(_1119_),
    .B2(_1120_),
    .ZN(_1134_));
 XNOR2_X2 _5868_ (.A(_3610_),
    .B(_1134_),
    .ZN(_1135_));
 XNOR2_X1 _5869_ (.A(_3606_),
    .B(_1103_),
    .ZN(_1136_));
 NAND2_X1 _5870_ (.A1(_1135_),
    .A2(_1136_),
    .ZN(_1137_));
 NOR2_X1 _5871_ (.A1(_3780_),
    .A2(_1137_),
    .ZN(_1138_));
 XNOR2_X2 _5872_ (.A(_3614_),
    .B(_1100_),
    .ZN(_1139_));
 NAND3_X1 _5873_ (.A1(_3660_),
    .A2(_3659_),
    .A3(_1139_),
    .ZN(_1140_));
 INV_X1 _5874_ (.A(_1140_),
    .ZN(_1141_));
 NAND3_X1 _5875_ (.A1(_1132_),
    .A2(_1138_),
    .A3(_1141_),
    .ZN(_1142_));
 NOR3_X2 _5876_ (.A1(_3770_),
    .A2(_3796_),
    .A3(_1142_),
    .ZN(_1143_));
 NAND2_X1 _5877_ (.A1(_1129_),
    .A2(_1143_),
    .ZN(_1144_));
 OAI21_X2 _5878_ (.A(_3670_),
    .B1(_3766_),
    .B2(_1144_),
    .ZN(_1145_));
 NOR4_X4 _5879_ (.A1(_1127_),
    .A2(_3617_),
    .A3(_3587_),
    .A4(_1125_),
    .ZN(_1146_));
 NOR3_X2 _5880_ (.A1(_3618_),
    .A2(_3587_),
    .A3(_3617_),
    .ZN(_1147_));
 NOR2_X1 _5881_ (.A1(_3588_),
    .A2(_3587_),
    .ZN(_1148_));
 OR3_X4 _5882_ (.A1(_1146_),
    .A2(_1147_),
    .A3(_1148_),
    .ZN(_1149_));
 OAI21_X1 _5883_ (.A(_3564_),
    .B1(_3401_),
    .B2(_0966_),
    .ZN(_1150_));
 AOI21_X1 _5884_ (.A(_0958_),
    .B1(_0959_),
    .B2(_1150_),
    .ZN(_1151_));
 OR2_X2 _5885_ (.A1(_1151_),
    .A2(_3559_),
    .ZN(_1152_));
 XOR2_X2 _5886_ (.A(_1059_),
    .B(_1152_),
    .Z(_1153_));
 NAND2_X1 _5887_ (.A1(_1149_),
    .A2(_1153_),
    .ZN(_1154_));
 NOR3_X4 _5888_ (.A1(_1147_),
    .A2(_1146_),
    .A3(_1148_),
    .ZN(_1155_));
 NAND2_X1 _5889_ (.A1(_1155_),
    .A2(net34),
    .ZN(_1156_));
 XNOR2_X2 _5890_ (.A(_0179_),
    .B(_0699_),
    .ZN(_1157_));
 XNOR2_X2 _5891_ (.A(_0712_),
    .B(_1157_),
    .ZN(_1158_));
 AND2_X1 _5892_ (.A1(_3382_),
    .A2(_3378_),
    .ZN(_1159_));
 OAI211_X2 _5893_ (.A(_0766_),
    .B(_1159_),
    .C1(_0768_),
    .C2(_0767_),
    .ZN(_1160_));
 AOI21_X2 _5894_ (.A(_3377_),
    .B1(_3381_),
    .B2(_3378_),
    .ZN(_1161_));
 AOI21_X2 _5895_ (.A(_1038_),
    .B1(_1160_),
    .B2(_1161_),
    .ZN(_1162_));
 AND3_X1 _5896_ (.A1(_1038_),
    .A2(_1160_),
    .A3(_1161_),
    .ZN(_1163_));
 OAI221_X2 _5897_ (.A(_1158_),
    .B1(_1162_),
    .B2(_1163_),
    .C1(_0714_),
    .C2(net213),
    .ZN(_1164_));
 NOR3_X1 _5898_ (.A1(net213),
    .A2(_3554_),
    .A3(_3542_),
    .ZN(_1165_));
 AOI21_X1 _5899_ (.A(_1040_),
    .B1(_1160_),
    .B2(_1161_),
    .ZN(_1166_));
 NAND4_X1 _5900_ (.A1(_0698_),
    .A2(_0741_),
    .A3(_1165_),
    .A4(_1166_),
    .ZN(_1167_));
 AND3_X1 _5901_ (.A1(_1040_),
    .A2(_1160_),
    .A3(_1161_),
    .ZN(_1168_));
 NAND4_X1 _5902_ (.A1(_0698_),
    .A2(_0741_),
    .A3(_1165_),
    .A4(_1168_),
    .ZN(_1169_));
 AND3_X4 _5903_ (.A1(_1164_),
    .A2(_1167_),
    .A3(_1169_),
    .ZN(_1170_));
 XOR2_X1 _5904_ (.A(_0712_),
    .B(_1157_),
    .Z(_1171_));
 OAI21_X1 _5905_ (.A(_1171_),
    .B1(_1166_),
    .B2(_1168_),
    .ZN(_1172_));
 OAI211_X2 _5906_ (.A(_1158_),
    .B(_1162_),
    .C1(_3396_),
    .C2(_0737_),
    .ZN(_1173_));
 OAI211_X2 _5907_ (.A(_1158_),
    .B(_1163_),
    .C1(_3396_),
    .C2(_0737_),
    .ZN(_1174_));
 AND3_X4 _5908_ (.A1(_1172_),
    .A2(_1173_),
    .A3(_1174_),
    .ZN(_1175_));
 AOI21_X2 _5909_ (.A(net18),
    .B1(_1170_),
    .B2(_1175_),
    .ZN(_1176_));
 INV_X1 _5910_ (.A(_3582_),
    .ZN(_1177_));
 XNOR2_X2 _5911_ (.A(_0203_),
    .B(_0450_),
    .ZN(_1178_));
 NAND3_X1 _5912_ (.A1(_3146_),
    .A2(_3145_),
    .A3(_1178_),
    .ZN(_1179_));
 NOR3_X2 _5913_ (.A1(_3230_),
    .A2(_3226_),
    .A3(_1179_),
    .ZN(_1180_));
 NAND4_X2 _5914_ (.A1(_0340_),
    .A2(_0563_),
    .A3(_0621_),
    .A4(_1180_),
    .ZN(_1181_));
 NOR4_X2 _5915_ (.A1(_3578_),
    .A2(_3546_),
    .A3(_3550_),
    .A4(_1181_),
    .ZN(_1182_));
 NAND3_X1 _5916_ (.A1(_0763_),
    .A2(_1177_),
    .A3(_1182_),
    .ZN(_1183_));
 AND2_X2 _5917_ (.A1(net18),
    .A2(_1183_),
    .ZN(_1184_));
 AND2_X2 _5918_ (.A1(_1170_),
    .A2(_1175_),
    .ZN(_1185_));
 AOI21_X4 _5919_ (.A(_1176_),
    .B1(_1184_),
    .B2(_1185_),
    .ZN(_1186_));
 MUX2_X2 _5920_ (.A(_1154_),
    .B(_1156_),
    .S(_1186_),
    .Z(_1187_));
 XNOR2_X2 _5921_ (.A(net131),
    .B(_1152_),
    .ZN(_1188_));
 NAND2_X1 _5922_ (.A1(_1155_),
    .A2(_1188_),
    .ZN(_1189_));
 NAND2_X1 _5923_ (.A1(_1149_),
    .A2(_1188_),
    .ZN(_1190_));
 MUX2_X2 _5924_ (.A(_1189_),
    .B(_1190_),
    .S(_1186_),
    .Z(_1191_));
 INV_X1 _5925_ (.A(_3235_),
    .ZN(_1192_));
 OAI21_X1 _5926_ (.A(_1192_),
    .B1(_0480_),
    .B2(_0632_),
    .ZN(_1193_));
 AOI21_X1 _5927_ (.A(_3231_),
    .B1(_1193_),
    .B2(_3232_),
    .ZN(_1194_));
 XOR2_X2 _5928_ (.A(_3228_),
    .B(_1194_),
    .Z(_1195_));
 INV_X1 _5929_ (.A(_1195_),
    .ZN(_3444_));
 NOR2_X1 _5930_ (.A1(_3452_),
    .A2(_3456_),
    .ZN(_1196_));
 NAND4_X2 _5931_ (.A1(_0476_),
    .A2(_0486_),
    .A3(_0487_),
    .A4(_1196_),
    .ZN(_1197_));
 OAI21_X1 _5932_ (.A(_0905_),
    .B1(_0638_),
    .B2(_0637_),
    .ZN(_1198_));
 NOR4_X2 _5933_ (.A1(_3570_),
    .A2(_3444_),
    .A3(_1197_),
    .A4(_1198_),
    .ZN(_1199_));
 NAND3_X1 _5934_ (.A1(_0947_),
    .A2(_1093_),
    .A3(_1199_),
    .ZN(_1200_));
 OAI211_X2 _5935_ (.A(_1077_),
    .B(_1081_),
    .C1(_1088_),
    .C2(_1092_),
    .ZN(_1201_));
 OAI21_X2 _5936_ (.A(net10),
    .B1(_1200_),
    .B2(_1201_),
    .ZN(_1202_));
 NOR2_X2 _5937_ (.A1(_1069_),
    .A2(_1066_),
    .ZN(_1203_));
 OAI21_X2 _5938_ (.A(_1203_),
    .B1(_1091_),
    .B2(_1090_),
    .ZN(_1204_));
 AND2_X2 _5939_ (.A1(_3576_),
    .A2(_1071_),
    .ZN(_1205_));
 NOR2_X2 _5940_ (.A1(_3575_),
    .A2(_1205_),
    .ZN(_1206_));
 AOI21_X1 _5941_ (.A(_1063_),
    .B1(_1204_),
    .B2(_1206_),
    .ZN(_1207_));
 AOI21_X1 _5942_ (.A(net18),
    .B1(_1204_),
    .B2(_1206_),
    .ZN(_1208_));
 MUX2_X2 _5943_ (.A(_1207_),
    .B(_1208_),
    .S(net131),
    .Z(_1209_));
 AND3_X1 _5944_ (.A1(_1063_),
    .A2(_1204_),
    .A3(_1206_),
    .ZN(_1210_));
 NAND2_X1 _5945_ (.A1(_3576_),
    .A2(_3584_),
    .ZN(_1211_));
 AOI21_X4 _5946_ (.A(_1211_),
    .B1(_1087_),
    .B2(_1085_),
    .ZN(_1212_));
 OR2_X2 _5947_ (.A1(_3575_),
    .A2(_1205_),
    .ZN(_1213_));
 NOR3_X1 _5948_ (.A1(net67),
    .A2(_1212_),
    .A3(_1213_),
    .ZN(_1214_));
 MUX2_X2 _5949_ (.A(_1210_),
    .B(_1214_),
    .S(net131),
    .Z(_1215_));
 NAND2_X4 _5950_ (.A1(_1170_),
    .A2(_1175_),
    .ZN(_1216_));
 NOR4_X2 _5951_ (.A1(_1202_),
    .A2(_1209_),
    .A3(_1215_),
    .A4(_1216_),
    .ZN(_1217_));
 OAI211_X2 _5952_ (.A(_0234_),
    .B(_1061_),
    .C1(_1212_),
    .C2(_1213_),
    .ZN(_1218_));
 OAI21_X1 _5953_ (.A(net67),
    .B1(_1212_),
    .B2(_1213_),
    .ZN(_1219_));
 MUX2_X2 _5954_ (.A(_1218_),
    .B(_1219_),
    .S(_1059_),
    .Z(_1220_));
 NAND3_X1 _5955_ (.A1(_1063_),
    .A2(_1204_),
    .A3(_1206_),
    .ZN(_1221_));
 NAND3_X1 _5956_ (.A1(_0234_),
    .A2(_1204_),
    .A3(_1206_),
    .ZN(_1222_));
 MUX2_X2 _5957_ (.A(_1221_),
    .B(_1222_),
    .S(_1059_),
    .Z(_1223_));
 AOI221_X2 _5958_ (.A(_1202_),
    .B1(_1220_),
    .B2(_1223_),
    .C1(_1170_),
    .C2(_1175_),
    .ZN(_1224_));
 OR2_X2 _5959_ (.A1(_1217_),
    .A2(_1224_),
    .ZN(_1225_));
 NOR4_X2 _5960_ (.A1(net10),
    .A2(_1209_),
    .A3(_1215_),
    .A4(_1185_),
    .ZN(_1226_));
 NAND3_X1 _5961_ (.A1(_0518_),
    .A2(_1170_),
    .A3(_1175_),
    .ZN(_1227_));
 AOI21_X1 _5962_ (.A(_1227_),
    .B1(_1223_),
    .B2(_1220_),
    .ZN(_1228_));
 OR2_X2 _5963_ (.A1(_1226_),
    .A2(_1228_),
    .ZN(_1229_));
 OAI211_X4 _5964_ (.A(_1187_),
    .B(_1191_),
    .C1(_1225_),
    .C2(_1229_),
    .ZN(_1230_));
 NOR2_X2 _5965_ (.A1(_1217_),
    .A2(_1224_),
    .ZN(_1231_));
 NOR2_X1 _5966_ (.A1(_1155_),
    .A2(_1188_),
    .ZN(_1232_));
 NOR2_X1 _5967_ (.A1(_1149_),
    .A2(_1188_),
    .ZN(_1233_));
 MUX2_X1 _5968_ (.A(_1232_),
    .B(_1233_),
    .S(_1186_),
    .Z(_1234_));
 NOR2_X1 _5969_ (.A1(_1149_),
    .A2(_1153_),
    .ZN(_1235_));
 NOR2_X1 _5970_ (.A1(_1155_),
    .A2(net34),
    .ZN(_1236_));
 MUX2_X1 _5971_ (.A(_1235_),
    .B(_1236_),
    .S(_1186_),
    .Z(_1237_));
 NAND2_X2 _5972_ (.A1(_1223_),
    .A2(_1220_),
    .ZN(_1238_));
 XNOR2_X2 _5973_ (.A(_1216_),
    .B(_1238_),
    .ZN(_1239_));
 OAI221_X2 _5974_ (.A(_1231_),
    .B1(_1237_),
    .B2(_1234_),
    .C1(_1239_),
    .C2(net10),
    .ZN(_1240_));
 NAND2_X4 _5975_ (.A1(_1240_),
    .A2(_1230_),
    .ZN(_1241_));
 XNOR2_X2 _5976_ (.A(_1241_),
    .B(_1145_),
    .ZN(_3623_));
 INV_X1 _5977_ (.A(_3433_),
    .ZN(_1242_));
 AOI21_X1 _5978_ (.A(_3445_),
    .B1(_0915_),
    .B2(_0863_),
    .ZN(_1243_));
 OAI21_X2 _5979_ (.A(_0850_),
    .B1(_1243_),
    .B2(_0865_),
    .ZN(_1244_));
 AOI21_X1 _5980_ (.A(_3437_),
    .B1(_1244_),
    .B2(_0867_),
    .ZN(_1245_));
 OAI21_X1 _5981_ (.A(_1242_),
    .B1(_1245_),
    .B2(_0982_),
    .ZN(_1246_));
 XNOR2_X2 _5982_ (.A(_0979_),
    .B(_1246_),
    .ZN(_3628_));
 INV_X1 _5983_ (.A(_1136_),
    .ZN(_3784_));
 INV_X1 _5984_ (.A(_3770_),
    .ZN(_1247_));
 AND2_X1 _5985_ (.A1(_3661_),
    .A2(_1139_),
    .ZN(_1248_));
 NAND2_X1 _5986_ (.A1(_1138_),
    .A2(_1248_),
    .ZN(_1249_));
 NOR3_X1 _5987_ (.A1(_3796_),
    .A2(_3776_),
    .A3(_1249_),
    .ZN(_1250_));
 NAND3_X1 _5988_ (.A1(_1129_),
    .A2(_1247_),
    .A3(_1250_),
    .ZN(_1251_));
 NAND2_X1 _5989_ (.A1(_3670_),
    .A2(_1251_),
    .ZN(_1252_));
 XNOR2_X1 _5990_ (.A(_1113_),
    .B(_1252_),
    .ZN(_3627_));
 NOR2_X1 _5991_ (.A1(net228),
    .A2(_1143_),
    .ZN(_1253_));
 XNOR2_X1 _5992_ (.A(_3792_),
    .B(_1253_),
    .ZN(_3665_));
 NOR2_X1 _5993_ (.A1(net228),
    .A2(_1250_),
    .ZN(_1254_));
 XNOR2_X1 _5994_ (.A(_3770_),
    .B(_1254_),
    .ZN(_3631_));
 NAND2_X1 _5995_ (.A1(_3670_),
    .A2(_1142_),
    .ZN(_1255_));
 XOR2_X2 _5996_ (.A(_3796_),
    .B(_1255_),
    .Z(_3635_));
 NAND2_X1 _5997_ (.A1(_3670_),
    .A2(_1249_),
    .ZN(_1256_));
 XNOR2_X1 _5998_ (.A(_1132_),
    .B(_1256_),
    .ZN(_3639_));
 OAI21_X1 _5999_ (.A(_3670_),
    .B1(_1137_),
    .B2(_1140_),
    .ZN(_1257_));
 XOR2_X2 _6000_ (.A(_3780_),
    .B(_1257_),
    .Z(_3643_));
 AOI21_X1 _6001_ (.A(_0901_),
    .B1(_1135_),
    .B2(_1248_),
    .ZN(_1258_));
 XNOR2_X1 _6002_ (.A(_3784_),
    .B(_1258_),
    .ZN(_3647_));
 INV_X1 _6003_ (.A(_1135_),
    .ZN(_3788_));
 NOR2_X1 _6004_ (.A1(_3686_),
    .A2(_1141_),
    .ZN(_1259_));
 XNOR2_X1 _6005_ (.A(_3788_),
    .B(_1259_),
    .ZN(_3651_));
 INV_X1 _6006_ (.A(_1139_),
    .ZN(_3714_));
 NOR2_X1 _6007_ (.A1(_3661_),
    .A2(_3686_),
    .ZN(_1260_));
 XNOR2_X1 _6008_ (.A(_3714_),
    .B(_1260_),
    .ZN(_3655_));
 INV_X1 _6009_ (.A(_3659_),
    .ZN(_3517_));
 MUX2_X1 _6010_ (.A(_3662_),
    .B(_3517_),
    .S(_0901_),
    .Z(_2959_));
 INV_X1 _6011_ (.A(_2959_),
    .ZN(_2963_));
 INV_X1 _6012_ (.A(_3667_),
    .ZN(_1261_));
 INV_X1 _6013_ (.A(_3637_),
    .ZN(_1262_));
 INV_X1 _6014_ (.A(_3645_),
    .ZN(_1263_));
 INV_X1 _6015_ (.A(_3653_),
    .ZN(_1264_));
 INV_X1 _6016_ (.A(_3663_),
    .ZN(_1265_));
 INV_X1 _6017_ (.A(_3664_),
    .ZN(_1266_));
 OAI21_X1 _6018_ (.A(_1265_),
    .B1(_1266_),
    .B2(_2958_),
    .ZN(_1267_));
 AOI21_X2 _6019_ (.A(_3657_),
    .B1(_1267_),
    .B2(_3658_),
    .ZN(_1268_));
 BUF_X1 _6020_ (.A(_3654_),
    .Z(_1269_));
 INV_X1 _6021_ (.A(_1269_),
    .ZN(_1270_));
 OAI21_X1 _6022_ (.A(_1264_),
    .B1(_1268_),
    .B2(_1270_),
    .ZN(_1271_));
 AOI21_X2 _6023_ (.A(_3649_),
    .B1(_1271_),
    .B2(_3650_),
    .ZN(_1272_));
 CLKBUF_X2 _6024_ (.A(_3646_),
    .Z(_1273_));
 INV_X1 _6025_ (.A(_1273_),
    .ZN(_1274_));
 OAI21_X1 _6026_ (.A(_1263_),
    .B1(_1272_),
    .B2(_1274_),
    .ZN(_1275_));
 AOI21_X2 _6027_ (.A(_3641_),
    .B1(_1275_),
    .B2(_3642_),
    .ZN(_1276_));
 CLKBUF_X2 _6028_ (.A(_3638_),
    .Z(_1277_));
 INV_X1 _6029_ (.A(_1277_),
    .ZN(_1278_));
 OAI21_X1 _6030_ (.A(_1262_),
    .B1(_1276_),
    .B2(_1278_),
    .ZN(_1279_));
 AOI21_X2 _6031_ (.A(_3633_),
    .B1(_1279_),
    .B2(_3634_),
    .ZN(_1280_));
 CLKBUF_X2 _6032_ (.A(_3668_),
    .Z(_1281_));
 INV_X1 _6033_ (.A(_1281_),
    .ZN(_1282_));
 OAI21_X1 _6034_ (.A(_1261_),
    .B1(_1280_),
    .B2(_1282_),
    .ZN(_1283_));
 AOI21_X2 _6035_ (.A(_3629_),
    .B1(_1283_),
    .B2(_3630_),
    .ZN(_1284_));
 XNOR2_X2 _6036_ (.A(_3626_),
    .B(_1284_),
    .ZN(_3852_));
 XNOR2_X2 _6037_ (.A(_1281_),
    .B(_1280_),
    .ZN(_3810_));
 XNOR2_X2 _6038_ (.A(_1277_),
    .B(_1276_),
    .ZN(_3818_));
 INV_X1 _6039_ (.A(_3649_),
    .ZN(_1285_));
 INV_X1 _6040_ (.A(_3657_),
    .ZN(_1286_));
 INV_X1 _6041_ (.A(_3658_),
    .ZN(_1287_));
 OAI21_X1 _6042_ (.A(_1286_),
    .B1(_2961_),
    .B2(_1287_),
    .ZN(_1288_));
 AOI21_X2 _6043_ (.A(_3653_),
    .B1(_1288_),
    .B2(_1269_),
    .ZN(_1289_));
 INV_X1 _6044_ (.A(_3650_),
    .ZN(_1290_));
 OAI21_X1 _6045_ (.A(_1285_),
    .B1(_1289_),
    .B2(_1290_),
    .ZN(_1291_));
 AOI21_X2 _6046_ (.A(_3645_),
    .B1(_1291_),
    .B2(_1273_),
    .ZN(_1292_));
 XNOR2_X2 _6047_ (.A(_3642_),
    .B(_1292_),
    .ZN(_3822_));
 INV_X1 _6048_ (.A(_3822_),
    .ZN(_3737_));
 XNOR2_X2 _6049_ (.A(_1273_),
    .B(_1272_),
    .ZN(_3826_));
 INV_X1 _6050_ (.A(_3826_),
    .ZN(_3736_));
 INV_X1 _6051_ (.A(_3677_),
    .ZN(_1293_));
 INV_X1 _6052_ (.A(_3683_),
    .ZN(_1294_));
 INV_X1 _6053_ (.A(_3690_),
    .ZN(_1295_));
 INV_X1 _6054_ (.A(_3696_),
    .ZN(_1296_));
 INV_X1 _6055_ (.A(_3702_),
    .ZN(_1297_));
 INV_X1 _6056_ (.A(_3708_),
    .ZN(_1298_));
 AOI21_X2 _6057_ (.A(_3711_),
    .B1(_3712_),
    .B2(_0005_),
    .ZN(_1299_));
 INV_X1 _6058_ (.A(_3709_),
    .ZN(_1300_));
 OAI21_X4 _6059_ (.A(_1298_),
    .B1(_1300_),
    .B2(_1299_),
    .ZN(_1301_));
 AOI21_X4 _6060_ (.A(_3705_),
    .B1(_3706_),
    .B2(_1301_),
    .ZN(_1302_));
 INV_X1 _6061_ (.A(_3703_),
    .ZN(_1303_));
 OAI21_X4 _6062_ (.A(_1297_),
    .B1(_1303_),
    .B2(_1302_),
    .ZN(_1304_));
 AOI21_X4 _6063_ (.A(_3699_),
    .B1(_1304_),
    .B2(_3700_),
    .ZN(_1305_));
 INV_X1 _6064_ (.A(_3697_),
    .ZN(_1306_));
 OAI21_X4 _6065_ (.A(_1296_),
    .B1(_1305_),
    .B2(_1306_),
    .ZN(_1307_));
 AOI21_X4 _6066_ (.A(_3693_),
    .B1(_3694_),
    .B2(_1307_),
    .ZN(_1308_));
 INV_X1 _6067_ (.A(_3691_),
    .ZN(_1309_));
 OAI21_X4 _6068_ (.A(_1295_),
    .B1(_1309_),
    .B2(_1308_),
    .ZN(_1310_));
 AOI21_X4 _6069_ (.A(_3687_),
    .B1(_3688_),
    .B2(_1310_),
    .ZN(_1311_));
 INV_X1 _6070_ (.A(_3684_),
    .ZN(_1312_));
 OAI21_X4 _6071_ (.A(_1294_),
    .B1(_1312_),
    .B2(_1311_),
    .ZN(_1313_));
 AOI21_X4 _6072_ (.A(_3680_),
    .B1(_1313_),
    .B2(_3681_),
    .ZN(_1314_));
 INV_X1 _6073_ (.A(_3678_),
    .ZN(_1315_));
 OAI21_X4 _6074_ (.A(_1293_),
    .B1(_1315_),
    .B2(_1314_),
    .ZN(_1316_));
 AND2_X1 _6075_ (.A1(_3672_),
    .A2(_3675_),
    .ZN(_1317_));
 NAND2_X4 _6076_ (.A1(_1317_),
    .A2(_1316_),
    .ZN(_1318_));
 AOI21_X4 _6077_ (.A(_3671_),
    .B1(_3674_),
    .B2(_3672_),
    .ZN(_1319_));
 NAND2_X4 _6078_ (.A1(_1318_),
    .A2(_1319_),
    .ZN(_3856_));
 INV_X8 _6079_ (.A(_3856_),
    .ZN(_1320_));
 BUF_X16 _6080_ (.A(_1320_),
    .Z(_1321_));
 BUF_X32 _6081_ (.A(_1321_),
    .Z(_3875_));
 XNOR2_X2 _6082_ (.A(_0867_),
    .B(_1244_),
    .ZN(_1322_));
 INV_X1 _6083_ (.A(_1322_),
    .ZN(_3632_));
 INV_X1 _6084_ (.A(_3716_),
    .ZN(_1323_));
 INV_X1 _6085_ (.A(_3519_),
    .ZN(_1324_));
 INV_X1 _6086_ (.A(_3526_),
    .ZN(_1325_));
 AOI21_X1 _6087_ (.A(_3530_),
    .B1(_2956_),
    .B2(_3531_),
    .ZN(_1326_));
 INV_X1 _6088_ (.A(_3527_),
    .ZN(_1327_));
 OAI21_X1 _6089_ (.A(_1325_),
    .B1(_1326_),
    .B2(_1327_),
    .ZN(_1328_));
 AOI21_X1 _6090_ (.A(_3522_),
    .B1(_1328_),
    .B2(_3523_),
    .ZN(_1329_));
 INV_X1 _6091_ (.A(_3520_),
    .ZN(_1330_));
 OAI21_X2 _6092_ (.A(_1324_),
    .B1(_1329_),
    .B2(_1330_),
    .ZN(_1331_));
 XNOR2_X2 _6093_ (.A(_1323_),
    .B(_1331_),
    .ZN(_3717_));
 INV_X1 _6094_ (.A(_3717_),
    .ZN(_3841_));
 INV_X1 _6095_ (.A(_3641_),
    .ZN(_1332_));
 INV_X1 _6096_ (.A(_3642_),
    .ZN(_1333_));
 OAI21_X1 _6097_ (.A(_1332_),
    .B1(_1292_),
    .B2(_1333_),
    .ZN(_1334_));
 AOI21_X2 _6098_ (.A(_3637_),
    .B1(_1334_),
    .B2(_1277_),
    .ZN(_1335_));
 XNOR2_X2 _6099_ (.A(_3634_),
    .B(_1335_),
    .ZN(_3814_));
 INV_X1 _6100_ (.A(_3633_),
    .ZN(_1336_));
 INV_X1 _6101_ (.A(_3634_),
    .ZN(_1337_));
 OAI21_X1 _6102_ (.A(_1336_),
    .B1(_1335_),
    .B2(_1337_),
    .ZN(_1338_));
 AOI21_X2 _6103_ (.A(_3667_),
    .B1(_1338_),
    .B2(_1281_),
    .ZN(_1339_));
 XNOR2_X2 _6104_ (.A(_3630_),
    .B(_1339_),
    .ZN(_3804_));
 INV_X1 _6105_ (.A(_3722_),
    .ZN(_1340_));
 INV_X1 _6106_ (.A(_3730_),
    .ZN(_1341_));
 AOI21_X1 _6107_ (.A(_3734_),
    .B1(_3735_),
    .B2(_2966_),
    .ZN(_1342_));
 INV_X1 _6108_ (.A(_3731_),
    .ZN(_1343_));
 OAI21_X2 _6109_ (.A(_1341_),
    .B1(_1342_),
    .B2(_1343_),
    .ZN(_1344_));
 AOI21_X1 _6110_ (.A(_3726_),
    .B1(_1344_),
    .B2(_3727_),
    .ZN(_1345_));
 INV_X1 _6111_ (.A(_3723_),
    .ZN(_1346_));
 OAI21_X2 _6112_ (.A(_1340_),
    .B1(_1345_),
    .B2(_1346_),
    .ZN(_1347_));
 XNOR2_X2 _6113_ (.A(_3720_),
    .B(_1347_),
    .ZN(_4010_));
 AOI21_X2 _6114_ (.A(_0518_),
    .B1(_0965_),
    .B2(_0969_),
    .ZN(_1348_));
 AND2_X1 _6115_ (.A1(_1153_),
    .A2(_1348_),
    .ZN(_1349_));
 AND2_X1 _6116_ (.A1(_1188_),
    .A2(_1348_),
    .ZN(_1350_));
 MUX2_X2 _6117_ (.A(_1349_),
    .B(_1350_),
    .S(_1186_),
    .Z(_1351_));
 NOR2_X1 _6118_ (.A1(_0517_),
    .A2(_1188_),
    .ZN(_1352_));
 NOR2_X1 _6119_ (.A1(_0517_),
    .A2(_1153_),
    .ZN(_1353_));
 MUX2_X2 _6120_ (.A(net67),
    .B(_1184_),
    .S(_1185_),
    .Z(_1354_));
 MUX2_X2 _6121_ (.A(_1352_),
    .B(_1353_),
    .S(_1354_),
    .Z(_1355_));
 NOR2_X1 _6122_ (.A1(_1351_),
    .A2(_1355_),
    .ZN(_3745_));
 XNOR2_X2 _6123_ (.A(_1354_),
    .B(_1153_),
    .ZN(_1356_));
 NAND4_X1 _6124_ (.A1(_0836_),
    .A2(_0965_),
    .A3(_0968_),
    .A4(_0976_),
    .ZN(_1357_));
 AND2_X1 _6125_ (.A1(net10),
    .A2(_1357_),
    .ZN(_1358_));
 XOR2_X2 _6126_ (.A(_1356_),
    .B(_1358_),
    .Z(_3749_));
 BUF_X1 _6127_ (.A(_3751_),
    .Z(_1359_));
 INV_X1 _6128_ (.A(_3567_),
    .ZN(_1360_));
 OR2_X1 _6129_ (.A1(_3433_),
    .A2(_0978_),
    .ZN(_1361_));
 AOI211_X2 _6130_ (.A(_0983_),
    .B(_1361_),
    .C1(_0995_),
    .C2(_0984_),
    .ZN(_1362_));
 OAI21_X1 _6131_ (.A(_3568_),
    .B1(_3572_),
    .B2(_0978_),
    .ZN(_1363_));
 OAI21_X1 _6132_ (.A(_1360_),
    .B1(_1362_),
    .B2(_1363_),
    .ZN(_1364_));
 AOI21_X2 _6133_ (.A(_1359_),
    .B1(_1364_),
    .B2(_3752_),
    .ZN(_1365_));
 XNOR2_X2 _6134_ (.A(net136),
    .B(_1365_),
    .ZN(_3754_));
 AOI21_X2 _6135_ (.A(_1145_),
    .B1(_1230_),
    .B2(net133),
    .ZN(_1366_));
 NOR2_X1 _6136_ (.A1(_1226_),
    .A2(_1228_),
    .ZN(_1367_));
 AOI211_X4 _6137_ (.A(_1234_),
    .B(_1237_),
    .C1(_1231_),
    .C2(_1367_),
    .ZN(_1368_));
 AOI211_X2 _6138_ (.A(_1225_),
    .B(_1229_),
    .C1(_1191_),
    .C2(_1187_),
    .ZN(_1369_));
 NOR3_X4 _6139_ (.A1(_1368_),
    .A2(_0899_),
    .A3(_1369_),
    .ZN(_1370_));
 NOR2_X1 _6140_ (.A1(_1366_),
    .A2(_1370_),
    .ZN(_3753_));
 NOR3_X1 _6141_ (.A1(_3433_),
    .A2(_3567_),
    .A3(_0978_),
    .ZN(_1371_));
 OAI21_X1 _6142_ (.A(_1371_),
    .B1(_1245_),
    .B2(_0982_),
    .ZN(_1372_));
 NOR3_X1 _6143_ (.A1(_3572_),
    .A2(_3567_),
    .A3(_0978_),
    .ZN(_1373_));
 INV_X1 _6144_ (.A(_3568_),
    .ZN(_1374_));
 AOI21_X1 _6145_ (.A(_1373_),
    .B1(_1360_),
    .B2(_1374_),
    .ZN(_1375_));
 AND3_X1 _6146_ (.A1(_3752_),
    .A2(_1372_),
    .A3(_1375_),
    .ZN(_1376_));
 AOI21_X2 _6147_ (.A(_3752_),
    .B1(_1372_),
    .B2(_1375_),
    .ZN(_1377_));
 NOR2_X4 _6148_ (.A1(_1376_),
    .A2(_1377_),
    .ZN(_3758_));
 NOR2_X1 _6149_ (.A1(_3766_),
    .A2(_1251_),
    .ZN(_1378_));
 NOR2_X1 _6150_ (.A1(net228),
    .A2(_1378_),
    .ZN(_1379_));
 AOI21_X2 _6151_ (.A(_1370_),
    .B1(_1379_),
    .B2(_1241_),
    .ZN(_3757_));
 INV_X1 _6152_ (.A(_3629_),
    .ZN(_1380_));
 INV_X1 _6153_ (.A(_2958_),
    .ZN(_1381_));
 AOI21_X1 _6154_ (.A(_3663_),
    .B1(_3664_),
    .B2(_1381_),
    .ZN(_1382_));
 OAI21_X1 _6155_ (.A(_1286_),
    .B1(_1382_),
    .B2(_1287_),
    .ZN(_1383_));
 AOI21_X1 _6156_ (.A(_3653_),
    .B1(_1383_),
    .B2(_1269_),
    .ZN(_1384_));
 OAI21_X1 _6157_ (.A(_1285_),
    .B1(_1384_),
    .B2(_1290_),
    .ZN(_1385_));
 AOI21_X1 _6158_ (.A(_3645_),
    .B1(_1385_),
    .B2(_1273_),
    .ZN(_1386_));
 OAI21_X1 _6159_ (.A(_1332_),
    .B1(_1386_),
    .B2(_1333_),
    .ZN(_1387_));
 AOI21_X1 _6160_ (.A(_3637_),
    .B1(_1387_),
    .B2(_1277_),
    .ZN(_1388_));
 OAI21_X1 _6161_ (.A(_1336_),
    .B1(_1388_),
    .B2(_1337_),
    .ZN(_1389_));
 AOI21_X1 _6162_ (.A(_3667_),
    .B1(_1389_),
    .B2(_1281_),
    .ZN(_1390_));
 INV_X1 _6163_ (.A(_3630_),
    .ZN(_1391_));
 OAI21_X1 _6164_ (.A(_1380_),
    .B1(_1390_),
    .B2(_1391_),
    .ZN(_1392_));
 BUF_X2 _6165_ (.A(_3760_),
    .Z(_1393_));
 AND2_X2 _6166_ (.A1(_1393_),
    .A2(_3626_),
    .ZN(_1394_));
 AOI221_X2 _6167_ (.A(_3759_),
    .B1(_1394_),
    .B2(_1392_),
    .C1(_3625_),
    .C2(_1393_),
    .ZN(_1395_));
 XNOR2_X2 _6168_ (.A(_1395_),
    .B(_3756_),
    .ZN(_3799_));
 AOI21_X2 _6169_ (.A(_1355_),
    .B1(_1358_),
    .B2(_1356_),
    .ZN(_3761_));
 INV_X1 _6170_ (.A(_3764_),
    .ZN(_1396_));
 AND2_X1 _6171_ (.A1(net136),
    .A2(_1396_),
    .ZN(_1397_));
 OAI21_X1 _6172_ (.A(_1397_),
    .B1(_1376_),
    .B2(_1359_),
    .ZN(_1398_));
 OR4_X1 _6173_ (.A1(_1396_),
    .A2(_3747_),
    .A3(_1359_),
    .A4(_1376_),
    .ZN(_1399_));
 NOR3_X1 _6174_ (.A1(net136),
    .A2(_1396_),
    .A3(_3747_),
    .ZN(_1400_));
 AOI21_X1 _6175_ (.A(_1400_),
    .B1(_3747_),
    .B2(_1396_),
    .ZN(_1401_));
 NAND3_X2 _6176_ (.A1(_1398_),
    .A2(_1399_),
    .A3(_1401_),
    .ZN(_3935_));
 BUF_X2 _6177_ (.A(_3768_),
    .Z(_1402_));
 INV_X1 _6178_ (.A(_3793_),
    .ZN(_1403_));
 INV_X1 _6179_ (.A(_3797_),
    .ZN(_1404_));
 INV_X1 _6180_ (.A(_3781_),
    .ZN(_1405_));
 INV_X1 _6181_ (.A(_3789_),
    .ZN(_1406_));
 AOI21_X1 _6182_ (.A(_3715_),
    .B1(_1331_),
    .B2(_3716_),
    .ZN(_1407_));
 INV_X1 _6183_ (.A(_3790_),
    .ZN(_1408_));
 OAI21_X1 _6184_ (.A(_1406_),
    .B1(_1407_),
    .B2(_1408_),
    .ZN(_1409_));
 AOI21_X1 _6185_ (.A(_3785_),
    .B1(_1409_),
    .B2(_3786_),
    .ZN(_1410_));
 INV_X1 _6186_ (.A(_3782_),
    .ZN(_1411_));
 OAI21_X2 _6187_ (.A(_1405_),
    .B1(_1410_),
    .B2(_1411_),
    .ZN(_1412_));
 AOI21_X1 _6188_ (.A(_3777_),
    .B1(_1412_),
    .B2(_3778_),
    .ZN(_1413_));
 INV_X1 _6189_ (.A(_3798_),
    .ZN(_1414_));
 OAI21_X1 _6190_ (.A(_1404_),
    .B1(_1413_),
    .B2(_1414_),
    .ZN(_1415_));
 AOI21_X1 _6191_ (.A(_3771_),
    .B1(_1415_),
    .B2(_3774_),
    .ZN(_1416_));
 INV_X1 _6192_ (.A(_3794_),
    .ZN(_1417_));
 OAI21_X1 _6193_ (.A(_1403_),
    .B1(_1416_),
    .B2(_1417_),
    .ZN(_1418_));
 XNOR2_X2 _6194_ (.A(_1402_),
    .B(_1418_),
    .ZN(_1419_));
 INV_X1 _6195_ (.A(_1419_),
    .ZN(_3944_));
 INV_X1 _6196_ (.A(_3777_),
    .ZN(_1420_));
 INV_X1 _6197_ (.A(_3785_),
    .ZN(_1421_));
 INV_X1 _6198_ (.A(_3715_),
    .ZN(_1422_));
 AOI21_X1 _6199_ (.A(_3519_),
    .B1(_0925_),
    .B2(_3520_),
    .ZN(_1423_));
 OAI21_X1 _6200_ (.A(_1422_),
    .B1(_1423_),
    .B2(_1323_),
    .ZN(_1424_));
 AOI21_X1 _6201_ (.A(_3789_),
    .B1(_1424_),
    .B2(_3790_),
    .ZN(_1425_));
 INV_X1 _6202_ (.A(_3786_),
    .ZN(_1426_));
 OAI21_X2 _6203_ (.A(_1421_),
    .B1(_1425_),
    .B2(_1426_),
    .ZN(_1427_));
 AOI21_X1 _6204_ (.A(_3781_),
    .B1(_1427_),
    .B2(_3782_),
    .ZN(_1428_));
 INV_X1 _6205_ (.A(_3778_),
    .ZN(_1429_));
 OAI21_X2 _6206_ (.A(_1420_),
    .B1(_1428_),
    .B2(_1429_),
    .ZN(_1430_));
 AND2_X1 _6207_ (.A1(_3798_),
    .A2(_3774_),
    .ZN(_1431_));
 AOI221_X2 _6208_ (.A(_3771_),
    .B1(_1431_),
    .B2(_1430_),
    .C1(_3797_),
    .C2(_3772_),
    .ZN(_1432_));
 XNOR2_X2 _6209_ (.A(_1417_),
    .B(_1432_),
    .ZN(_1433_));
 INV_X1 _6210_ (.A(_1433_),
    .ZN(_3948_));
 XNOR2_X1 _6211_ (.A(_3774_),
    .B(_1415_),
    .ZN(_1434_));
 INV_X1 _6212_ (.A(_1434_),
    .ZN(_3952_));
 XNOR2_X2 _6213_ (.A(_1414_),
    .B(_1430_),
    .ZN(_3970_));
 XNOR2_X2 _6214_ (.A(_1429_),
    .B(_1412_),
    .ZN(_3956_));
 XNOR2_X2 _6215_ (.A(_1411_),
    .B(_1427_),
    .ZN(_3960_));
 XNOR2_X1 _6216_ (.A(_3786_),
    .B(_1409_),
    .ZN(_1435_));
 INV_X1 _6217_ (.A(_1435_),
    .ZN(_3964_));
 AOI21_X2 _6218_ (.A(_3763_),
    .B1(_3764_),
    .B2(_3747_),
    .ZN(_1436_));
 INV_X1 _6219_ (.A(_1436_),
    .ZN(_1437_));
 NOR3_X2 _6220_ (.A1(_3567_),
    .A2(_1359_),
    .A3(_1437_),
    .ZN(_1438_));
 OAI21_X2 _6221_ (.A(_1438_),
    .B1(_1363_),
    .B2(_1362_),
    .ZN(_1439_));
 NAND2_X1 _6222_ (.A1(_3748_),
    .A2(_3764_),
    .ZN(_1440_));
 NOR2_X1 _6223_ (.A1(_3752_),
    .A2(_1359_),
    .ZN(_1441_));
 OAI21_X2 _6224_ (.A(_1436_),
    .B1(_1440_),
    .B2(_1441_),
    .ZN(_1442_));
 AND2_X4 _6225_ (.A1(_1439_),
    .A2(_1442_),
    .ZN(_1443_));
 AND4_X2 _6226_ (.A1(_1220_),
    .A2(_1223_),
    .A3(_1216_),
    .A4(_1443_),
    .ZN(_1444_));
 NAND4_X2 _6227_ (.A1(_1170_),
    .A2(_1175_),
    .A3(_1439_),
    .A4(_1442_),
    .ZN(_1445_));
 AOI21_X4 _6228_ (.A(_1445_),
    .B1(_1223_),
    .B2(_1220_),
    .ZN(_1446_));
 NOR4_X4 _6229_ (.A1(_1209_),
    .A2(_1215_),
    .A3(_1216_),
    .A4(_1443_),
    .ZN(_1447_));
 AOI221_X2 _6230_ (.A(_1185_),
    .B1(_1439_),
    .B2(_1442_),
    .C1(_1223_),
    .C2(_1220_),
    .ZN(_1448_));
 NOR4_X4 _6231_ (.A1(_1444_),
    .A2(_1446_),
    .A3(_1447_),
    .A4(_1448_),
    .ZN(_1449_));
 NAND2_X1 _6232_ (.A1(_0519_),
    .A2(net34),
    .ZN(_1450_));
 NAND2_X1 _6233_ (.A1(_0519_),
    .A2(_1188_),
    .ZN(_1451_));
 MUX2_X2 _6234_ (.A(_1450_),
    .B(_1451_),
    .S(_1354_),
    .Z(_1452_));
 NAND2_X1 _6235_ (.A1(net34),
    .A2(_1348_),
    .ZN(_1453_));
 NAND2_X1 _6236_ (.A1(_1188_),
    .A2(_1348_),
    .ZN(_1454_));
 MUX2_X2 _6237_ (.A(_1453_),
    .B(_1454_),
    .S(_1186_),
    .Z(_1455_));
 AOI21_X4 _6238_ (.A(_1449_),
    .B1(_1452_),
    .B2(_1455_),
    .ZN(_1456_));
 OR4_X4 _6239_ (.A1(_1444_),
    .A2(_1446_),
    .A3(_1447_),
    .A4(_1448_),
    .ZN(_1457_));
 NOR3_X4 _6240_ (.A1(_1351_),
    .A2(_1355_),
    .A3(_1457_),
    .ZN(_1458_));
 NOR3_X4 _6241_ (.A1(_0899_),
    .A2(_1456_),
    .A3(_1458_),
    .ZN(_1459_));
 OAI21_X4 _6242_ (.A(_1457_),
    .B1(_1355_),
    .B2(_1351_),
    .ZN(_1460_));
 NAND3_X4 _6243_ (.A1(_1455_),
    .A2(_1452_),
    .A3(_1449_),
    .ZN(_1461_));
 NOR3_X1 _6244_ (.A1(_3644_),
    .A2(_3648_),
    .A3(_3640_),
    .ZN(_1462_));
 NAND3_X1 _6245_ (.A1(_0917_),
    .A2(_1322_),
    .A3(_1462_),
    .ZN(_1463_));
 OR3_X2 _6246_ (.A1(_3666_),
    .A2(_3628_),
    .A3(_1463_),
    .ZN(_1464_));
 NOR4_X4 _6247_ (.A1(_3624_),
    .A2(_3754_),
    .A3(_3758_),
    .A4(_1464_),
    .ZN(_1465_));
 INV_X2 _6248_ (.A(_3935_),
    .ZN(_1466_));
 AOI221_X2 _6249_ (.A(_0900_),
    .B1(_1460_),
    .B2(_1461_),
    .C1(_1465_),
    .C2(_1466_),
    .ZN(_1467_));
 OAI21_X2 _6250_ (.A(_1403_),
    .B1(_1432_),
    .B2(_1417_),
    .ZN(_1468_));
 AOI21_X4 _6251_ (.A(_3767_),
    .B1(_1468_),
    .B2(_1402_),
    .ZN(_1469_));
 AOI21_X4 _6252_ (.A(_1469_),
    .B1(_1240_),
    .B2(_1230_),
    .ZN(_1470_));
 AOI21_X2 _6253_ (.A(_3767_),
    .B1(_3793_),
    .B2(_1402_),
    .ZN(_1471_));
 NAND2_X1 _6254_ (.A1(_1402_),
    .A2(_3794_),
    .ZN(_1472_));
 OAI21_X4 _6255_ (.A(_1471_),
    .B1(_1472_),
    .B2(net140),
    .ZN(_1473_));
 NOR3_X4 _6256_ (.A1(_1473_),
    .A2(net121),
    .A3(_1368_),
    .ZN(_1474_));
 OAI22_X4 _6257_ (.A1(_1459_),
    .A2(_1467_),
    .B1(_1474_),
    .B2(_1470_),
    .ZN(_1475_));
 NAND3_X4 _6258_ (.A1(net219),
    .A2(_1460_),
    .A3(_1461_),
    .ZN(_1476_));
 AOI21_X4 _6259_ (.A(_0900_),
    .B1(_1466_),
    .B2(_1465_),
    .ZN(_1477_));
 OAI21_X4 _6260_ (.A(_1477_),
    .B1(_1458_),
    .B2(_1456_),
    .ZN(_1478_));
 OAI21_X4 _6261_ (.A(_1473_),
    .B1(net121),
    .B2(_1368_),
    .ZN(_1479_));
 NAND3_X4 _6262_ (.A1(_1230_),
    .A2(_1240_),
    .A3(_1469_),
    .ZN(_1480_));
 NAND4_X4 _6263_ (.A1(_1476_),
    .A2(_1478_),
    .A3(_1479_),
    .A4(_1480_),
    .ZN(_1481_));
 INV_X1 _6264_ (.A(_3842_),
    .ZN(_3539_));
 NOR2_X2 _6265_ (.A1(_3539_),
    .A2(_3717_),
    .ZN(_1482_));
 XNOR2_X1 _6266_ (.A(_3790_),
    .B(_1424_),
    .ZN(_1483_));
 INV_X1 _6267_ (.A(_1483_),
    .ZN(_3900_));
 NOR2_X1 _6268_ (.A1(_3964_),
    .A2(_3900_),
    .ZN(_1484_));
 INV_X1 _6269_ (.A(_1484_),
    .ZN(_1485_));
 NOR4_X1 _6270_ (.A1(_3970_),
    .A2(_3956_),
    .A3(_3960_),
    .A4(_1485_),
    .ZN(_1486_));
 AND2_X1 _6271_ (.A1(_1434_),
    .A2(_1486_),
    .ZN(_1487_));
 AND3_X1 _6272_ (.A1(_1433_),
    .A2(_1482_),
    .A3(_1487_),
    .ZN(_1488_));
 AOI221_X2 _6273_ (.A(_1320_),
    .B1(_1481_),
    .B2(_1475_),
    .C1(_1488_),
    .C2(_1419_),
    .ZN(_1489_));
 AOI22_X4 _6274_ (.A1(_1476_),
    .A2(_1478_),
    .B1(_1479_),
    .B2(_1480_),
    .ZN(_1490_));
 NOR4_X4 _6275_ (.A1(_1470_),
    .A2(_1467_),
    .A3(_1459_),
    .A4(_1474_),
    .ZN(_1491_));
 NOR3_X4 _6276_ (.A1(net1),
    .A2(_1490_),
    .A3(_1491_),
    .ZN(_1492_));
 NOR2_X1 _6277_ (.A1(_1489_),
    .A2(_1492_),
    .ZN(_3800_));
 OAI21_X1 _6278_ (.A(_1380_),
    .B1(_1339_),
    .B2(_1391_),
    .ZN(_1493_));
 AOI21_X2 _6279_ (.A(_3625_),
    .B1(_1493_),
    .B2(_3626_),
    .ZN(_1494_));
 XNOR2_X2 _6280_ (.A(_1393_),
    .B(_1494_),
    .ZN(_3847_));
 BUF_X1 _6281_ (.A(_3843_),
    .Z(_1495_));
 NAND4_X1 _6282_ (.A1(_1495_),
    .A2(_1419_),
    .A3(_1433_),
    .A4(_1487_),
    .ZN(_1496_));
 AND2_X1 _6283_ (.A1(net1),
    .A2(_1496_),
    .ZN(_1497_));
 NAND2_X4 _6284_ (.A1(_1475_),
    .A2(_1481_),
    .ZN(_1498_));
 AOI21_X1 _6285_ (.A(_1492_),
    .B1(_1497_),
    .B2(_1498_),
    .ZN(_3848_));
 NOR2_X1 _6286_ (.A1(_1489_),
    .A2(_1492_),
    .ZN(_3851_));
 XOR2_X2 _6287_ (.A(_1498_),
    .B(_1497_),
    .Z(_3803_));
 NOR2_X1 _6288_ (.A1(net229),
    .A2(_1488_),
    .ZN(_1499_));
 XNOR2_X1 _6289_ (.A(_3944_),
    .B(_1499_),
    .ZN(_3809_));
 AOI21_X1 _6290_ (.A(net229),
    .B1(_1487_),
    .B2(_1495_),
    .ZN(_1500_));
 XNOR2_X1 _6291_ (.A(_3948_),
    .B(_1500_),
    .ZN(_3813_));
 AOI21_X1 _6292_ (.A(net229),
    .B1(_1482_),
    .B2(_1486_),
    .ZN(_1501_));
 XNOR2_X1 _6293_ (.A(_3952_),
    .B(_1501_),
    .ZN(_3817_));
 NOR3_X1 _6294_ (.A1(_3956_),
    .A2(_3960_),
    .A3(_1485_),
    .ZN(_1502_));
 AOI21_X1 _6295_ (.A(net229),
    .B1(_1502_),
    .B2(_1495_),
    .ZN(_1503_));
 XNOR2_X1 _6296_ (.A(_3970_),
    .B(_1503_),
    .ZN(_3821_));
 NOR2_X1 _6297_ (.A1(_3960_),
    .A2(_1485_),
    .ZN(_1504_));
 AOI21_X1 _6298_ (.A(_3875_),
    .B1(_1482_),
    .B2(_1504_),
    .ZN(_1505_));
 XNOR2_X1 _6299_ (.A(_3956_),
    .B(_1505_),
    .ZN(_3825_));
 AOI21_X1 _6300_ (.A(net226),
    .B1(_1484_),
    .B2(_1495_),
    .ZN(_1506_));
 XNOR2_X1 _6301_ (.A(_3960_),
    .B(_1506_),
    .ZN(_3829_));
 AOI21_X1 _6302_ (.A(_1321_),
    .B1(_1482_),
    .B2(_1483_),
    .ZN(_1507_));
 XNOR2_X1 _6303_ (.A(_3964_),
    .B(_1507_),
    .ZN(_3833_));
 NOR2_X1 _6304_ (.A1(_1495_),
    .A2(_3875_),
    .ZN(_1508_));
 XNOR2_X1 _6305_ (.A(_3900_),
    .B(_1508_),
    .ZN(_3837_));
 MUX2_X1 _6306_ (.A(_3844_),
    .B(_3717_),
    .S(_1321_),
    .Z(_2969_));
 INV_X1 _6307_ (.A(_2969_),
    .ZN(_2973_));
 INV_X1 _6308_ (.A(_3849_),
    .ZN(_1509_));
 AOI21_X1 _6309_ (.A(_3805_),
    .B1(_3811_),
    .B2(_3806_),
    .ZN(_1510_));
 BUF_X8 clone17 (.A(_0235_),
    .Z(net17));
 BUF_X2 _6311_ (.A(_3812_),
    .Z(_1512_));
 NAND2_X1 _6312_ (.A1(_3808_),
    .A2(_1512_),
    .ZN(_1513_));
 INV_X1 _6313_ (.A(_3815_),
    .ZN(_1514_));
 CLKBUF_X2 _6314_ (.A(_3816_),
    .Z(_1515_));
 INV_X1 _6315_ (.A(_3820_),
    .ZN(_1516_));
 INV_X1 _6316_ (.A(_3827_),
    .ZN(_1517_));
 INV_X1 _6317_ (.A(_3835_),
    .ZN(_1518_));
 INV_X1 _6318_ (.A(_3845_),
    .ZN(_1519_));
 INV_X1 _6319_ (.A(_3846_),
    .ZN(_1520_));
 OAI21_X1 _6320_ (.A(_1519_),
    .B1(_1520_),
    .B2(_2968_),
    .ZN(_1521_));
 AOI21_X1 _6321_ (.A(_3839_),
    .B1(_1521_),
    .B2(_3840_),
    .ZN(_1522_));
 INV_X1 _6322_ (.A(_3836_),
    .ZN(_1523_));
 OAI21_X1 _6323_ (.A(_1518_),
    .B1(_1522_),
    .B2(_1523_),
    .ZN(_1524_));
 AOI21_X2 _6324_ (.A(_3831_),
    .B1(_1524_),
    .B2(_3832_),
    .ZN(_1525_));
 INV_X1 _6325_ (.A(_3828_),
    .ZN(_1526_));
 OAI21_X1 _6326_ (.A(_1517_),
    .B1(_1525_),
    .B2(_1526_),
    .ZN(_1527_));
 AOI21_X2 _6327_ (.A(_3823_),
    .B1(_1527_),
    .B2(_3824_),
    .ZN(_1528_));
 NOR2_X1 _6328_ (.A1(_1516_),
    .A2(_1528_),
    .ZN(_1529_));
 OAI21_X1 _6329_ (.A(_1515_),
    .B1(_3819_),
    .B2(_1529_),
    .ZN(_1530_));
 AND2_X1 _6330_ (.A1(_1514_),
    .A2(_1530_),
    .ZN(_1531_));
 OAI21_X1 _6331_ (.A(_1510_),
    .B1(_1513_),
    .B2(_1531_),
    .ZN(_1532_));
 CLKBUF_X2 _6332_ (.A(_3854_),
    .Z(_1533_));
 AOI21_X1 _6333_ (.A(_3853_),
    .B1(_1532_),
    .B2(_1533_),
    .ZN(_1534_));
 INV_X1 _6334_ (.A(_3850_),
    .ZN(_1535_));
 OAI21_X1 _6335_ (.A(_1509_),
    .B1(_1534_),
    .B2(_1535_),
    .ZN(_1536_));
 XOR2_X2 _6336_ (.A(_3802_),
    .B(_1536_),
    .Z(_4015_));
 INV_X1 _6337_ (.A(_3805_),
    .ZN(_1537_));
 INV_X1 _6338_ (.A(_3823_),
    .ZN(_1538_));
 INV_X1 _6339_ (.A(_3831_),
    .ZN(_1539_));
 INV_X1 _6340_ (.A(_3839_),
    .ZN(_1540_));
 INV_X1 _6341_ (.A(_3840_),
    .ZN(_1541_));
 OAI21_X1 _6342_ (.A(_1540_),
    .B1(_1541_),
    .B2(_2970_),
    .ZN(_1542_));
 AOI21_X2 _6343_ (.A(_3835_),
    .B1(_1542_),
    .B2(_3836_),
    .ZN(_1543_));
 INV_X1 _6344_ (.A(_3832_),
    .ZN(_1544_));
 OAI21_X1 _6345_ (.A(_1539_),
    .B1(_1543_),
    .B2(_1544_),
    .ZN(_1545_));
 AOI21_X2 _6346_ (.A(_3827_),
    .B1(_1545_),
    .B2(_3828_),
    .ZN(_1546_));
 INV_X1 _6347_ (.A(_3824_),
    .ZN(_1547_));
 OAI21_X1 _6348_ (.A(_1538_),
    .B1(_1546_),
    .B2(_1547_),
    .ZN(_1548_));
 AOI21_X2 _6349_ (.A(_3819_),
    .B1(_1548_),
    .B2(_3820_),
    .ZN(_1549_));
 INV_X1 _6350_ (.A(_1515_),
    .ZN(_1550_));
 OAI21_X1 _6351_ (.A(_1514_),
    .B1(_1549_),
    .B2(_1550_),
    .ZN(_1551_));
 AOI21_X2 _6352_ (.A(_3811_),
    .B1(_1551_),
    .B2(_1512_),
    .ZN(_1552_));
 INV_X1 _6353_ (.A(net138),
    .ZN(_1553_));
 OAI21_X1 _6354_ (.A(_1537_),
    .B1(_1552_),
    .B2(_1553_),
    .ZN(_1554_));
 AOI21_X2 _6355_ (.A(_3853_),
    .B1(_1554_),
    .B2(_1533_),
    .ZN(_1555_));
 XNOR2_X2 _6356_ (.A(_3850_),
    .B(_1555_),
    .ZN(_4019_));
 NAND4_X1 _6357_ (.A1(_1515_),
    .A2(_3808_),
    .A3(_1512_),
    .A4(_1529_),
    .ZN(_1556_));
 INV_X1 _6358_ (.A(_1512_),
    .ZN(_1557_));
 AOI21_X1 _6359_ (.A(_3815_),
    .B1(_3819_),
    .B2(_1515_),
    .ZN(_1558_));
 NOR2_X1 _6360_ (.A1(_1557_),
    .A2(_1558_),
    .ZN(_1559_));
 OAI21_X1 _6361_ (.A(_3806_),
    .B1(_3811_),
    .B2(_1559_),
    .ZN(_1560_));
 NAND3_X2 _6362_ (.A1(_1556_),
    .A2(_1537_),
    .A3(_1560_),
    .ZN(_1561_));
 XOR2_X2 _6363_ (.A(_1533_),
    .B(_1561_),
    .Z(_4023_));
 XNOR2_X2 _6364_ (.A(net138),
    .B(_1552_),
    .ZN(_3977_));
 XNOR2_X2 _6365_ (.A(_1512_),
    .B(_1531_),
    .ZN(_4027_));
 XNOR2_X2 _6366_ (.A(_3820_),
    .B(_1528_),
    .ZN(_3985_));
 INV_X1 _6367_ (.A(_3985_),
    .ZN(_3926_));
 XNOR2_X2 _6368_ (.A(_3824_),
    .B(_1546_),
    .ZN(_3990_));
 INV_X1 _6369_ (.A(_3990_),
    .ZN(_3927_));
 INV_X1 _6370_ (.A(_3857_),
    .ZN(_1562_));
 INV_X1 _6371_ (.A(_3863_),
    .ZN(_1563_));
 INV_X1 _6372_ (.A(_3869_),
    .ZN(_1564_));
 INV_X1 _6373_ (.A(_3876_),
    .ZN(_1565_));
 INV_X1 _6374_ (.A(_3882_),
    .ZN(_1566_));
 INV_X1 _6375_ (.A(_3888_),
    .ZN(_1567_));
 INV_X1 _6376_ (.A(_3894_),
    .ZN(_1568_));
 BUF_X1 _6377_ (.A(_3898_),
    .Z(_1569_));
 AOI21_X1 _6378_ (.A(_3897_),
    .B1(_1569_),
    .B2(_2940_),
    .ZN(_1570_));
 INV_X2 _6379_ (.A(_3895_),
    .ZN(_1571_));
 OAI21_X4 _6380_ (.A(_1568_),
    .B1(_1571_),
    .B2(_1570_),
    .ZN(_1572_));
 AOI21_X4 _6381_ (.A(_3891_),
    .B1(_3892_),
    .B2(_1572_),
    .ZN(_1573_));
 INV_X1 _6382_ (.A(_3889_),
    .ZN(_1574_));
 OAI21_X4 _6383_ (.A(_1567_),
    .B1(_1573_),
    .B2(_1574_),
    .ZN(_1575_));
 AOI21_X4 _6384_ (.A(_3885_),
    .B1(_3886_),
    .B2(_1575_),
    .ZN(_1576_));
 INV_X1 _6385_ (.A(_3883_),
    .ZN(_1577_));
 OAI21_X4 _6386_ (.A(_1566_),
    .B1(_1576_),
    .B2(_1577_),
    .ZN(_1578_));
 AOI21_X4 _6387_ (.A(_3879_),
    .B1(_3880_),
    .B2(_1578_),
    .ZN(_1579_));
 INV_X1 _6388_ (.A(_3877_),
    .ZN(_1580_));
 OAI21_X4 _6389_ (.A(_1565_),
    .B1(_1579_),
    .B2(_1580_),
    .ZN(_1581_));
 AOI21_X4 _6390_ (.A(_3872_),
    .B1(_3873_),
    .B2(_1581_),
    .ZN(_1582_));
 INV_X1 _6391_ (.A(_3870_),
    .ZN(_1583_));
 OAI21_X4 _6392_ (.A(_1564_),
    .B1(_1582_),
    .B2(_1583_),
    .ZN(_1584_));
 AOI21_X4 _6393_ (.A(_3866_),
    .B1(_1584_),
    .B2(_3867_),
    .ZN(_1585_));
 INV_X1 _6394_ (.A(_3864_),
    .ZN(_1586_));
 OAI21_X4 _6395_ (.A(_1563_),
    .B1(_1585_),
    .B2(_1586_),
    .ZN(_1587_));
 AOI21_X4 _6396_ (.A(_3860_),
    .B1(_1587_),
    .B2(_3861_),
    .ZN(_1588_));
 INV_X2 _6397_ (.A(_3858_),
    .ZN(_1589_));
 OAI21_X4 _6398_ (.A(_1562_),
    .B1(_1589_),
    .B2(_1588_),
    .ZN(_1590_));
 INV_X8 _6399_ (.A(_1590_),
    .ZN(_1591_));
 BUF_X16 _6400_ (.A(_1591_),
    .Z(_4053_));
 INV_X1 _6401_ (.A(_3719_),
    .ZN(_1592_));
 INV_X1 _6402_ (.A(_3726_),
    .ZN(_1593_));
 INV_X1 _6403_ (.A(_3734_),
    .ZN(_1594_));
 AOI21_X1 _6404_ (.A(_3740_),
    .B1(_3741_),
    .B2(_2964_),
    .ZN(_1595_));
 INV_X1 _6405_ (.A(_3735_),
    .ZN(_1596_));
 OAI21_X2 _6406_ (.A(_1594_),
    .B1(_1595_),
    .B2(_1596_),
    .ZN(_1597_));
 AOI21_X1 _6407_ (.A(_3730_),
    .B1(_1597_),
    .B2(_3731_),
    .ZN(_1598_));
 INV_X1 _6408_ (.A(_3727_),
    .ZN(_1599_));
 OAI21_X2 _6409_ (.A(_1593_),
    .B1(_1598_),
    .B2(_1599_),
    .ZN(_1600_));
 AOI21_X1 _6410_ (.A(_3722_),
    .B1(_1600_),
    .B2(_3723_),
    .ZN(_1601_));
 INV_X1 _6411_ (.A(_3720_),
    .ZN(_1602_));
 OAI21_X2 _6412_ (.A(_1592_),
    .B1(_1601_),
    .B2(_1602_),
    .ZN(_1603_));
 XNOR2_X2 _6413_ (.A(_3902_),
    .B(_1603_),
    .ZN(_4009_));
 XNOR2_X2 _6414_ (.A(_1515_),
    .B(_1549_),
    .ZN(_3981_));
 INV_X1 _6415_ (.A(_3908_),
    .ZN(_1604_));
 INV_X1 _6416_ (.A(_3916_),
    .ZN(_1605_));
 INV_X1 _6417_ (.A(_3924_),
    .ZN(_1606_));
 AOI21_X2 _6418_ (.A(_3930_),
    .B1(_2974_),
    .B2(_3931_),
    .ZN(_1607_));
 INV_X1 _6419_ (.A(_3925_),
    .ZN(_1608_));
 OAI21_X4 _6420_ (.A(_1606_),
    .B1(_1608_),
    .B2(_1607_),
    .ZN(_1609_));
 AOI21_X4 _6421_ (.A(_3920_),
    .B1(_1609_),
    .B2(_3921_),
    .ZN(_1610_));
 INV_X1 _6422_ (.A(_3917_),
    .ZN(_1611_));
 OAI21_X4 _6423_ (.A(_1605_),
    .B1(_1611_),
    .B2(_1610_),
    .ZN(_1612_));
 AOI21_X4 _6424_ (.A(_3912_),
    .B1(_3913_),
    .B2(_1612_),
    .ZN(_1613_));
 INV_X1 _6425_ (.A(_3909_),
    .ZN(_1614_));
 OAI21_X4 _6426_ (.A(_1604_),
    .B1(_1613_),
    .B2(_1614_),
    .ZN(_1615_));
 XNOR2_X2 _6427_ (.A(_3906_),
    .B(_1615_),
    .ZN(_4172_));
 INV_X1 _6428_ (.A(_4172_),
    .ZN(_3933_));
 AOI21_X1 _6429_ (.A(_1370_),
    .B1(_1379_),
    .B2(_1241_),
    .ZN(_3936_));
 BUF_X2 _6430_ (.A(_3938_),
    .Z(_1616_));
 INV_X1 _6431_ (.A(_3759_),
    .ZN(_1617_));
 INV_X1 _6432_ (.A(_1393_),
    .ZN(_1618_));
 OAI21_X1 _6433_ (.A(_1617_),
    .B1(_1494_),
    .B2(_1618_),
    .ZN(_1619_));
 AOI21_X1 _6434_ (.A(_3755_),
    .B1(_1619_),
    .B2(_3756_),
    .ZN(_1620_));
 XOR2_X2 _6435_ (.A(_1616_),
    .B(_1620_),
    .Z(_1621_));
 INV_X1 _6436_ (.A(_1621_),
    .ZN(_3939_));
 AOI21_X1 _6437_ (.A(_1492_),
    .B1(_1497_),
    .B2(_1498_),
    .ZN(_3940_));
 INV_X1 _6438_ (.A(_3949_),
    .ZN(_1622_));
 INV_X1 _6439_ (.A(_3971_),
    .ZN(_1623_));
 INV_X1 _6440_ (.A(_3961_),
    .ZN(_1624_));
 INV_X1 _6441_ (.A(_3901_),
    .ZN(_1625_));
 AOI21_X1 _6442_ (.A(_3719_),
    .B1(_1347_),
    .B2(_3720_),
    .ZN(_1626_));
 INV_X1 _6443_ (.A(_3902_),
    .ZN(_1627_));
 OAI21_X2 _6444_ (.A(_1625_),
    .B1(_1626_),
    .B2(_1627_),
    .ZN(_1628_));
 AOI21_X1 _6445_ (.A(_3965_),
    .B1(_1628_),
    .B2(_3966_),
    .ZN(_1629_));
 INV_X1 _6446_ (.A(_3962_),
    .ZN(_1630_));
 OAI21_X2 _6447_ (.A(_1624_),
    .B1(_1629_),
    .B2(_1630_),
    .ZN(_1631_));
 AOI21_X1 _6448_ (.A(_3957_),
    .B1(_1631_),
    .B2(_3958_),
    .ZN(_1632_));
 INV_X1 _6449_ (.A(_3972_),
    .ZN(_1633_));
 OAI21_X2 _6450_ (.A(_1623_),
    .B1(_1632_),
    .B2(_1633_),
    .ZN(_1634_));
 AOI21_X1 _6451_ (.A(_3953_),
    .B1(_1634_),
    .B2(_3968_),
    .ZN(_1635_));
 INV_X1 _6452_ (.A(_3950_),
    .ZN(_1636_));
 OAI21_X2 _6453_ (.A(_1622_),
    .B1(_1635_),
    .B2(_1636_),
    .ZN(_1637_));
 XNOR2_X2 _6454_ (.A(_3946_),
    .B(_1637_),
    .ZN(_1638_));
 INV_X1 _6455_ (.A(_1638_),
    .ZN(_4112_));
 INV_X1 _6456_ (.A(_3953_),
    .ZN(_1639_));
 INV_X1 _6457_ (.A(_3957_),
    .ZN(_1640_));
 INV_X1 _6458_ (.A(_3965_),
    .ZN(_1641_));
 AOI21_X2 _6459_ (.A(_3901_),
    .B1(_1603_),
    .B2(_3902_),
    .ZN(_1642_));
 INV_X2 _6460_ (.A(_3966_),
    .ZN(_1643_));
 OAI21_X4 _6461_ (.A(_1641_),
    .B1(_1642_),
    .B2(_1643_),
    .ZN(_1644_));
 AOI21_X2 _6462_ (.A(_3961_),
    .B1(_1644_),
    .B2(_3962_),
    .ZN(_1645_));
 INV_X2 _6463_ (.A(_3958_),
    .ZN(_1646_));
 OAI21_X4 _6464_ (.A(_1640_),
    .B1(_1645_),
    .B2(_1646_),
    .ZN(_1647_));
 AOI21_X4 _6465_ (.A(_3971_),
    .B1(_1647_),
    .B2(_3972_),
    .ZN(_1648_));
 INV_X1 _6466_ (.A(_3954_),
    .ZN(_1649_));
 OAI21_X4 _6467_ (.A(_1639_),
    .B1(_1649_),
    .B2(_1648_),
    .ZN(_1650_));
 XNOR2_X2 _6468_ (.A(_3950_),
    .B(_1650_),
    .ZN(_1651_));
 INV_X1 _6469_ (.A(_1651_),
    .ZN(_4128_));
 XNOR2_X2 _6470_ (.A(_3968_),
    .B(_1634_),
    .ZN(_1652_));
 INV_X1 _6471_ (.A(_1652_),
    .ZN(_4116_));
 XNOR2_X2 _6472_ (.A(_1633_),
    .B(_1647_),
    .ZN(_4134_));
 XNOR2_X2 _6473_ (.A(_1646_),
    .B(_1631_),
    .ZN(_4120_));
 XNOR2_X2 _6474_ (.A(_3962_),
    .B(_1644_),
    .ZN(_1653_));
 INV_X1 _6475_ (.A(_1653_),
    .ZN(_4124_));
 OAI21_X1 _6476_ (.A(_1509_),
    .B1(_1555_),
    .B2(_1535_),
    .ZN(_1654_));
 AOI21_X2 _6477_ (.A(_3801_),
    .B1(_1654_),
    .B2(_3802_),
    .ZN(_1655_));
 XNOR2_X2 _6478_ (.A(_3942_),
    .B(_1655_),
    .ZN(_3974_));
 XNOR2_X2 _6479_ (.A(_3966_),
    .B(_1628_),
    .ZN(_1656_));
 INV_X2 _6480_ (.A(_1656_),
    .ZN(_4075_));
 BUF_X8 _6481_ (.A(_1590_),
    .Z(_1657_));
 BUF_X16 _6482_ (.A(_1657_),
    .Z(_4031_));
 NAND3_X1 _6483_ (.A1(_4011_),
    .A2(_1653_),
    .A3(_1656_),
    .ZN(_1658_));
 NOR3_X1 _6484_ (.A1(_4134_),
    .A2(_4120_),
    .A3(_1658_),
    .ZN(_1659_));
 NAND3_X1 _6485_ (.A1(_1651_),
    .A2(_1652_),
    .A3(_1659_),
    .ZN(_1660_));
 OAI21_X1 _6486_ (.A(net4),
    .B1(_4112_),
    .B2(_1660_),
    .ZN(_1661_));
 AOI21_X1 _6487_ (.A(_3759_),
    .B1(_3625_),
    .B2(_1393_),
    .ZN(_1662_));
 NAND2_X1 _6488_ (.A1(_3626_),
    .A2(_1393_),
    .ZN(_1663_));
 OAI21_X1 _6489_ (.A(_1662_),
    .B1(_1663_),
    .B2(_1284_),
    .ZN(_1664_));
 AND2_X1 _6490_ (.A1(_3756_),
    .A2(_1616_),
    .ZN(_1665_));
 AOI221_X2 _6491_ (.A(_3937_),
    .B1(_1664_),
    .B2(_1665_),
    .C1(_3755_),
    .C2(_1616_),
    .ZN(_1666_));
 OAI21_X2 _6492_ (.A(_1666_),
    .B1(_1458_),
    .B2(_1456_),
    .ZN(_1667_));
 AOI21_X1 _6493_ (.A(_3937_),
    .B1(_3755_),
    .B2(_1616_),
    .ZN(_1668_));
 NAND2_X1 _6494_ (.A1(_3756_),
    .A2(_1616_),
    .ZN(_1669_));
 OAI21_X4 _6495_ (.A(_1668_),
    .B1(_1669_),
    .B2(_1395_),
    .ZN(_1670_));
 NAND3_X4 _6496_ (.A1(_1670_),
    .A2(_1461_),
    .A3(_1460_),
    .ZN(_1671_));
 OAI211_X4 _6497_ (.A(_1667_),
    .B(_1671_),
    .C1(_1366_),
    .C2(_1370_),
    .ZN(_1672_));
 AND2_X1 _6498_ (.A1(_1129_),
    .A2(_1143_),
    .ZN(_1673_));
 AOI21_X2 _6499_ (.A(_0900_),
    .B1(_1113_),
    .B2(_1673_),
    .ZN(_1674_));
 OAI21_X1 _6500_ (.A(_1674_),
    .B1(_1368_),
    .B2(_1369_),
    .ZN(_1675_));
 AOI21_X2 _6501_ (.A(_1670_),
    .B1(_1461_),
    .B2(_1460_),
    .ZN(_1676_));
 NOR3_X1 _6502_ (.A1(_1456_),
    .A2(_1458_),
    .A3(_1666_),
    .ZN(_1677_));
 OAI221_X4 _6503_ (.A(_1675_),
    .B1(_1676_),
    .B2(_1677_),
    .C1(_1241_),
    .C2(_3670_),
    .ZN(_1678_));
 NOR3_X2 _6504_ (.A1(_3818_),
    .A2(_3822_),
    .A3(_3826_),
    .ZN(_1679_));
 NOR3_X2 _6505_ (.A1(_3810_),
    .A2(_3814_),
    .A3(_3804_),
    .ZN(_1680_));
 NAND2_X1 _6506_ (.A1(_1679_),
    .A2(_1680_),
    .ZN(_1681_));
 OR2_X1 _6507_ (.A1(_3852_),
    .A2(_1681_),
    .ZN(_1682_));
 NOR3_X4 _6508_ (.A1(_3799_),
    .A2(_3847_),
    .A3(_1682_),
    .ZN(_1683_));
 AOI21_X4 _6509_ (.A(_1320_),
    .B1(_1621_),
    .B2(_1683_),
    .ZN(_1684_));
 AND3_X2 _6510_ (.A1(_1672_),
    .A2(_1678_),
    .A3(_1684_),
    .ZN(_1685_));
 AOI21_X4 _6511_ (.A(net1),
    .B1(_1672_),
    .B2(_1678_),
    .ZN(_1686_));
 INV_X1 _6512_ (.A(_3945_),
    .ZN(_1687_));
 AND2_X4 _6513_ (.A1(_3950_),
    .A2(_1650_),
    .ZN(_1688_));
 OAI21_X4 _6514_ (.A(_3946_),
    .B1(_3949_),
    .B2(_1688_),
    .ZN(_1689_));
 AND2_X4 _6515_ (.A1(_1687_),
    .A2(_1689_),
    .ZN(_1690_));
 AOI21_X4 _6516_ (.A(_1690_),
    .B1(_1481_),
    .B2(_1475_),
    .ZN(_1691_));
 NAND2_X4 _6517_ (.A1(_1687_),
    .A2(_1689_),
    .ZN(_1692_));
 NOR3_X4 _6518_ (.A1(_1491_),
    .A2(_1692_),
    .A3(_1490_),
    .ZN(_1693_));
 OAI22_X4 _6519_ (.A1(_1685_),
    .A2(_1686_),
    .B1(_1691_),
    .B2(_1693_),
    .ZN(_1694_));
 NAND3_X4 _6520_ (.A1(_1672_),
    .A2(_1678_),
    .A3(_1684_),
    .ZN(_1695_));
 NAND3_X1 _6521_ (.A1(net219),
    .A2(_1230_),
    .A3(_1240_),
    .ZN(_1696_));
 AOI211_X4 _6522_ (.A(_1676_),
    .B(_1677_),
    .C1(_1675_),
    .C2(_1696_),
    .ZN(_1697_));
 AOI221_X2 _6523_ (.A(_1370_),
    .B1(_1667_),
    .B2(_1671_),
    .C1(_1241_),
    .C2(_1674_),
    .ZN(_1698_));
 OAI21_X4 _6524_ (.A(_1320_),
    .B1(_1697_),
    .B2(net125),
    .ZN(_1699_));
 OAI21_X4 _6525_ (.A(_1692_),
    .B1(_1491_),
    .B2(_1490_),
    .ZN(_1700_));
 NAND3_X4 _6526_ (.A1(_1475_),
    .A2(_1481_),
    .A3(_1690_),
    .ZN(_1701_));
 NAND4_X4 _6527_ (.A1(_1695_),
    .A2(_1699_),
    .A3(_1700_),
    .A4(_1701_),
    .ZN(_1702_));
 NAND2_X4 _6528_ (.A1(_1694_),
    .A2(_1702_),
    .ZN(_1703_));
 MUX2_X1 _6529_ (.A(net221),
    .B(_1661_),
    .S(_1703_),
    .Z(_3973_));
 AOI22_X4 _6530_ (.A1(_1695_),
    .A2(_1699_),
    .B1(_1700_),
    .B2(_1701_),
    .ZN(_1704_));
 NOR4_X4 _6531_ (.A1(_1691_),
    .A2(_1686_),
    .A3(_1685_),
    .A4(_1693_),
    .ZN(_1705_));
 NOR3_X4 _6532_ (.A1(_1590_),
    .A2(_1704_),
    .A3(_1705_),
    .ZN(_1706_));
 INV_X1 _6533_ (.A(_4134_),
    .ZN(_1707_));
 NAND2_X1 _6534_ (.A1(_4010_),
    .A2(_4009_),
    .ZN(_1708_));
 NOR4_X2 _6535_ (.A1(_4120_),
    .A2(_4124_),
    .A3(_4075_),
    .A4(_1708_),
    .ZN(_1709_));
 NAND3_X2 _6536_ (.A1(_1652_),
    .A2(_1707_),
    .A3(_1709_),
    .ZN(_1710_));
 NAND2_X1 _6537_ (.A1(_1638_),
    .A2(_1651_),
    .ZN(_1711_));
 OAI21_X4 _6538_ (.A(net4),
    .B1(_1710_),
    .B2(_1711_),
    .ZN(_1712_));
 AOI21_X4 _6539_ (.A(_1712_),
    .B1(_1702_),
    .B2(_1694_),
    .ZN(_1713_));
 NOR2_X1 _6540_ (.A1(_1706_),
    .A2(_1713_),
    .ZN(_4016_));
 MUX2_X1 _6541_ (.A(net221),
    .B(_1661_),
    .S(_1703_),
    .Z(_4020_));
 NOR2_X1 _6542_ (.A1(_1706_),
    .A2(_1713_),
    .ZN(_4024_));
 MUX2_X1 _6543_ (.A(net221),
    .B(_1661_),
    .S(_1703_),
    .Z(_3978_));
 XNOR2_X2 _6544_ (.A(_1703_),
    .B(_1712_),
    .ZN(_4028_));
 NAND2_X1 _6545_ (.A1(net225),
    .A2(_1660_),
    .ZN(_1714_));
 XNOR2_X1 _6546_ (.A(_1638_),
    .B(_1714_),
    .ZN(_3982_));
 NAND2_X1 _6547_ (.A1(net225),
    .A2(_1710_),
    .ZN(_1715_));
 XNOR2_X1 _6548_ (.A(_1651_),
    .B(_1715_),
    .ZN(_3986_));
 NOR2_X1 _6549_ (.A1(_4053_),
    .A2(_1659_),
    .ZN(_1716_));
 XNOR2_X1 _6550_ (.A(_4116_),
    .B(_1716_),
    .ZN(_3989_));
 NOR2_X1 _6551_ (.A1(_4053_),
    .A2(_1709_),
    .ZN(_1717_));
 XNOR2_X1 _6552_ (.A(_4134_),
    .B(_1717_),
    .ZN(_3993_));
 NAND2_X1 _6553_ (.A1(_1657_),
    .A2(_1658_),
    .ZN(_1718_));
 XOR2_X1 _6554_ (.A(_4120_),
    .B(_1718_),
    .Z(_3997_));
 OAI21_X1 _6555_ (.A(_1657_),
    .B1(_4075_),
    .B2(_1708_),
    .ZN(_1719_));
 XNOR2_X1 _6556_ (.A(_1653_),
    .B(_1719_),
    .ZN(_4002_));
 NOR2_X4 _6557_ (.A1(_4011_),
    .A2(_4053_),
    .ZN(_1720_));
 XNOR2_X2 _6558_ (.A(_4075_),
    .B(_1720_),
    .ZN(_4005_));
 NOR2_X4 _6559_ (.A1(_4009_),
    .A2(_4031_),
    .ZN(_1721_));
 AOI21_X4 _6560_ (.A(_1721_),
    .B1(_4031_),
    .B2(_4012_),
    .ZN(_2979_));
 INV_X1 _6561_ (.A(_4017_),
    .ZN(_1722_));
 INV_X1 _6562_ (.A(_4025_),
    .ZN(_1723_));
 INV_X1 _6563_ (.A(_4029_),
    .ZN(_1724_));
 INV_X1 _6564_ (.A(_3987_),
    .ZN(_1725_));
 INV_X1 _6565_ (.A(_3995_),
    .ZN(_1726_));
 INV_X1 _6566_ (.A(_4003_),
    .ZN(_1727_));
 AOI21_X2 _6567_ (.A(_4007_),
    .B1(_4008_),
    .B2(_2981_),
    .ZN(_1728_));
 INV_X1 _6568_ (.A(_4004_),
    .ZN(_1729_));
 OAI21_X2 _6569_ (.A(_1727_),
    .B1(_1728_),
    .B2(_1729_),
    .ZN(_1730_));
 AOI21_X2 _6570_ (.A(_3999_),
    .B1(_1730_),
    .B2(_4000_),
    .ZN(_1731_));
 INV_X1 _6571_ (.A(_3996_),
    .ZN(_1732_));
 OAI21_X2 _6572_ (.A(_1726_),
    .B1(_1731_),
    .B2(_1732_),
    .ZN(_1733_));
 AOI21_X2 _6573_ (.A(_3991_),
    .B1(_1733_),
    .B2(_3992_),
    .ZN(_1734_));
 INV_X1 _6574_ (.A(_3988_),
    .ZN(_1735_));
 OAI21_X2 _6575_ (.A(_1725_),
    .B1(_1734_),
    .B2(_1735_),
    .ZN(_1736_));
 AOI21_X2 _6576_ (.A(_3983_),
    .B1(_1736_),
    .B2(_3984_),
    .ZN(_1737_));
 INV_X2 _6577_ (.A(_4030_),
    .ZN(_1738_));
 OAI21_X2 _6578_ (.A(_1724_),
    .B1(_1737_),
    .B2(_1738_),
    .ZN(_1739_));
 AOI21_X1 _6579_ (.A(_3979_),
    .B1(_1739_),
    .B2(net163),
    .ZN(_1740_));
 INV_X1 _6580_ (.A(_4026_),
    .ZN(_1741_));
 OAI21_X2 _6581_ (.A(_1723_),
    .B1(_1740_),
    .B2(_1741_),
    .ZN(_1742_));
 AOI21_X1 _6582_ (.A(_4021_),
    .B1(_1742_),
    .B2(_4022_),
    .ZN(_1743_));
 INV_X1 _6583_ (.A(_4018_),
    .ZN(_1744_));
 OAI21_X1 _6584_ (.A(_1722_),
    .B1(_1743_),
    .B2(_1744_),
    .ZN(_1745_));
 XNOR2_X1 _6585_ (.A(_3976_),
    .B(_1745_),
    .ZN(_1746_));
 INV_X1 _6586_ (.A(_1746_),
    .ZN(_4139_));
 INV_X1 _6587_ (.A(_2983_),
    .ZN(_2980_));
 INV_X1 _6588_ (.A(_4013_),
    .ZN(_1747_));
 INV_X2 _6589_ (.A(_4014_),
    .ZN(_1748_));
 OAI21_X4 _6590_ (.A(_1747_),
    .B1(_2983_),
    .B2(_1748_),
    .ZN(_1749_));
 AOI21_X4 _6591_ (.A(_4007_),
    .B1(_1749_),
    .B2(_4008_),
    .ZN(_1750_));
 OAI21_X4 _6592_ (.A(_1727_),
    .B1(_1750_),
    .B2(_1729_),
    .ZN(_1751_));
 AOI21_X4 _6593_ (.A(_3999_),
    .B1(_4000_),
    .B2(_1751_),
    .ZN(_1752_));
 OAI21_X4 _6594_ (.A(_1726_),
    .B1(_1752_),
    .B2(_1732_),
    .ZN(_1753_));
 AOI21_X4 _6595_ (.A(_3991_),
    .B1(_1753_),
    .B2(_3992_),
    .ZN(_1754_));
 OAI21_X4 _6596_ (.A(_1725_),
    .B1(_1754_),
    .B2(_1735_),
    .ZN(_1755_));
 AOI21_X4 _6597_ (.A(_3983_),
    .B1(_1755_),
    .B2(_3984_),
    .ZN(_1756_));
 OAI21_X4 _6598_ (.A(_1724_),
    .B1(_1738_),
    .B2(_1756_),
    .ZN(_1757_));
 AOI21_X4 _6599_ (.A(_3979_),
    .B1(_1757_),
    .B2(_3980_),
    .ZN(_1758_));
 OAI21_X4 _6600_ (.A(_1723_),
    .B1(_1741_),
    .B2(_1758_),
    .ZN(_1759_));
 AOI21_X4 _6601_ (.A(_4021_),
    .B1(_1759_),
    .B2(_4022_),
    .ZN(_1760_));
 XNOR2_X2 _6602_ (.A(_4018_),
    .B(_1760_),
    .ZN(_4179_));
 XOR2_X2 _6603_ (.A(_4022_),
    .B(_1742_),
    .Z(_4183_));
 XNOR2_X2 _6604_ (.A(_4026_),
    .B(_1758_),
    .ZN(_4186_));
 XOR2_X2 _6605_ (.A(net164),
    .B(_1739_),
    .Z(_4142_));
 XNOR2_X2 _6606_ (.A(_4030_),
    .B(_1756_),
    .ZN(_4190_));
 XOR2_X2 _6607_ (.A(_3984_),
    .B(_1736_),
    .Z(_4146_));
 XNOR2_X2 _6608_ (.A(_3988_),
    .B(_1754_),
    .ZN(_4194_));
 INV_X1 _6609_ (.A(_4033_),
    .ZN(_1761_));
 INV_X1 _6610_ (.A(_4039_),
    .ZN(_1762_));
 INV_X1 _6611_ (.A(_4045_),
    .ZN(_1763_));
 INV_X1 _6612_ (.A(_4051_),
    .ZN(_1764_));
 INV_X1 _6613_ (.A(_4058_),
    .ZN(_1765_));
 INV_X1 _6614_ (.A(_4064_),
    .ZN(_1766_));
 INV_X1 _6615_ (.A(_4070_),
    .ZN(_1767_));
 BUF_X2 clone3 (.A(_1790_),
    .Z(net3));
 BUF_X4 _6617_ (.A(_0005_),
    .Z(_1769_));
 AOI21_X2 _6618_ (.A(_4073_),
    .B1(_4074_),
    .B2(_1769_),
    .ZN(_1770_));
 INV_X2 _6619_ (.A(_4071_),
    .ZN(_1771_));
 OAI21_X4 _6620_ (.A(_1767_),
    .B1(_1771_),
    .B2(_1770_),
    .ZN(_1772_));
 AOI21_X4 _6621_ (.A(_4067_),
    .B1(_1772_),
    .B2(_4068_),
    .ZN(_1773_));
 INV_X1 _6622_ (.A(_4065_),
    .ZN(_1774_));
 OAI21_X4 _6623_ (.A(_1766_),
    .B1(_1774_),
    .B2(_1773_),
    .ZN(_1775_));
 AOI21_X4 _6624_ (.A(_4061_),
    .B1(_1775_),
    .B2(_4062_),
    .ZN(_1776_));
 INV_X1 _6625_ (.A(_4059_),
    .ZN(_1777_));
 OAI21_X4 _6626_ (.A(_1765_),
    .B1(_1776_),
    .B2(_1777_),
    .ZN(_1778_));
 AOI21_X4 _6627_ (.A(_4055_),
    .B1(_1778_),
    .B2(_4056_),
    .ZN(_1779_));
 INV_X1 _6628_ (.A(_4052_),
    .ZN(_1780_));
 OAI21_X4 _6629_ (.A(_1764_),
    .B1(_1779_),
    .B2(_1780_),
    .ZN(_1781_));
 AOI21_X4 _6630_ (.A(_4048_),
    .B1(_1781_),
    .B2(_4049_),
    .ZN(_1782_));
 INV_X1 _6631_ (.A(_4046_),
    .ZN(_1783_));
 OAI21_X4 _6632_ (.A(_1763_),
    .B1(_1782_),
    .B2(_1783_),
    .ZN(_1784_));
 AOI21_X4 _6633_ (.A(_4042_),
    .B1(_4043_),
    .B2(_1784_),
    .ZN(_1785_));
 INV_X1 _6634_ (.A(_4040_),
    .ZN(_1786_));
 OAI21_X4 _6635_ (.A(_1762_),
    .B1(_1785_),
    .B2(_1786_),
    .ZN(_1787_));
 AOI21_X4 _6636_ (.A(_4036_),
    .B1(_1787_),
    .B2(_4037_),
    .ZN(_1788_));
 INV_X1 _6637_ (.A(_4034_),
    .ZN(_1789_));
 OAI21_X4 _6638_ (.A(_1761_),
    .B1(_1788_),
    .B2(_1789_),
    .ZN(_1790_));
 BUF_X8 _6639_ (.A(_1790_),
    .Z(_1791_));
 INV_X8 _6640_ (.A(_1791_),
    .ZN(_4223_));
 INV_X1 _6641_ (.A(_3905_),
    .ZN(_1792_));
 INV_X1 _6642_ (.A(_3912_),
    .ZN(_1793_));
 INV_X1 _6643_ (.A(_3920_),
    .ZN(_1794_));
 AOI21_X1 _6644_ (.A(_3924_),
    .B1(_2976_),
    .B2(_3925_),
    .ZN(_1795_));
 INV_X1 _6645_ (.A(_3921_),
    .ZN(_1796_));
 OAI21_X1 _6646_ (.A(_1794_),
    .B1(_1795_),
    .B2(_1796_),
    .ZN(_1797_));
 AOI21_X1 _6647_ (.A(_3916_),
    .B1(_1797_),
    .B2(_3917_),
    .ZN(_1798_));
 INV_X1 _6648_ (.A(_3913_),
    .ZN(_1799_));
 OAI21_X1 _6649_ (.A(_1793_),
    .B1(_1798_),
    .B2(_1799_),
    .ZN(_1800_));
 AOI21_X2 _6650_ (.A(_3908_),
    .B1(_1800_),
    .B2(_3909_),
    .ZN(_1801_));
 INV_X1 _6651_ (.A(_3906_),
    .ZN(_1802_));
 OAI21_X2 _6652_ (.A(_1792_),
    .B1(_1801_),
    .B2(_1802_),
    .ZN(_1803_));
 XNOR2_X2 _6653_ (.A(net144),
    .B(_1803_),
    .ZN(_4173_));
 INV_X1 _6654_ (.A(_4173_),
    .ZN(_4080_));
 INV_X1 _6655_ (.A(_4194_),
    .ZN(_4104_));
 INV_X1 _6656_ (.A(_4146_),
    .ZN(_4103_));
 INV_X1 _6657_ (.A(_4249_),
    .ZN(_1804_));
 INV_X1 _6658_ (.A(_4089_),
    .ZN(_1805_));
 INV_X1 _6659_ (.A(_4097_),
    .ZN(_1806_));
 AOI21_X1 _6660_ (.A(_4101_),
    .B1(_4102_),
    .B2(_2986_),
    .ZN(_1807_));
 INV_X1 _6661_ (.A(_4098_),
    .ZN(_1808_));
 OAI21_X1 _6662_ (.A(_1806_),
    .B1(_1807_),
    .B2(_1808_),
    .ZN(_1809_));
 AOI21_X1 _6663_ (.A(_4093_),
    .B1(_1809_),
    .B2(_4094_),
    .ZN(_1810_));
 INV_X1 _6664_ (.A(_4090_),
    .ZN(_1811_));
 OAI21_X1 _6665_ (.A(_1805_),
    .B1(_1810_),
    .B2(_1811_),
    .ZN(_1812_));
 AOI21_X1 _6666_ (.A(_4085_),
    .B1(_1812_),
    .B2(_4086_),
    .ZN(_1813_));
 INV_X1 _6667_ (.A(_4250_),
    .ZN(_1814_));
 OAI21_X2 _6668_ (.A(_1804_),
    .B1(_1813_),
    .B2(_1814_),
    .ZN(_1815_));
 XOR2_X2 _6669_ (.A(_4082_),
    .B(_1815_),
    .Z(_4110_));
 INV_X1 _6670_ (.A(_4110_),
    .ZN(_4278_));
 INV_X1 _6671_ (.A(_4136_),
    .ZN(_1816_));
 INV_X1 _6672_ (.A(_4126_),
    .ZN(_1817_));
 AOI21_X2 _6673_ (.A(_4077_),
    .B1(_1803_),
    .B2(_4078_),
    .ZN(_1818_));
 INV_X2 _6674_ (.A(_4127_),
    .ZN(_1819_));
 OAI21_X4 _6675_ (.A(_1817_),
    .B1(_1818_),
    .B2(_1819_),
    .ZN(_1820_));
 AOI21_X2 _6676_ (.A(_4122_),
    .B1(_1820_),
    .B2(net232),
    .ZN(_1821_));
 INV_X1 _6677_ (.A(_4137_),
    .ZN(_1822_));
 OAI21_X2 _6678_ (.A(_1816_),
    .B1(_1821_),
    .B2(_1822_),
    .ZN(_1823_));
 AOI21_X1 _6679_ (.A(_4118_),
    .B1(_1823_),
    .B2(_4133_),
    .ZN(_1824_));
 INV_X1 _6680_ (.A(_1824_),
    .ZN(_1825_));
 AOI21_X1 _6681_ (.A(_4130_),
    .B1(_1825_),
    .B2(_4131_),
    .ZN(_1826_));
 XOR2_X2 _6682_ (.A(_4115_),
    .B(_1826_),
    .Z(_1827_));
 INV_X1 _6683_ (.A(_1827_),
    .ZN(_4399_));
 INV_X1 _6684_ (.A(_4118_),
    .ZN(_1828_));
 INV_X1 _6685_ (.A(_4122_),
    .ZN(_1829_));
 INV_X1 _6686_ (.A(_4077_),
    .ZN(_1830_));
 AOI21_X4 _6687_ (.A(_3905_),
    .B1(_1615_),
    .B2(_3906_),
    .ZN(_1831_));
 INV_X1 _6688_ (.A(_4078_),
    .ZN(_1832_));
 OAI21_X4 _6689_ (.A(_1830_),
    .B1(_1831_),
    .B2(_1832_),
    .ZN(_1833_));
 AOI21_X4 _6690_ (.A(_4126_),
    .B1(_4127_),
    .B2(_1833_),
    .ZN(_1834_));
 INV_X1 _6691_ (.A(_4123_),
    .ZN(_1835_));
 OAI21_X4 _6692_ (.A(_1829_),
    .B1(_1834_),
    .B2(_1835_),
    .ZN(_1836_));
 AOI21_X2 _6693_ (.A(_4136_),
    .B1(_1836_),
    .B2(_4137_),
    .ZN(_1837_));
 INV_X1 _6694_ (.A(_4119_),
    .ZN(_1838_));
 OAI21_X4 _6695_ (.A(_1828_),
    .B1(_1837_),
    .B2(_1838_),
    .ZN(_1839_));
 XNOR2_X1 _6696_ (.A(_4131_),
    .B(_1839_),
    .ZN(_1840_));
 INV_X2 _6697_ (.A(_1840_),
    .ZN(_4383_));
 XOR2_X2 _6698_ (.A(_4133_),
    .B(_1823_),
    .Z(_4367_));
 XNOR2_X2 _6699_ (.A(_4137_),
    .B(_1836_),
    .ZN(_1841_));
 INV_X1 _6700_ (.A(_1841_),
    .ZN(_4351_));
 XNOR2_X2 _6701_ (.A(_4123_),
    .B(_1820_),
    .ZN(_1842_));
 INV_X1 _6702_ (.A(_1842_),
    .ZN(_4283_));
 XNOR2_X1 _6703_ (.A(_1833_),
    .B(_4127_),
    .ZN(_1843_));
 INV_X2 _6704_ (.A(_1843_),
    .ZN(_4242_));
 BUF_X16 _6705_ (.A(_1791_),
    .Z(_4198_));
 NAND3_X1 _6706_ (.A1(_1842_),
    .A2(_4174_),
    .A3(_1843_),
    .ZN(_1844_));
 NOR3_X1 _6707_ (.A1(_4367_),
    .A2(_4351_),
    .A3(_1844_),
    .ZN(_1845_));
 NAND3_X1 _6708_ (.A1(_1827_),
    .A2(_1840_),
    .A3(_1845_),
    .ZN(_1846_));
 NAND2_X1 _6709_ (.A1(net3),
    .A2(_1846_),
    .ZN(_1847_));
 INV_X1 _6710_ (.A(_3941_),
    .ZN(_1848_));
 AOI21_X1 _6711_ (.A(_3853_),
    .B1(_1561_),
    .B2(_1533_),
    .ZN(_1849_));
 OAI21_X1 _6712_ (.A(_1509_),
    .B1(_1849_),
    .B2(_1535_),
    .ZN(_1850_));
 AND2_X1 _6713_ (.A1(_3802_),
    .A2(_1850_),
    .ZN(_1851_));
 OAI21_X2 _6714_ (.A(_3942_),
    .B1(_3801_),
    .B2(_1851_),
    .ZN(_1852_));
 NAND2_X1 _6715_ (.A1(_1848_),
    .A2(_1852_),
    .ZN(_1853_));
 AOI21_X2 _6716_ (.A(_1853_),
    .B1(_1678_),
    .B2(_1672_),
    .ZN(_1854_));
 AND2_X2 _6717_ (.A1(_1848_),
    .A2(_1852_),
    .ZN(_1855_));
 NOR3_X2 _6718_ (.A1(_1697_),
    .A2(net126),
    .A3(_1855_),
    .ZN(_1856_));
 AOI21_X2 _6719_ (.A(_1320_),
    .B1(_1419_),
    .B2(_1488_),
    .ZN(_1857_));
 OAI21_X1 _6720_ (.A(_1857_),
    .B1(_1491_),
    .B2(_1490_),
    .ZN(_1858_));
 NAND3_X1 _6721_ (.A1(_1320_),
    .A2(_1475_),
    .A3(_1481_),
    .ZN(_1859_));
 AOI211_X4 _6722_ (.A(_1854_),
    .B(_1856_),
    .C1(_1858_),
    .C2(_1859_),
    .ZN(_1860_));
 OAI21_X2 _6723_ (.A(_1855_),
    .B1(net126),
    .B2(_1697_),
    .ZN(_1861_));
 NAND3_X2 _6724_ (.A1(_1672_),
    .A2(_1678_),
    .A3(_1853_),
    .ZN(_1862_));
 AOI221_X2 _6725_ (.A(_1492_),
    .B1(_1861_),
    .B2(_1862_),
    .C1(_1857_),
    .C2(_1498_),
    .ZN(_1863_));
 NOR3_X4 _6726_ (.A1(net4),
    .A2(_1860_),
    .A3(_1863_),
    .ZN(_1864_));
 INV_X1 _6727_ (.A(_3981_),
    .ZN(_1865_));
 NAND3_X2 _6728_ (.A1(_3926_),
    .A2(_3927_),
    .A3(_1865_),
    .ZN(_1866_));
 NOR3_X1 _6729_ (.A1(_4023_),
    .A2(_3977_),
    .A3(_4027_),
    .ZN(_1867_));
 INV_X1 _6730_ (.A(_1867_),
    .ZN(_1868_));
 OR2_X1 _6731_ (.A1(_4019_),
    .A2(_1868_),
    .ZN(_1869_));
 OR2_X2 _6732_ (.A1(_4015_),
    .A2(_1869_),
    .ZN(_1870_));
 NOR3_X4 _6733_ (.A1(_3974_),
    .A2(_1866_),
    .A3(_1870_),
    .ZN(_1871_));
 OAI221_X4 _6734_ (.A(_1858_),
    .B1(_1854_),
    .B2(_1856_),
    .C1(_1498_),
    .C2(net1),
    .ZN(_1872_));
 OAI211_X4 _6735_ (.A(_1861_),
    .B(_1862_),
    .C1(net145),
    .C2(_1492_),
    .ZN(_1873_));
 AOI211_X2 _6736_ (.A(_1591_),
    .B(_1871_),
    .C1(_1872_),
    .C2(_1873_),
    .ZN(_1874_));
 INV_X1 _6737_ (.A(_4114_),
    .ZN(_1875_));
 AND2_X4 _6738_ (.A1(_4131_),
    .A2(_1839_),
    .ZN(_1876_));
 OAI21_X4 _6739_ (.A(_4115_),
    .B1(_4130_),
    .B2(_1876_),
    .ZN(_1877_));
 AND2_X4 _6740_ (.A1(_1875_),
    .A2(_1877_),
    .ZN(_1878_));
 AOI21_X4 _6741_ (.A(_1878_),
    .B1(_1702_),
    .B2(_1694_),
    .ZN(_1879_));
 NAND2_X4 _6742_ (.A1(_1875_),
    .A2(_1877_),
    .ZN(_1880_));
 NOR3_X4 _6743_ (.A1(_1880_),
    .A2(_1705_),
    .A3(_1704_),
    .ZN(_1881_));
 OAI22_X4 _6744_ (.A1(_1864_),
    .A2(_1874_),
    .B1(_1879_),
    .B2(_1881_),
    .ZN(_1882_));
 NAND3_X4 _6745_ (.A1(net220),
    .A2(_1873_),
    .A3(_1872_),
    .ZN(_1883_));
 NOR2_X2 _6746_ (.A1(_1591_),
    .A2(_1871_),
    .ZN(_1884_));
 OAI21_X4 _6747_ (.A(_1884_),
    .B1(_1863_),
    .B2(_1860_),
    .ZN(_1885_));
 OAI21_X4 _6748_ (.A(_1880_),
    .B1(net134),
    .B2(_1704_),
    .ZN(_1886_));
 NAND3_X4 _6749_ (.A1(_1694_),
    .A2(_1702_),
    .A3(_1878_),
    .ZN(_1887_));
 NAND4_X4 _6750_ (.A1(_1883_),
    .A2(_1885_),
    .A3(_1886_),
    .A4(_1887_),
    .ZN(_1888_));
 NAND2_X4 _6751_ (.A1(_1882_),
    .A2(_1888_),
    .ZN(_1889_));
 MUX2_X1 _6752_ (.A(net69),
    .B(_1847_),
    .S(_1889_),
    .Z(_4138_));
 AOI22_X4 _6753_ (.A1(_1883_),
    .A2(_1885_),
    .B1(_1886_),
    .B2(_1887_),
    .ZN(_1890_));
 NOR4_X4 _6754_ (.A1(_1879_),
    .A2(_1874_),
    .A3(_1864_),
    .A4(_1881_),
    .ZN(_1891_));
 NOR3_X4 _6755_ (.A1(net3),
    .A2(_1890_),
    .A3(_1891_),
    .ZN(_1892_));
 NOR3_X2 _6756_ (.A1(_3933_),
    .A2(_4080_),
    .A3(_4242_),
    .ZN(_1893_));
 NAND3_X1 _6757_ (.A1(_1841_),
    .A2(_1842_),
    .A3(_1893_),
    .ZN(_1894_));
 OR3_X2 _6758_ (.A1(_4383_),
    .A2(net181),
    .A3(_1894_),
    .ZN(_1895_));
 OAI21_X2 _6759_ (.A(net3),
    .B1(_4399_),
    .B2(_1895_),
    .ZN(_1896_));
 AOI21_X4 _6760_ (.A(_1896_),
    .B1(net195),
    .B2(_1888_),
    .ZN(_1897_));
 NOR2_X1 _6761_ (.A1(_1892_),
    .A2(_1897_),
    .ZN(_4178_));
 MUX2_X1 _6762_ (.A(net69),
    .B(_1847_),
    .S(_1889_),
    .Z(_4182_));
 NOR2_X1 _6763_ (.A1(_1892_),
    .A2(_1897_),
    .ZN(_4187_));
 MUX2_X1 _6764_ (.A(net69),
    .B(_1847_),
    .S(_1889_),
    .Z(_4143_));
 NOR2_X1 _6765_ (.A1(_1892_),
    .A2(_1897_),
    .ZN(_4191_));
 XNOR2_X2 _6766_ (.A(_1889_),
    .B(_1847_),
    .ZN(_4147_));
 NAND2_X1 _6767_ (.A1(net277),
    .A2(_1895_),
    .ZN(_1898_));
 XNOR2_X1 _6768_ (.A(_1827_),
    .B(_1898_),
    .ZN(_4195_));
 NOR2_X1 _6769_ (.A1(_1845_),
    .A2(_4223_),
    .ZN(_1899_));
 XNOR2_X2 _6770_ (.A(_4383_),
    .B(_1899_),
    .ZN(_4151_));
 NAND2_X1 _6771_ (.A1(_1791_),
    .A2(_1894_),
    .ZN(_1900_));
 XOR2_X2 _6772_ (.A(net181),
    .B(_1900_),
    .Z(_4157_));
 NAND2_X1 _6773_ (.A1(net277),
    .A2(_1844_),
    .ZN(_1901_));
 XNOR2_X1 _6774_ (.A(_1841_),
    .B(_1901_),
    .ZN(_4160_));
 NOR2_X1 _6775_ (.A1(_4223_),
    .A2(_1893_),
    .ZN(_1902_));
 XNOR2_X1 _6776_ (.A(_4283_),
    .B(_1902_),
    .ZN(_4165_));
 NOR2_X4 _6777_ (.A1(_4174_),
    .A2(_4223_),
    .ZN(_1903_));
 XNOR2_X2 _6778_ (.A(_4242_),
    .B(_1903_),
    .ZN(_4169_));
 NOR2_X1 _6779_ (.A1(_4198_),
    .A2(_4173_),
    .ZN(_1904_));
 AOI21_X2 _6780_ (.A(_1904_),
    .B1(net277),
    .B2(_4175_),
    .ZN(_2989_));
 INV_X1 _6781_ (.A(_4141_),
    .ZN(_1905_));
 INV_X1 _6782_ (.A(_4188_),
    .ZN(_1906_));
 INV_X1 _6783_ (.A(_4192_),
    .ZN(_1907_));
 INV_X1 _6784_ (.A(_4196_),
    .ZN(_1908_));
 INV_X1 _6785_ (.A(_4158_),
    .ZN(_1909_));
 INV_X1 _6786_ (.A(_4166_),
    .ZN(_1910_));
 AOI21_X1 _6787_ (.A(_4170_),
    .B1(_4171_),
    .B2(_2990_),
    .ZN(_1911_));
 INV_X1 _6788_ (.A(_4167_),
    .ZN(_1912_));
 OAI21_X2 _6789_ (.A(_1910_),
    .B1(_1911_),
    .B2(_1912_),
    .ZN(_1913_));
 AOI21_X1 _6790_ (.A(_4162_),
    .B1(_1913_),
    .B2(_4163_),
    .ZN(_1914_));
 INV_X1 _6791_ (.A(_4159_),
    .ZN(_1915_));
 OAI21_X2 _6792_ (.A(_1909_),
    .B1(_1914_),
    .B2(_1915_),
    .ZN(_1916_));
 AOI21_X1 _6793_ (.A(_4152_),
    .B1(_1916_),
    .B2(_4155_),
    .ZN(_1917_));
 INV_X1 _6794_ (.A(_4197_),
    .ZN(_1918_));
 OAI21_X2 _6795_ (.A(_1908_),
    .B1(_1917_),
    .B2(_1918_),
    .ZN(_1919_));
 AOI21_X1 _6796_ (.A(_4148_),
    .B1(_1919_),
    .B2(_4149_),
    .ZN(_1920_));
 INV_X1 _6797_ (.A(_4193_),
    .ZN(_1921_));
 OAI21_X2 _6798_ (.A(_1907_),
    .B1(_1920_),
    .B2(_1921_),
    .ZN(_1922_));
 AOI21_X1 _6799_ (.A(_4144_),
    .B1(_1922_),
    .B2(_4145_),
    .ZN(_1923_));
 INV_X1 _6800_ (.A(_4189_),
    .ZN(_1924_));
 OAI21_X2 _6801_ (.A(_1906_),
    .B1(_1923_),
    .B2(_1924_),
    .ZN(_1925_));
 AOI21_X1 _6802_ (.A(_4184_),
    .B1(_1925_),
    .B2(_4185_),
    .ZN(_1926_));
 INV_X1 _6803_ (.A(_1926_),
    .ZN(_1927_));
 AOI21_X2 _6804_ (.A(_4180_),
    .B1(_1927_),
    .B2(_4181_),
    .ZN(_1928_));
 XNOR2_X2 _6805_ (.A(_1905_),
    .B(_1928_),
    .ZN(_1929_));
 INV_X1 _6806_ (.A(_1929_),
    .ZN(_4483_));
 INV_X1 _6807_ (.A(_2992_),
    .ZN(_2988_));
 INV_X1 _6808_ (.A(_4184_),
    .ZN(_1930_));
 INV_X1 _6809_ (.A(_4145_),
    .ZN(_1931_));
 INV_X1 _6810_ (.A(_4148_),
    .ZN(_1932_));
 AOI21_X2 _6811_ (.A(_4152_),
    .B1(_4153_),
    .B2(_4158_),
    .ZN(_1933_));
 NAND2_X2 _6812_ (.A1(_4159_),
    .A2(_4155_),
    .ZN(_1934_));
 INV_X1 _6813_ (.A(_4176_),
    .ZN(_1935_));
 INV_X1 _6814_ (.A(_4177_),
    .ZN(_1936_));
 OAI21_X4 _6815_ (.A(_1935_),
    .B1(_1936_),
    .B2(_2992_),
    .ZN(_1937_));
 AOI21_X4 _6816_ (.A(_4170_),
    .B1(_4171_),
    .B2(_1937_),
    .ZN(_1938_));
 OAI21_X4 _6817_ (.A(_1910_),
    .B1(_1938_),
    .B2(_1912_),
    .ZN(_1939_));
 AOI21_X4 _6818_ (.A(_4162_),
    .B1(_4163_),
    .B2(_1939_),
    .ZN(_1940_));
 OAI21_X4 _6819_ (.A(_1933_),
    .B1(_1940_),
    .B2(_1934_),
    .ZN(_1941_));
 AOI21_X4 _6820_ (.A(_4196_),
    .B1(_1941_),
    .B2(_4197_),
    .ZN(_1942_));
 INV_X2 _6821_ (.A(_4149_),
    .ZN(_1943_));
 OAI21_X4 _6822_ (.A(_1932_),
    .B1(_1942_),
    .B2(_1943_),
    .ZN(_1944_));
 AOI21_X2 _6823_ (.A(_4192_),
    .B1(_1944_),
    .B2(_4193_),
    .ZN(_1945_));
 NOR2_X2 _6824_ (.A1(_1931_),
    .A2(_1945_),
    .ZN(_1946_));
 OAI21_X2 _6825_ (.A(_4189_),
    .B1(_4144_),
    .B2(_1946_),
    .ZN(_1947_));
 INV_X2 _6826_ (.A(_1947_),
    .ZN(_1948_));
 OAI21_X2 _6827_ (.A(_4185_),
    .B1(_4188_),
    .B2(_1948_),
    .ZN(_1949_));
 NAND2_X2 _6828_ (.A1(_1949_),
    .A2(_1930_),
    .ZN(_1950_));
 XOR2_X2 _6829_ (.A(_4181_),
    .B(_1950_),
    .Z(_4475_));
 XNOR2_X2 _6830_ (.A(_4185_),
    .B(_1925_),
    .ZN(_1951_));
 INV_X1 _6831_ (.A(_1951_),
    .ZN(_4467_));
 NOR3_X1 _6832_ (.A1(_4189_),
    .A2(_4144_),
    .A3(_1946_),
    .ZN(_1952_));
 NOR2_X2 _6833_ (.A1(_1948_),
    .A2(_1952_),
    .ZN(_4459_));
 XNOR2_X2 _6834_ (.A(_4145_),
    .B(_1922_),
    .ZN(_1953_));
 INV_X1 _6835_ (.A(_1953_),
    .ZN(_4451_));
 XNOR2_X2 _6836_ (.A(_1943_),
    .B(_1919_),
    .ZN(_4438_));
 INV_X1 _6837_ (.A(_4200_),
    .ZN(_1954_));
 INV_X1 _6838_ (.A(_4204_),
    .ZN(_1955_));
 INV_X1 _6839_ (.A(_4206_),
    .ZN(_1956_));
 INV_X1 _6840_ (.A(_4210_),
    .ZN(_1957_));
 INV_X1 _6841_ (.A(_4212_),
    .ZN(_1958_));
 INV_X1 _6842_ (.A(_4216_),
    .ZN(_1959_));
 INV_X1 _6843_ (.A(_4218_),
    .ZN(_1960_));
 INV_X1 _6844_ (.A(_4222_),
    .ZN(_1961_));
 INV_X1 _6845_ (.A(_4225_),
    .ZN(_1962_));
 INV_X1 _6846_ (.A(_4231_),
    .ZN(_1963_));
 INV_X1 _6847_ (.A(_4237_),
    .ZN(_1964_));
 AOI21_X2 _6848_ (.A(_4240_),
    .B1(_4241_),
    .B2(_2940_),
    .ZN(_1965_));
 INV_X1 _6849_ (.A(_4238_),
    .ZN(_1966_));
 OAI21_X2 _6850_ (.A(_1964_),
    .B1(_1965_),
    .B2(_1966_),
    .ZN(_1967_));
 AOI21_X1 _6851_ (.A(_4234_),
    .B1(_1967_),
    .B2(_4235_),
    .ZN(_1968_));
 INV_X1 _6852_ (.A(_4232_),
    .ZN(_1969_));
 OAI21_X2 _6853_ (.A(_1963_),
    .B1(_1968_),
    .B2(_1969_),
    .ZN(_1970_));
 AND2_X2 _6854_ (.A1(_4229_),
    .A2(_1970_),
    .ZN(_1971_));
 OAI21_X2 _6855_ (.A(_4226_),
    .B1(_4228_),
    .B2(_1971_),
    .ZN(_1972_));
 AOI21_X4 _6856_ (.A(_1961_),
    .B1(_1972_),
    .B2(_1962_),
    .ZN(_1973_));
 OAI21_X4 _6857_ (.A(_4219_),
    .B1(_4221_),
    .B2(_1973_),
    .ZN(_1974_));
 AOI21_X4 _6858_ (.A(_1959_),
    .B1(_1974_),
    .B2(_1960_),
    .ZN(_1975_));
 OAI21_X4 _6859_ (.A(_4213_),
    .B1(_4215_),
    .B2(_1975_),
    .ZN(_1976_));
 AOI21_X4 _6860_ (.A(_1957_),
    .B1(_1976_),
    .B2(_1958_),
    .ZN(_1977_));
 OAI21_X4 _6861_ (.A(_4207_),
    .B1(_4209_),
    .B2(_1977_),
    .ZN(_1978_));
 AOI21_X4 _6862_ (.A(_1955_),
    .B1(_1978_),
    .B2(_1956_),
    .ZN(_1979_));
 OAI21_X4 _6863_ (.A(_4201_),
    .B1(_4203_),
    .B2(_1979_),
    .ZN(_1980_));
 NAND2_X4 _6864_ (.A1(_1980_),
    .A2(_1954_),
    .ZN(_1981_));
 INV_X2 _6865_ (.A(_1981_),
    .ZN(_1982_));
 BUF_X8 _6866_ (.A(_1982_),
    .Z(_1983_));
 BUF_X8 _6867_ (.A(_1983_),
    .Z(_4335_));
 INV_X1 _6868_ (.A(_4140_),
    .ZN(_1984_));
 AOI21_X4 _6869_ (.A(_4180_),
    .B1(_1950_),
    .B2(_4181_),
    .ZN(_1985_));
 OAI21_X4 _6870_ (.A(_1984_),
    .B1(_1905_),
    .B2(_1985_),
    .ZN(_1986_));
 NOR2_X1 _6871_ (.A1(_1710_),
    .A2(_1711_),
    .ZN(_1987_));
 NOR2_X1 _6872_ (.A1(_1591_),
    .A2(_1987_),
    .ZN(_1988_));
 OAI21_X2 _6873_ (.A(_1988_),
    .B1(_1705_),
    .B2(_1704_),
    .ZN(_1989_));
 OAI21_X4 _6874_ (.A(_1722_),
    .B1(_1760_),
    .B2(_1744_),
    .ZN(_1990_));
 AOI21_X4 _6875_ (.A(_3975_),
    .B1(_1990_),
    .B2(_3976_),
    .ZN(_1991_));
 INV_X4 _6876_ (.A(_1991_),
    .ZN(_1992_));
 AOI21_X2 _6877_ (.A(_1992_),
    .B1(_1872_),
    .B2(_1873_),
    .ZN(_1993_));
 NOR3_X2 _6878_ (.A1(_1860_),
    .A2(_1863_),
    .A3(_1991_),
    .ZN(_1994_));
 OAI221_X2 _6879_ (.A(_1989_),
    .B1(_1993_),
    .B2(_1994_),
    .C1(_1703_),
    .C2(net4),
    .ZN(_1995_));
 OAI21_X2 _6880_ (.A(_1991_),
    .B1(_1863_),
    .B2(_1860_),
    .ZN(_1996_));
 NAND3_X4 _6881_ (.A1(_1873_),
    .A2(_1872_),
    .A3(_1992_),
    .ZN(_1997_));
 OAI211_X4 _6882_ (.A(_1996_),
    .B(_1997_),
    .C1(_1706_),
    .C2(_1713_),
    .ZN(_1998_));
 AOI21_X4 _6883_ (.A(net147),
    .B1(_1995_),
    .B2(_1998_),
    .ZN(_1999_));
 NAND3_X1 _6884_ (.A1(net220),
    .A2(_1694_),
    .A3(_1702_),
    .ZN(_2000_));
 AOI211_X4 _6885_ (.A(_1993_),
    .B(_1994_),
    .C1(_2000_),
    .C2(_1989_),
    .ZN(_2001_));
 AOI221_X4 _6886_ (.A(_1706_),
    .B1(_1997_),
    .B2(_1996_),
    .C1(_1988_),
    .C2(_1703_),
    .ZN(_2002_));
 INV_X4 _6887_ (.A(_1986_),
    .ZN(_2003_));
 NOR3_X4 _6888_ (.A1(_2003_),
    .A2(_2002_),
    .A3(_2001_),
    .ZN(_2004_));
 OAI22_X4 _6889_ (.A1(_1892_),
    .A2(net196),
    .B1(_1999_),
    .B2(_2004_),
    .ZN(_2005_));
 NAND3_X4 _6890_ (.A1(_4223_),
    .A2(net148),
    .A3(net233),
    .ZN(_2006_));
 INV_X1 _6891_ (.A(_1896_),
    .ZN(_2007_));
 OAI21_X4 _6892_ (.A(_2007_),
    .B1(net183),
    .B2(_1890_),
    .ZN(_2008_));
 OAI21_X4 _6893_ (.A(_2003_),
    .B1(_2002_),
    .B2(_2001_),
    .ZN(_2009_));
 NAND3_X4 _6894_ (.A1(_1998_),
    .A2(_1995_),
    .A3(_1986_),
    .ZN(_2010_));
 NAND4_X4 _6895_ (.A1(_2009_),
    .A2(_2008_),
    .A3(_2006_),
    .A4(_2010_),
    .ZN(_2011_));
 NAND2_X4 _6896_ (.A1(_2005_),
    .A2(_2011_),
    .ZN(_2012_));
 BUF_X8 _6897_ (.A(_2012_),
    .Z(_2013_));
 INV_X2 _6898_ (.A(_2013_),
    .ZN(_4259_));
 INV_X1 _6899_ (.A(_4245_),
    .ZN(_2014_));
 INV_X1 _6900_ (.A(_4085_),
    .ZN(_2015_));
 INV_X1 _6901_ (.A(_4093_),
    .ZN(_2016_));
 INV_X1 _6902_ (.A(_4101_),
    .ZN(_2017_));
 AOI21_X2 _6903_ (.A(_4107_),
    .B1(_2984_),
    .B2(_4108_),
    .ZN(_2018_));
 INV_X1 _6904_ (.A(_4102_),
    .ZN(_2019_));
 OAI21_X4 _6905_ (.A(_2017_),
    .B1(_2019_),
    .B2(_2018_),
    .ZN(_2020_));
 AOI21_X4 _6906_ (.A(_4097_),
    .B1(_2020_),
    .B2(_4098_),
    .ZN(_2021_));
 INV_X1 _6907_ (.A(_4094_),
    .ZN(_2022_));
 OAI21_X4 _6908_ (.A(_2016_),
    .B1(_2021_),
    .B2(_2022_),
    .ZN(_2023_));
 AOI21_X4 _6909_ (.A(_4089_),
    .B1(_2023_),
    .B2(_4090_),
    .ZN(_2024_));
 INV_X1 _6910_ (.A(_4086_),
    .ZN(_2025_));
 OAI21_X4 _6911_ (.A(_2015_),
    .B1(_2024_),
    .B2(_2025_),
    .ZN(_2026_));
 NAND3_X2 _6912_ (.A1(_4250_),
    .A2(_4247_),
    .A3(_2026_),
    .ZN(_2027_));
 AOI21_X2 _6913_ (.A(_4081_),
    .B1(_4082_),
    .B2(_4249_),
    .ZN(_2028_));
 NAND2_X2 _6914_ (.A1(_2028_),
    .A2(_2027_),
    .ZN(_2029_));
 XNOR2_X2 _6915_ (.A(_2014_),
    .B(_2029_),
    .ZN(_4251_));
 INV_X2 _6916_ (.A(_4251_),
    .ZN(_4277_));
 INV_X1 _6917_ (.A(_4256_),
    .ZN(_2030_));
 INV_X1 _6918_ (.A(_4297_),
    .ZN(_2031_));
 INV_X1 _6919_ (.A(_4264_),
    .ZN(_2032_));
 INV_X1 _6920_ (.A(_4272_),
    .ZN(_2033_));
 AOI21_X2 _6921_ (.A(_4274_),
    .B1(_4275_),
    .B2(_3005_),
    .ZN(_2034_));
 INV_X2 _6922_ (.A(_4273_),
    .ZN(_2035_));
 OAI21_X4 _6923_ (.A(_2033_),
    .B1(_2034_),
    .B2(_2035_),
    .ZN(_2036_));
 AOI21_X1 _6924_ (.A(_4268_),
    .B1(_2036_),
    .B2(_4269_),
    .ZN(_2037_));
 INV_X1 _6925_ (.A(_4265_),
    .ZN(_2038_));
 OAI21_X2 _6926_ (.A(_2032_),
    .B1(_2037_),
    .B2(_2038_),
    .ZN(_2039_));
 AOI21_X2 _6927_ (.A(_4301_),
    .B1(_2039_),
    .B2(_4302_),
    .ZN(_2040_));
 INV_X1 _6928_ (.A(_4298_),
    .ZN(_2041_));
 OAI21_X4 _6929_ (.A(_2031_),
    .B1(_2041_),
    .B2(_2040_),
    .ZN(_2042_));
 AOI21_X4 _6930_ (.A(_4293_),
    .B1(net98),
    .B2(_2042_),
    .ZN(_2043_));
 INV_X1 _6931_ (.A(_4257_),
    .ZN(_2044_));
 OAI21_X4 _6932_ (.A(_2030_),
    .B1(_2043_),
    .B2(_2044_),
    .ZN(_2045_));
 XNOR2_X2 _6933_ (.A(net235),
    .B(_4254_),
    .ZN(_4304_));
 BUF_X16 _6934_ (.A(_1981_),
    .Z(_2046_));
 BUF_X16 _6935_ (.A(_2046_),
    .Z(_4307_));
 NOR2_X1 _6936_ (.A1(_4307_),
    .A2(_4277_),
    .ZN(_2047_));
 AOI21_X2 _6937_ (.A(_2047_),
    .B1(_4307_),
    .B2(_4280_),
    .ZN(_2998_));
 INV_X1 _6938_ (.A(_2998_),
    .ZN(_2995_));
 INV_X1 _6939_ (.A(_4244_),
    .ZN(_2048_));
 AOI21_X1 _6940_ (.A(_4081_),
    .B1(_1815_),
    .B2(_4247_),
    .ZN(_2049_));
 OAI21_X2 _6941_ (.A(_2048_),
    .B1(_2049_),
    .B2(_2014_),
    .ZN(_2050_));
 XOR2_X2 _6942_ (.A(_4286_),
    .B(_2050_),
    .Z(_4287_));
 BUF_X2 _6943_ (.A(_4290_),
    .Z(_2051_));
 XNOR2_X2 _6944_ (.A(_4193_),
    .B(_1944_),
    .ZN(_2052_));
 INV_X1 _6945_ (.A(_2052_),
    .ZN(_2053_));
 NOR2_X1 _6946_ (.A1(_4438_),
    .A2(_2053_),
    .ZN(_2054_));
 NAND2_X1 _6947_ (.A1(_1953_),
    .A2(_2054_),
    .ZN(_2055_));
 NOR2_X1 _6948_ (.A1(_4459_),
    .A2(_2055_),
    .ZN(_2056_));
 NAND2_X1 _6949_ (.A1(_1951_),
    .A2(_2056_),
    .ZN(_2057_));
 NOR2_X2 _6950_ (.A1(_4475_),
    .A2(_2057_),
    .ZN(_2058_));
 AOI21_X2 _6951_ (.A(_1982_),
    .B1(_2058_),
    .B2(_1929_),
    .ZN(_2059_));
 INV_X1 _6952_ (.A(_4293_),
    .ZN(_2060_));
 INV_X1 _6953_ (.A(_4301_),
    .ZN(_2061_));
 INV_X1 _6954_ (.A(_4268_),
    .ZN(_2062_));
 AOI21_X4 _6955_ (.A(_4272_),
    .B1(net274),
    .B2(_3007_),
    .ZN(_2063_));
 INV_X1 _6956_ (.A(_4269_),
    .ZN(_2064_));
 OAI21_X4 _6957_ (.A(_2062_),
    .B1(_2063_),
    .B2(_2064_),
    .ZN(_2065_));
 AOI21_X2 _6958_ (.A(_4264_),
    .B1(_2065_),
    .B2(_4265_),
    .ZN(_2066_));
 INV_X1 _6959_ (.A(_4302_),
    .ZN(_2067_));
 OAI21_X4 _6960_ (.A(_2061_),
    .B1(_2066_),
    .B2(_2067_),
    .ZN(_2068_));
 AOI21_X4 _6961_ (.A(_4297_),
    .B1(_2068_),
    .B2(_4298_),
    .ZN(_2069_));
 INV_X2 _6962_ (.A(_4294_),
    .ZN(_2070_));
 OAI21_X4 _6963_ (.A(_2060_),
    .B1(_2069_),
    .B2(_2070_),
    .ZN(_2071_));
 AND2_X4 _6964_ (.A1(_4257_),
    .A2(_2071_),
    .ZN(_2072_));
 NAND2_X4 _6965_ (.A1(_4251_),
    .A2(_2072_),
    .ZN(_2073_));
 NOR2_X4 _6966_ (.A1(_2073_),
    .A2(_2059_),
    .ZN(_2074_));
 NAND2_X2 _6967_ (.A1(_1929_),
    .A2(_2058_),
    .ZN(_4258_));
 NAND2_X4 _6968_ (.A1(_1981_),
    .A2(_4258_),
    .ZN(_2075_));
 NAND2_X4 _6969_ (.A1(_4277_),
    .A2(_2072_),
    .ZN(_2076_));
 NOR2_X4 _6970_ (.A1(_2075_),
    .A2(_2076_),
    .ZN(_2077_));
 OAI211_X4 _6971_ (.A(net186),
    .B(net178),
    .C1(_2074_),
    .C2(_2077_),
    .ZN(_2078_));
 AOI22_X4 _6972_ (.A1(_2006_),
    .A2(_2008_),
    .B1(_2009_),
    .B2(_2010_),
    .ZN(_2079_));
 NOR4_X4 _6973_ (.A1(_1892_),
    .A2(net197),
    .A3(_1999_),
    .A4(net124),
    .ZN(_2080_));
 NOR2_X4 _6974_ (.A1(_2046_),
    .A2(_2076_),
    .ZN(_2081_));
 NOR2_X4 _6975_ (.A1(_1983_),
    .A2(_2073_),
    .ZN(_2082_));
 OAI22_X4 _6976_ (.A1(_2079_),
    .A2(_2080_),
    .B1(_2081_),
    .B2(_2082_),
    .ZN(_2083_));
 AOI21_X1 _6977_ (.A(_4253_),
    .B1(_4256_),
    .B2(_4254_),
    .ZN(_2084_));
 NAND3_X4 _6978_ (.A1(_2078_),
    .A2(net247),
    .A3(_2084_),
    .ZN(_2085_));
 XNOR2_X2 _6979_ (.A(_2051_),
    .B(_2085_),
    .ZN(_4303_));
 INV_X4 _6980_ (.A(net265),
    .ZN(_4546_));
 INV_X1 _6981_ (.A(_4312_),
    .ZN(_2086_));
 INV_X1 _6982_ (.A(_4318_),
    .ZN(_2087_));
 INV_X1 _6983_ (.A(_4319_),
    .ZN(_2088_));
 INV_X1 _6984_ (.A(_4324_),
    .ZN(_2089_));
 INV_X1 _6985_ (.A(_4330_),
    .ZN(_2090_));
 INV_X1 _6986_ (.A(_4331_),
    .ZN(_2091_));
 INV_X1 _6987_ (.A(_4337_),
    .ZN(_2092_));
 INV_X1 _6988_ (.A(_4235_),
    .ZN(_2093_));
 XNOR2_X1 _6989_ (.A(_2093_),
    .B(_1967_),
    .ZN(_2094_));
 AOI21_X1 _6990_ (.A(_4340_),
    .B1(_2094_),
    .B2(_4341_),
    .ZN(_2095_));
 INV_X1 _6991_ (.A(_4338_),
    .ZN(_2096_));
 OAI21_X1 _6992_ (.A(_2092_),
    .B1(_2095_),
    .B2(_2096_),
    .ZN(_2097_));
 AOI21_X1 _6993_ (.A(_4333_),
    .B1(_2097_),
    .B2(_4334_),
    .ZN(_2098_));
 OAI21_X1 _6994_ (.A(_2090_),
    .B1(_2091_),
    .B2(_2098_),
    .ZN(_2099_));
 AOI21_X1 _6995_ (.A(_4327_),
    .B1(_2099_),
    .B2(_4328_),
    .ZN(_2100_));
 INV_X1 _6996_ (.A(_4325_),
    .ZN(_2101_));
 OAI21_X1 _6997_ (.A(_2089_),
    .B1(_2100_),
    .B2(_2101_),
    .ZN(_2102_));
 AOI21_X1 _6998_ (.A(_4321_),
    .B1(_2102_),
    .B2(_4322_),
    .ZN(_2103_));
 OAI21_X1 _6999_ (.A(_2087_),
    .B1(_2088_),
    .B2(_2103_),
    .ZN(_2104_));
 AOI21_X1 _7000_ (.A(_4315_),
    .B1(_2104_),
    .B2(_4316_),
    .ZN(_2105_));
 INV_X1 _7001_ (.A(_4313_),
    .ZN(_2106_));
 OAI21_X2 _7002_ (.A(_2086_),
    .B1(_2105_),
    .B2(_2106_),
    .ZN(_2107_));
 AOI21_X4 _7003_ (.A(_4309_),
    .B1(_2107_),
    .B2(_4310_),
    .ZN(_2108_));
 MUX2_X1 _7004_ (.A(_4306_),
    .B(_4546_),
    .S(_2108_),
    .Z(_3000_));
 INV_X1 _7005_ (.A(_4354_),
    .ZN(_2109_));
 AOI21_X4 _7006_ (.A(_4244_),
    .B1(_2029_),
    .B2(_4245_),
    .ZN(_2110_));
 INV_X4 _7007_ (.A(_2110_),
    .ZN(_2111_));
 AOI21_X4 _7008_ (.A(_4285_),
    .B1(_2111_),
    .B2(_4286_),
    .ZN(_2112_));
 XNOR2_X1 _7009_ (.A(_2109_),
    .B(_2112_),
    .ZN(_2113_));
 INV_X1 _7010_ (.A(_2113_),
    .ZN(_4355_));
 BUF_X2 _7011_ (.A(_4358_),
    .Z(_2114_));
 INV_X1 _7012_ (.A(_4253_),
    .ZN(_2115_));
 NAND2_X2 _7013_ (.A1(_4251_),
    .A2(_2045_),
    .ZN(_2116_));
 NOR2_X2 _7014_ (.A1(_2059_),
    .A2(_2116_),
    .ZN(_2117_));
 NAND2_X2 _7015_ (.A1(_4277_),
    .A2(_2045_),
    .ZN(_2118_));
 NOR2_X2 _7016_ (.A1(_2075_),
    .A2(_2118_),
    .ZN(_2119_));
 OAI211_X2 _7017_ (.A(net186),
    .B(net178),
    .C1(_2117_),
    .C2(_2119_),
    .ZN(_2120_));
 NOR2_X1 _7018_ (.A1(_2046_),
    .A2(_2118_),
    .ZN(_2121_));
 NOR2_X2 _7019_ (.A1(_1983_),
    .A2(_2116_),
    .ZN(_2122_));
 OAI22_X1 _7020_ (.A1(_2079_),
    .A2(_2080_),
    .B1(_2121_),
    .B2(_2122_),
    .ZN(_2123_));
 NAND3_X1 _7021_ (.A1(_2123_),
    .A2(_2120_),
    .A3(_2115_),
    .ZN(_2124_));
 AOI21_X2 _7022_ (.A(_4289_),
    .B1(_2124_),
    .B2(_2051_),
    .ZN(_2125_));
 XNOR2_X2 _7023_ (.A(_2125_),
    .B(_2114_),
    .ZN(_4550_));
 INV_X1 _7024_ (.A(_4353_),
    .ZN(_2126_));
 AOI21_X1 _7025_ (.A(_4285_),
    .B1(_2050_),
    .B2(_4286_),
    .ZN(_2127_));
 OAI21_X2 _7026_ (.A(_2126_),
    .B1(_2127_),
    .B2(_2109_),
    .ZN(_2128_));
 XNOR2_X2 _7027_ (.A(_4370_),
    .B(_2128_),
    .ZN(_2129_));
 INV_X1 _7028_ (.A(_2129_),
    .ZN(_4372_));
 BUF_X2 _7029_ (.A(_4374_),
    .Z(_2130_));
 OR3_X1 _7030_ (.A1(_2051_),
    .A2(_4289_),
    .A3(_4357_),
    .ZN(_2131_));
 NOR2_X1 _7031_ (.A1(_4289_),
    .A2(_4357_),
    .ZN(_2132_));
 NAND2_X1 _7032_ (.A1(_2084_),
    .A2(_2132_),
    .ZN(_2133_));
 NAND2_X2 _7033_ (.A1(_2078_),
    .A2(_2083_),
    .ZN(_2134_));
 OAI221_X2 _7034_ (.A(_2131_),
    .B1(_2134_),
    .B2(_2133_),
    .C1(_2114_),
    .C2(_4357_),
    .ZN(_2135_));
 XNOR2_X2 _7035_ (.A(net188),
    .B(_2130_),
    .ZN(_4554_));
 OAI21_X4 _7036_ (.A(_2126_),
    .B1(_2109_),
    .B2(_2112_),
    .ZN(_2136_));
 AOI21_X4 _7037_ (.A(_4369_),
    .B1(_4370_),
    .B2(_2136_),
    .ZN(_2137_));
 XNOR2_X2 _7038_ (.A(_4386_),
    .B(net132),
    .ZN(_4387_));
 BUF_X2 _7039_ (.A(_4390_),
    .Z(_2138_));
 BUF_X2 _7040_ (.A(_4373_),
    .Z(_2139_));
 NAND4_X2 _7041_ (.A1(_2051_),
    .A2(_2114_),
    .A3(_4251_),
    .A4(_2045_),
    .ZN(_2140_));
 NOR2_X2 _7042_ (.A1(_2059_),
    .A2(_2140_),
    .ZN(_2141_));
 NAND4_X2 _7043_ (.A1(_2051_),
    .A2(_2114_),
    .A3(_4277_),
    .A4(_2045_),
    .ZN(_2142_));
 NOR2_X2 _7044_ (.A1(_2075_),
    .A2(_2142_),
    .ZN(_2143_));
 OAI211_X2 _7045_ (.A(net187),
    .B(net178),
    .C1(_2141_),
    .C2(_2143_),
    .ZN(_2144_));
 NOR2_X2 _7046_ (.A1(_2046_),
    .A2(_2142_),
    .ZN(_2145_));
 NOR2_X2 _7047_ (.A1(_1983_),
    .A2(_2140_),
    .ZN(_2146_));
 OAI22_X2 _7048_ (.A1(_2079_),
    .A2(_2080_),
    .B1(_2145_),
    .B2(_2146_),
    .ZN(_2147_));
 AOI21_X1 _7049_ (.A(_4289_),
    .B1(_4253_),
    .B2(_2051_),
    .ZN(_2148_));
 INV_X1 _7050_ (.A(_2148_),
    .ZN(_2149_));
 AOI21_X1 _7051_ (.A(_4357_),
    .B1(_2149_),
    .B2(_2114_),
    .ZN(_2150_));
 NAND3_X1 _7052_ (.A1(_2144_),
    .A2(_2147_),
    .A3(_2150_),
    .ZN(_2151_));
 AOI21_X2 _7053_ (.A(_2139_),
    .B1(_2151_),
    .B2(_2130_),
    .ZN(_2152_));
 XOR2_X2 _7054_ (.A(_2138_),
    .B(_2152_),
    .Z(_2153_));
 INV_X2 _7055_ (.A(_2153_),
    .ZN(_4558_));
 INV_X1 _7056_ (.A(_4385_),
    .ZN(_2154_));
 AOI21_X1 _7057_ (.A(_4369_),
    .B1(_2128_),
    .B2(_4370_),
    .ZN(_2155_));
 INV_X1 _7058_ (.A(_4386_),
    .ZN(_2156_));
 OAI21_X1 _7059_ (.A(_2154_),
    .B1(_2155_),
    .B2(_2156_),
    .ZN(_2157_));
 XOR2_X2 _7060_ (.A(_4402_),
    .B(_2157_),
    .Z(_4403_));
 CLKBUF_X2 _7061_ (.A(_4406_),
    .Z(_2158_));
 INV_X2 _7062_ (.A(_2158_),
    .ZN(_2159_));
 AND3_X1 _7063_ (.A1(_2130_),
    .A2(_2138_),
    .A3(_2159_),
    .ZN(_2160_));
 BUF_X2 _7064_ (.A(_4389_),
    .Z(_2161_));
 NOR3_X1 _7065_ (.A1(_2159_),
    .A2(_2139_),
    .A3(_2161_),
    .ZN(_2162_));
 MUX2_X1 _7066_ (.A(_2160_),
    .B(_2162_),
    .S(_2135_),
    .Z(_2163_));
 NOR4_X4 _7067_ (.A1(_2130_),
    .A2(_2159_),
    .A3(_2139_),
    .A4(_2161_),
    .ZN(_2164_));
 NOR3_X2 _7068_ (.A1(_2138_),
    .A2(_2159_),
    .A3(_2161_),
    .ZN(_2165_));
 NAND3_X1 _7069_ (.A1(_2138_),
    .A2(_2159_),
    .A3(_2139_),
    .ZN(_2166_));
 INV_X1 _7070_ (.A(_2161_),
    .ZN(_2167_));
 OAI21_X2 _7071_ (.A(_2166_),
    .B1(_2167_),
    .B2(_2158_),
    .ZN(_2168_));
 NOR4_X4 _7072_ (.A1(_2168_),
    .A2(_2164_),
    .A3(_2165_),
    .A4(_2163_),
    .ZN(_2169_));
 INV_X2 _7073_ (.A(net111),
    .ZN(_4561_));
 INV_X1 _7074_ (.A(_4190_),
    .ZN(_2170_));
 NAND3_X1 _7075_ (.A1(_2170_),
    .A2(_4103_),
    .A3(_4104_),
    .ZN(_2171_));
 OR2_X1 _7076_ (.A1(_4142_),
    .A2(_2171_),
    .ZN(_2172_));
 OR2_X1 _7077_ (.A1(_4183_),
    .A2(_4186_),
    .ZN(_2173_));
 OR3_X1 _7078_ (.A1(_4179_),
    .A2(_2172_),
    .A3(_2173_),
    .ZN(_2174_));
 OAI21_X1 _7079_ (.A(_1790_),
    .B1(_2174_),
    .B2(_4139_),
    .ZN(_2175_));
 OR3_X4 _7080_ (.A1(_2001_),
    .A2(_2002_),
    .A3(_2175_),
    .ZN(_2176_));
 OAI21_X4 _7081_ (.A(_4223_),
    .B1(_2001_),
    .B2(_2002_),
    .ZN(_2177_));
 OAI21_X4 _7082_ (.A(_2154_),
    .B1(_2137_),
    .B2(_2156_),
    .ZN(_2178_));
 AOI21_X4 _7083_ (.A(_4401_),
    .B1(_2178_),
    .B2(_4402_),
    .ZN(_2179_));
 INV_X4 _7084_ (.A(_2179_),
    .ZN(_2180_));
 OAI21_X4 _7085_ (.A(_2180_),
    .B1(net183),
    .B2(_1890_),
    .ZN(_2181_));
 NAND3_X4 _7086_ (.A1(net148),
    .A2(net233),
    .A3(_2179_),
    .ZN(_2182_));
 AOI22_X4 _7087_ (.A1(_2176_),
    .A2(_2177_),
    .B1(_2181_),
    .B2(_2182_),
    .ZN(_2183_));
 AND4_X4 _7088_ (.A1(_2181_),
    .A2(_2177_),
    .A3(_2182_),
    .A4(_2176_),
    .ZN(_2184_));
 OR2_X4 _7089_ (.A1(_2184_),
    .A2(_2183_),
    .ZN(_2185_));
 BUF_X8 _7090_ (.A(_2185_),
    .Z(_4424_));
 NOR2_X2 _7091_ (.A1(_4307_),
    .A2(_4424_),
    .ZN(_2186_));
 INV_X1 _7092_ (.A(_4403_),
    .ZN(_2187_));
 INV_X1 _7093_ (.A(_4279_),
    .ZN(_2188_));
 NOR3_X1 _7094_ (.A1(_2188_),
    .A2(_4287_),
    .A3(_4355_),
    .ZN(_2189_));
 NAND2_X1 _7095_ (.A1(_2129_),
    .A2(_2189_),
    .ZN(_2190_));
 OAI21_X2 _7096_ (.A(_2046_),
    .B1(_4387_),
    .B2(_2190_),
    .ZN(_2191_));
 AOI21_X2 _7097_ (.A(_4335_),
    .B1(_2187_),
    .B2(_2191_),
    .ZN(_2192_));
 AOI21_X1 _7098_ (.A(_2186_),
    .B1(_2192_),
    .B2(_4424_),
    .ZN(_4439_));
 MUX2_X1 _7099_ (.A(_4260_),
    .B(_2012_),
    .S(_1983_),
    .Z(_2193_));
 XOR2_X2 _7100_ (.A(net68),
    .B(_2193_),
    .Z(_2194_));
 OR2_X1 _7101_ (.A1(_2130_),
    .A2(_2139_),
    .ZN(_2195_));
 AOI21_X1 _7102_ (.A(_2161_),
    .B1(_2195_),
    .B2(_2138_),
    .ZN(_2196_));
 INV_X1 _7103_ (.A(_2150_),
    .ZN(_2197_));
 NOR3_X1 _7104_ (.A1(_2139_),
    .A2(_2161_),
    .A3(_2197_),
    .ZN(_2198_));
 AND2_X2 _7105_ (.A1(_2144_),
    .A2(_2147_),
    .ZN(_2199_));
 AOI21_X4 _7106_ (.A(_2196_),
    .B1(_2198_),
    .B2(_2199_),
    .ZN(_2200_));
 AOI21_X1 _7107_ (.A(_4405_),
    .B1(_2200_),
    .B2(_2158_),
    .ZN(_2201_));
 XNOR2_X2 _7108_ (.A(_2194_),
    .B(_2201_),
    .ZN(_4416_));
 NOR3_X2 _7109_ (.A1(_4110_),
    .A2(_4251_),
    .A3(_4287_),
    .ZN(_2202_));
 NAND3_X1 _7110_ (.A1(_2113_),
    .A2(_2129_),
    .A3(_2202_),
    .ZN(_2203_));
 NOR3_X4 _7111_ (.A1(_4403_),
    .A2(_4387_),
    .A3(_2203_),
    .ZN(_2204_));
 INV_X1 _7112_ (.A(_2204_),
    .ZN(_4423_));
 NAND2_X1 _7113_ (.A1(_2046_),
    .A2(_4423_),
    .ZN(_2205_));
 MUX2_X2 _7114_ (.A(_2046_),
    .B(_2205_),
    .S(_2185_),
    .Z(_4458_));
 INV_X1 _7115_ (.A(_4429_),
    .ZN(_2206_));
 INV_X1 _7116_ (.A(_4397_),
    .ZN(_2207_));
 INV_X1 _7117_ (.A(_4365_),
    .ZN(_2208_));
 INV_X1 _7118_ (.A(_4281_),
    .ZN(_2209_));
 INV_X1 _7119_ (.A(_4282_),
    .ZN(_2210_));
 OAI21_X1 _7120_ (.A(_2209_),
    .B1(_2210_),
    .B2(_2994_),
    .ZN(_2211_));
 AOI21_X2 _7121_ (.A(_4349_),
    .B1(_2211_),
    .B2(net96),
    .ZN(_2212_));
 INV_X1 _7122_ (.A(_4366_),
    .ZN(_2213_));
 OAI21_X1 _7123_ (.A(_2208_),
    .B1(_2212_),
    .B2(_2213_),
    .ZN(_2214_));
 AOI21_X2 _7124_ (.A(_4381_),
    .B1(_2214_),
    .B2(_4382_),
    .ZN(_2215_));
 INV_X1 _7125_ (.A(_4398_),
    .ZN(_2216_));
 OAI21_X4 _7126_ (.A(_2207_),
    .B1(_2215_),
    .B2(_2216_),
    .ZN(_2217_));
 AOI21_X4 _7127_ (.A(_4413_),
    .B1(_4414_),
    .B2(_2217_),
    .ZN(_2218_));
 INV_X2 _7128_ (.A(net93),
    .ZN(_2219_));
 OAI21_X4 _7129_ (.A(_2206_),
    .B1(_2218_),
    .B2(_2219_),
    .ZN(_2220_));
 AOI21_X4 _7130_ (.A(_4440_),
    .B1(_4441_),
    .B2(_2220_),
    .ZN(_2221_));
 NAND2_X1 _7131_ (.A1(_2052_),
    .A2(net160),
    .ZN(_2222_));
 INV_X1 _7132_ (.A(_2222_),
    .ZN(_2223_));
 NOR2_X4 _7133_ (.A1(_2221_),
    .A2(_2052_),
    .ZN(_2224_));
 NOR2_X2 _7134_ (.A1(_2223_),
    .A2(net285),
    .ZN(_2225_));
 XOR2_X2 _7135_ (.A(_4458_),
    .B(_2225_),
    .Z(_4447_));
 INV_X2 _7136_ (.A(_4447_),
    .ZN(_4491_));
 INV_X1 _7137_ (.A(_2108_),
    .ZN(_2226_));
 BUF_X4 _7138_ (.A(_2226_),
    .Z(_2227_));
 NOR2_X4 _7139_ (.A1(_2227_),
    .A2(net118),
    .ZN(_2228_));
 INV_X4 _7140_ (.A(_4304_),
    .ZN(_4542_));
 NOR3_X4 _7141_ (.A1(net193),
    .A2(_4546_),
    .A3(_4542_),
    .ZN(_2229_));
 NOR2_X4 _7142_ (.A1(net190),
    .A2(_4558_),
    .ZN(_2230_));
 NAND3_X1 _7143_ (.A1(net111),
    .A2(net291),
    .A3(_2230_),
    .ZN(_2231_));
 AND2_X1 _7144_ (.A1(_2227_),
    .A2(net113),
    .ZN(_2232_));
 AOI21_X1 _7145_ (.A(_2228_),
    .B1(_2231_),
    .B2(_2232_),
    .ZN(_4446_));
 AOI21_X1 _7146_ (.A(_2186_),
    .B1(_2192_),
    .B2(net68),
    .ZN(_4450_));
 INV_X1 _7147_ (.A(_4453_),
    .ZN(_2233_));
 INV_X1 _7148_ (.A(_4441_),
    .ZN(_2234_));
 INV_X1 _7149_ (.A(_4413_),
    .ZN(_2235_));
 INV_X1 _7150_ (.A(_4381_),
    .ZN(_2236_));
 INV_X1 _7151_ (.A(_4349_),
    .ZN(_2237_));
 INV_X2 _7152_ (.A(_4350_),
    .ZN(_2238_));
 OAI21_X4 _7153_ (.A(_2237_),
    .B1(_2238_),
    .B2(_2996_),
    .ZN(_2239_));
 AOI21_X4 _7154_ (.A(_4365_),
    .B1(_4366_),
    .B2(_2239_),
    .ZN(_2240_));
 INV_X1 _7155_ (.A(_4382_),
    .ZN(_2241_));
 OAI21_X4 _7156_ (.A(_2236_),
    .B1(_2241_),
    .B2(_2240_),
    .ZN(_2242_));
 AOI21_X4 _7157_ (.A(_4397_),
    .B1(_2242_),
    .B2(_4398_),
    .ZN(_2243_));
 INV_X1 _7158_ (.A(_4414_),
    .ZN(_2244_));
 OAI21_X4 _7159_ (.A(_2235_),
    .B1(_2244_),
    .B2(_2243_),
    .ZN(_2245_));
 AOI21_X4 _7160_ (.A(_4429_),
    .B1(_2245_),
    .B2(net209),
    .ZN(_2246_));
 NOR2_X4 _7161_ (.A1(_2234_),
    .A2(_2246_),
    .ZN(_2247_));
 NOR2_X4 _7162_ (.A1(_2247_),
    .A2(_4440_),
    .ZN(_2248_));
 NAND2_X1 _7163_ (.A1(_2052_),
    .A2(net135),
    .ZN(_2249_));
 NOR2_X1 _7164_ (.A1(_2052_),
    .A2(_2248_),
    .ZN(_2250_));
 OAI21_X1 _7165_ (.A(_2249_),
    .B1(_2250_),
    .B2(_4458_),
    .ZN(_2251_));
 XNOR2_X2 _7166_ (.A(_2233_),
    .B(_2251_),
    .ZN(_4490_));
 INV_X1 _7167_ (.A(_4490_),
    .ZN(_4454_));
 NOR2_X4 _7168_ (.A1(net193),
    .A2(_4554_),
    .ZN(_2252_));
 NAND4_X4 _7169_ (.A1(net119),
    .A2(_2153_),
    .A3(_2169_),
    .A4(_2252_),
    .ZN(_4415_));
 AOI21_X1 _7170_ (.A(_2228_),
    .B1(_2232_),
    .B2(net245),
    .ZN(_4455_));
 NOR4_X4 _7171_ (.A1(_2224_),
    .A2(net222),
    .A3(net146),
    .A4(_2046_),
    .ZN(_2253_));
 NOR3_X4 _7172_ (.A1(_1983_),
    .A2(net216),
    .A3(_2224_),
    .ZN(_2254_));
 AOI21_X4 _7173_ (.A(_2253_),
    .B1(_2254_),
    .B2(net68),
    .ZN(_2255_));
 NOR2_X2 _7174_ (.A1(_2233_),
    .A2(_2223_),
    .ZN(_2256_));
 AOI21_X4 _7175_ (.A(_4452_),
    .B1(_2255_),
    .B2(_2256_),
    .ZN(_2257_));
 XOR2_X2 _7176_ (.A(_4461_),
    .B(_2257_),
    .Z(_2258_));
 INV_X2 _7177_ (.A(net217),
    .ZN(_4463_));
 AOI21_X1 _7178_ (.A(_2228_),
    .B1(_2231_),
    .B2(_2232_),
    .ZN(_4462_));
 AOI21_X1 _7179_ (.A(_2186_),
    .B1(_2192_),
    .B2(_4424_),
    .ZN(_4466_));
 AOI21_X1 _7180_ (.A(_4460_),
    .B1(_4452_),
    .B2(_4461_),
    .ZN(_2259_));
 NOR3_X1 _7181_ (.A1(_1983_),
    .A2(_2053_),
    .A3(net215),
    .ZN(_2260_));
 OAI21_X1 _7182_ (.A(_2260_),
    .B1(net146),
    .B2(net222),
    .ZN(_2261_));
 AND2_X1 _7183_ (.A1(_4453_),
    .A2(_4461_),
    .ZN(_2262_));
 NAND2_X1 _7184_ (.A1(_1983_),
    .A2(_2052_),
    .ZN(_2263_));
 OAI211_X2 _7185_ (.A(_2261_),
    .B(_2262_),
    .C1(_2263_),
    .C2(net68),
    .ZN(_2264_));
 INV_X2 _7186_ (.A(_2248_),
    .ZN(_2265_));
 NOR3_X2 _7187_ (.A1(_2265_),
    .A2(net214),
    .A3(_1983_),
    .ZN(_2266_));
 OAI21_X1 _7188_ (.A(_2266_),
    .B1(net146),
    .B2(net222),
    .ZN(_2267_));
 NAND2_X1 _7189_ (.A1(_1983_),
    .A2(_2248_),
    .ZN(_2268_));
 OAI221_X1 _7190_ (.A(_2267_),
    .B1(_2268_),
    .B2(_2185_),
    .C1(_2265_),
    .C2(_2053_),
    .ZN(_2269_));
 OAI21_X2 _7191_ (.A(_2259_),
    .B1(_2269_),
    .B2(_2264_),
    .ZN(_2270_));
 XNOR2_X2 _7192_ (.A(_4469_),
    .B(_2270_),
    .ZN(_2271_));
 INV_X2 _7193_ (.A(_2271_),
    .ZN(_4471_));
 AOI21_X1 _7194_ (.A(_2228_),
    .B1(_2232_),
    .B2(net245),
    .ZN(_4470_));
 MUX2_X1 _7195_ (.A(_4307_),
    .B(_2205_),
    .S(_4424_),
    .Z(_4474_));
 BUF_X2 _7196_ (.A(_4477_),
    .Z(_2272_));
 BUF_X2 _7197_ (.A(_4468_),
    .Z(_2273_));
 OR3_X1 _7198_ (.A1(_4452_),
    .A2(_4460_),
    .A3(_2273_),
    .ZN(_2274_));
 AOI21_X2 _7199_ (.A(_2274_),
    .B1(_2256_),
    .B2(_2255_),
    .ZN(_2275_));
 OR2_X1 _7200_ (.A1(_4461_),
    .A2(_4460_),
    .ZN(_2276_));
 AOI21_X2 _7201_ (.A(_2273_),
    .B1(_2276_),
    .B2(_4469_),
    .ZN(_2277_));
 OR2_X1 _7202_ (.A1(_2275_),
    .A2(_2277_),
    .ZN(_2278_));
 XOR2_X2 _7203_ (.A(_2272_),
    .B(_2278_),
    .Z(_2279_));
 INV_X2 _7204_ (.A(_2279_),
    .ZN(_4479_));
 AOI21_X1 _7205_ (.A(_2228_),
    .B1(_2231_),
    .B2(_2232_),
    .ZN(_4478_));
 AOI21_X1 _7206_ (.A(_2186_),
    .B1(_2192_),
    .B2(net68),
    .ZN(_4482_));
 INV_X2 _7207_ (.A(_4485_),
    .ZN(_2280_));
 BUF_X2 _7208_ (.A(_4476_),
    .Z(_2281_));
 NOR3_X1 _7209_ (.A1(_2280_),
    .A2(_2273_),
    .A3(_2281_),
    .ZN(_2282_));
 AND3_X1 _7210_ (.A1(_4469_),
    .A2(_2272_),
    .A3(_2280_),
    .ZN(_2283_));
 MUX2_X1 _7211_ (.A(_2282_),
    .B(_2283_),
    .S(_2270_),
    .Z(_2284_));
 NOR4_X2 _7212_ (.A1(_4469_),
    .A2(_2280_),
    .A3(_2273_),
    .A4(_2281_),
    .ZN(_2285_));
 NOR3_X1 _7213_ (.A1(_2272_),
    .A2(_2280_),
    .A3(_2281_),
    .ZN(_2286_));
 NAND3_X1 _7214_ (.A1(_2272_),
    .A2(_2280_),
    .A3(_2273_),
    .ZN(_2287_));
 INV_X1 _7215_ (.A(_2281_),
    .ZN(_2288_));
 OAI21_X1 _7216_ (.A(_2287_),
    .B1(_2288_),
    .B2(_4485_),
    .ZN(_2289_));
 OR4_X4 _7217_ (.A1(_2284_),
    .A2(_2285_),
    .A3(_2286_),
    .A4(_2289_),
    .ZN(_4487_));
 AOI21_X1 _7218_ (.A(_2228_),
    .B1(_2227_),
    .B2(_4417_),
    .ZN(_4486_));
 NAND2_X1 _7219_ (.A1(_4425_),
    .A2(_2046_),
    .ZN(_2290_));
 OAI21_X2 _7220_ (.A(_2290_),
    .B1(_2185_),
    .B2(_2046_),
    .ZN(_2291_));
 XNOR2_X2 _7221_ (.A(net276),
    .B(_2291_),
    .ZN(_2292_));
 NAND2_X1 _7222_ (.A1(_2272_),
    .A2(_4485_),
    .ZN(_2293_));
 OR4_X1 _7223_ (.A1(_2275_),
    .A2(_2277_),
    .A3(_2292_),
    .A4(_2293_),
    .ZN(_2294_));
 XNOR2_X1 _7224_ (.A(_4259_),
    .B(_2291_),
    .ZN(_2295_));
 NOR2_X1 _7225_ (.A1(_2280_),
    .A2(_2288_),
    .ZN(_2296_));
 OAI21_X1 _7226_ (.A(_2295_),
    .B1(_2296_),
    .B2(_4484_),
    .ZN(_2297_));
 NOR2_X1 _7227_ (.A1(_2281_),
    .A2(_4484_),
    .ZN(_2298_));
 OAI211_X2 _7228_ (.A(_2292_),
    .B(_2298_),
    .C1(_2275_),
    .C2(_2277_),
    .ZN(_2299_));
 NOR3_X1 _7229_ (.A1(_2272_),
    .A2(_2281_),
    .A3(_4484_),
    .ZN(_2300_));
 NOR2_X1 _7230_ (.A1(_4485_),
    .A2(_4484_),
    .ZN(_2301_));
 OAI21_X1 _7231_ (.A(_2292_),
    .B1(_2300_),
    .B2(_2301_),
    .ZN(_2302_));
 AND4_X1 _7232_ (.A1(_2294_),
    .A2(_2297_),
    .A3(_2299_),
    .A4(_2302_),
    .ZN(_2303_));
 BUF_X4 _7233_ (.A(_2303_),
    .Z(_4523_));
 INV_X2 _7234_ (.A(_3012_),
    .ZN(_4497_));
 INV_X1 _7235_ (.A(net56),
    .ZN(_4498_));
 INV_X1 _7236_ (.A(_3149_),
    .ZN(_2912_));
 INV_X1 _7237_ (.A(_2921_),
    .ZN(_2936_));
 INV_X1 _7238_ (.A(_2953_),
    .ZN(_2960_));
 INV_X1 _7239_ (.A(_2991_),
    .ZN(_2993_));
 INV_X1 _7240_ (.A(net5),
    .ZN(_3013_));
 INV_X4 _7241_ (.A(net14),
    .ZN(_2896_));
 INV_X1 _7242_ (.A(net16),
    .ZN(_3027_));
 INV_X2 _7243_ (.A(net15),
    .ZN(_3035_));
 OAI21_X4 _7244_ (.A(_0002_),
    .B1(_0003_),
    .B2(_4502_),
    .ZN(_2304_));
 NAND2_X2 _7245_ (.A1(_3290_),
    .A2(_0205_),
    .ZN(_2305_));
 OR4_X4 _7246_ (.A1(net51),
    .A2(net50),
    .A3(_2305_),
    .A4(_0007_),
    .ZN(_2306_));
 NOR2_X4 _7247_ (.A1(_2306_),
    .A2(net52),
    .ZN(_2307_));
 AOI21_X4 _7248_ (.A(_2304_),
    .B1(_2307_),
    .B2(_0010_),
    .ZN(_2308_));
 NOR2_X1 _7249_ (.A1(_0009_),
    .A2(_2304_),
    .ZN(_2309_));
 OR2_X4 _7250_ (.A1(_2308_),
    .A2(_2309_),
    .ZN(_2310_));
 XNOR2_X2 _7251_ (.A(_2310_),
    .B(_4501_),
    .ZN(_2908_));
 INV_X1 _7252_ (.A(net20),
    .ZN(_3057_));
 INV_X1 _7253_ (.A(net19),
    .ZN(_3065_));
 INV_X1 _7254_ (.A(net21),
    .ZN(_3073_));
 AOI21_X2 _7255_ (.A(_2308_),
    .B1(_0042_),
    .B2(_0045_),
    .ZN(_2311_));
 XNOR2_X2 _7256_ (.A(net44),
    .B(_2311_),
    .ZN(_3105_));
 OAI21_X1 _7257_ (.A(_0042_),
    .B1(_0044_),
    .B2(net42),
    .ZN(_2312_));
 XNOR2_X2 _7258_ (.A(net43),
    .B(_2312_),
    .ZN(_3108_));
 XOR2_X2 _7259_ (.A(net42),
    .B(_2308_),
    .Z(_3111_));
 NOR2_X1 _7260_ (.A1(net54),
    .A2(net53),
    .ZN(_2313_));
 AOI21_X1 _7261_ (.A(_2304_),
    .B1(_2313_),
    .B2(_0043_),
    .ZN(_2314_));
 XOR2_X2 _7262_ (.A(net55),
    .B(_2314_),
    .Z(_3114_));
 INV_X1 _7263_ (.A(net53),
    .ZN(_2315_));
 AOI21_X1 _7264_ (.A(_2304_),
    .B1(_2307_),
    .B2(_2315_),
    .ZN(_2316_));
 XOR2_X2 _7265_ (.A(net54),
    .B(_2316_),
    .Z(_3117_));
 NOR2_X1 _7266_ (.A1(_0043_),
    .A2(_2304_),
    .ZN(_2317_));
 XNOR2_X1 _7267_ (.A(_2315_),
    .B(_2317_),
    .ZN(_3120_));
 NAND2_X1 _7268_ (.A1(_0042_),
    .A2(_2306_),
    .ZN(_2318_));
 XNOR2_X1 _7269_ (.A(net52),
    .B(_2318_),
    .ZN(_3123_));
 NOR2_X1 _7270_ (.A1(net50),
    .A2(_0007_),
    .ZN(_2319_));
 AOI21_X1 _7271_ (.A(_2304_),
    .B1(_2319_),
    .B2(_0006_),
    .ZN(_2320_));
 XOR2_X2 _7272_ (.A(net51),
    .B(_2320_),
    .Z(_3126_));
 OAI21_X1 _7273_ (.A(_0042_),
    .B1(_2305_),
    .B2(_0007_),
    .ZN(_2321_));
 XNOR2_X1 _7274_ (.A(net50),
    .B(_2321_),
    .ZN(_3129_));
 NOR2_X1 _7275_ (.A1(_0006_),
    .A2(_2304_),
    .ZN(_2322_));
 XOR2_X2 _7276_ (.A(_0007_),
    .B(_2322_),
    .Z(_2925_));
 OR2_X1 _7277_ (.A1(_2906_),
    .A2(_0015_),
    .ZN(_2323_));
 NOR2_X1 _7278_ (.A1(_0170_),
    .A2(_2323_),
    .ZN(_2324_));
 AOI21_X1 _7279_ (.A(_2324_),
    .B1(_0182_),
    .B2(_2909_),
    .ZN(_2325_));
 NOR2_X1 _7280_ (.A1(_0048_),
    .A2(_2325_),
    .ZN(_2326_));
 OAI22_X1 _7281_ (.A1(_0021_),
    .A2(_0186_),
    .B1(_2323_),
    .B2(_0037_),
    .ZN(_2327_));
 AOI21_X1 _7282_ (.A(_2326_),
    .B1(_2327_),
    .B2(_0048_),
    .ZN(_2328_));
 OAI21_X1 _7283_ (.A(_0191_),
    .B1(_3090_),
    .B2(_2328_),
    .ZN(_2329_));
 XNOR2_X1 _7284_ (.A(_3086_),
    .B(_2329_),
    .ZN(_3134_));
 NOR2_X1 _7285_ (.A1(_3147_),
    .A2(_3261_),
    .ZN(_2330_));
 XNOR2_X1 _7286_ (.A(_1178_),
    .B(_2330_),
    .ZN(_3142_));
 INV_X1 _7287_ (.A(net22),
    .ZN(_3157_));
 INV_X1 _7288_ (.A(net23),
    .ZN(_3165_));
 INV_X1 _7289_ (.A(net6),
    .ZN(_3181_));
 INV_X1 _7290_ (.A(net24),
    .ZN(_3189_));
 NOR2_X1 _7291_ (.A1(_3324_),
    .A2(_1047_),
    .ZN(_2331_));
 INV_X1 _7292_ (.A(_3050_),
    .ZN(_2332_));
 NOR2_X1 _7293_ (.A1(_0020_),
    .A2(_0175_),
    .ZN(_2333_));
 NOR3_X1 _7294_ (.A1(_2909_),
    .A2(_0031_),
    .A3(_0173_),
    .ZN(_2334_));
 NOR2_X1 _7295_ (.A1(_2333_),
    .A2(_2334_),
    .ZN(_2335_));
 NOR2_X4 _7296_ (.A1(_2332_),
    .A2(_2335_),
    .ZN(_2336_));
 AOI21_X1 _7297_ (.A(net227),
    .B1(_2331_),
    .B2(_2336_),
    .ZN(_2337_));
 XNOR2_X1 _7298_ (.A(_0395_),
    .B(_2337_),
    .ZN(_3201_));
 OAI21_X1 _7299_ (.A(_0191_),
    .B1(_1047_),
    .B2(_1052_),
    .ZN(_2338_));
 XNOR2_X1 _7300_ (.A(_3324_),
    .B(_2338_),
    .ZN(_3205_));
 NOR3_X1 _7301_ (.A1(_2909_),
    .A2(_0095_),
    .A3(_0323_),
    .ZN(_2339_));
 OAI21_X1 _7302_ (.A(_2336_),
    .B1(_2339_),
    .B2(_1045_),
    .ZN(_2340_));
 NAND2_X1 _7303_ (.A1(_0191_),
    .A2(_2340_),
    .ZN(_2341_));
 XNOR2_X1 _7304_ (.A(_3174_),
    .B(_2341_),
    .ZN(_3209_));
 OAI21_X1 _7305_ (.A(_0191_),
    .B1(_3082_),
    .B2(_1052_),
    .ZN(_2342_));
 XNOR2_X1 _7306_ (.A(_3178_),
    .B(_2342_),
    .ZN(_3213_));
 NOR2_X1 _7307_ (.A1(_2929_),
    .A2(_2336_),
    .ZN(_2343_));
 XOR2_X1 _7308_ (.A(_3082_),
    .B(_2343_),
    .Z(_3217_));
 INV_X1 _7309_ (.A(_3109_),
    .ZN(_2344_));
 INV_X1 _7310_ (.A(_3121_),
    .ZN(_2345_));
 INV_X1 _7311_ (.A(_3127_),
    .ZN(_2346_));
 AOI21_X1 _7312_ (.A(_3130_),
    .B1(_0227_),
    .B2(_2926_),
    .ZN(_2347_));
 INV_X1 _7313_ (.A(_3128_),
    .ZN(_2348_));
 OAI21_X1 _7314_ (.A(_2346_),
    .B1(_2347_),
    .B2(_2348_),
    .ZN(_2349_));
 AOI21_X1 _7315_ (.A(_3124_),
    .B1(_2349_),
    .B2(_3125_),
    .ZN(_2350_));
 INV_X1 _7316_ (.A(_0218_),
    .ZN(_2351_));
 OAI21_X2 _7317_ (.A(_2345_),
    .B1(_2350_),
    .B2(_2351_),
    .ZN(_2352_));
 AOI21_X1 _7318_ (.A(_3118_),
    .B1(_2352_),
    .B2(_0221_),
    .ZN(_2353_));
 OAI21_X2 _7319_ (.A(_0217_),
    .B1(_2353_),
    .B2(_0223_),
    .ZN(_2354_));
 AOI21_X1 _7320_ (.A(_3112_),
    .B1(_2354_),
    .B2(_0214_),
    .ZN(_2355_));
 OAI21_X2 _7321_ (.A(_2344_),
    .B1(_2355_),
    .B2(_0213_),
    .ZN(_2356_));
 AOI21_X1 _7322_ (.A(_3106_),
    .B1(_2356_),
    .B2(_0208_),
    .ZN(_2357_));
 INV_X1 _7323_ (.A(_2357_),
    .ZN(_2358_));
 AOI21_X1 _7324_ (.A(_3103_),
    .B1(_3104_),
    .B2(_2358_),
    .ZN(_2359_));
 XOR2_X2 _7325_ (.A(_0207_),
    .B(_2359_),
    .Z(_3251_));
 OR2_X1 _7326_ (.A1(_3109_),
    .A2(_1062_),
    .ZN(_2360_));
 AOI21_X1 _7327_ (.A(_3106_),
    .B1(_2360_),
    .B2(_0208_),
    .ZN(_2361_));
 XNOR2_X1 _7328_ (.A(_3104_),
    .B(_2361_),
    .ZN(_3254_));
 XOR2_X2 _7329_ (.A(_0208_),
    .B(_2356_),
    .Z(_3257_));
 NOR2_X1 _7330_ (.A1(_3110_),
    .A2(_3112_),
    .ZN(_2362_));
 NOR2_X1 _7331_ (.A1(_0231_),
    .A2(_0226_),
    .ZN(_2363_));
 OAI21_X1 _7332_ (.A(_0214_),
    .B1(_2363_),
    .B2(_0224_),
    .ZN(_2364_));
 AOI21_X1 _7333_ (.A(_1062_),
    .B1(_2362_),
    .B2(_2364_),
    .ZN(_3260_));
 XOR2_X2 _7334_ (.A(_0214_),
    .B(_2354_),
    .Z(_3264_));
 INV_X1 _7335_ (.A(_3125_),
    .ZN(_2365_));
 NOR2_X1 _7336_ (.A1(_2365_),
    .A2(_0231_),
    .ZN(_2366_));
 NAND3_X1 _7337_ (.A1(_0218_),
    .A2(_0221_),
    .A3(_2366_),
    .ZN(_2367_));
 NAND2_X1 _7338_ (.A1(_0222_),
    .A2(_2367_),
    .ZN(_2368_));
 XNOR2_X1 _7339_ (.A(_0223_),
    .B(_2368_),
    .ZN(_3267_));
 XOR2_X2 _7340_ (.A(_0221_),
    .B(_2352_),
    .Z(_3270_));
 NOR2_X1 _7341_ (.A1(_3124_),
    .A2(_2366_),
    .ZN(_2369_));
 XNOR2_X1 _7342_ (.A(_0218_),
    .B(_2369_),
    .ZN(_3273_));
 XNOR2_X1 _7343_ (.A(_2365_),
    .B(_2349_),
    .ZN(_3276_));
 XNOR2_X1 _7344_ (.A(_2348_),
    .B(_0230_),
    .ZN(_3279_));
 XOR2_X2 _7345_ (.A(_2926_),
    .B(_0227_),
    .Z(_3282_));
 INV_X1 _7346_ (.A(_3230_),
    .ZN(_2370_));
 NAND3_X1 _7347_ (.A1(_3147_),
    .A2(_2370_),
    .A3(_1178_),
    .ZN(_2371_));
 NAND2_X1 _7348_ (.A1(net224),
    .A2(_2371_),
    .ZN(_2372_));
 XNOR2_X1 _7349_ (.A(_3226_),
    .B(_2372_),
    .ZN(_3295_));
 AND2_X1 _7350_ (.A1(_0476_),
    .A2(_1196_),
    .ZN(_2373_));
 NOR2_X1 _7351_ (.A1(_3483_),
    .A2(_2373_),
    .ZN(_2374_));
 XNOR2_X1 _7352_ (.A(_1195_),
    .B(_2374_),
    .ZN(_3303_));
 XOR2_X2 _7353_ (.A(_3144_),
    .B(_2932_),
    .Z(_3306_));
 INV_X1 _7354_ (.A(net8),
    .ZN(_3327_));
 INV_X1 _7355_ (.A(net7),
    .ZN(_3335_));
 AND2_X1 _7356_ (.A1(_0395_),
    .A2(_2331_),
    .ZN(_2375_));
 INV_X1 _7357_ (.A(_2375_),
    .ZN(_2376_));
 NOR2_X1 _7358_ (.A1(_3388_),
    .A2(_2376_),
    .ZN(_2377_));
 AOI21_X2 _7359_ (.A(_0053_),
    .B1(_2377_),
    .B2(_2336_),
    .ZN(_2378_));
 XOR2_X2 _7360_ (.A(_3392_),
    .B(_2378_),
    .Z(_3347_));
 INV_X1 _7361_ (.A(net12),
    .ZN(_3359_));
 INV_X1 _7362_ (.A(net11),
    .ZN(_3367_));
 INV_X1 _7363_ (.A(_2336_),
    .ZN(_2379_));
 OAI21_X1 _7364_ (.A(_0191_),
    .B1(_1055_),
    .B2(_2379_),
    .ZN(_2380_));
 XNOR2_X1 _7365_ (.A(_3380_),
    .B(_2380_),
    .ZN(_3395_));
 NOR2_X1 _7366_ (.A1(net17),
    .A2(_1182_),
    .ZN(_2381_));
 XNOR2_X1 _7367_ (.A(_1177_),
    .B(_2381_),
    .ZN(_3403_));
 NOR2_X1 _7368_ (.A1(_3546_),
    .A2(_3550_),
    .ZN(_2382_));
 OR3_X1 _7369_ (.A1(_3222_),
    .A2(_3226_),
    .A3(_2371_),
    .ZN(_2383_));
 OR3_X1 _7370_ (.A1(_3352_),
    .A2(_3356_),
    .A3(_2383_),
    .ZN(_2384_));
 INV_X1 _7371_ (.A(_2384_),
    .ZN(_2385_));
 AOI21_X1 _7372_ (.A(_0235_),
    .B1(_2382_),
    .B2(_2385_),
    .ZN(_2386_));
 XNOR2_X1 _7373_ (.A(_0774_),
    .B(_2386_),
    .ZN(_3407_));
 OAI21_X1 _7374_ (.A(net224),
    .B1(_3550_),
    .B2(_1181_),
    .ZN(_2387_));
 XNOR2_X1 _7375_ (.A(_3546_),
    .B(_2387_),
    .ZN(_3411_));
 NAND2_X1 _7376_ (.A1(net224),
    .A2(_2384_),
    .ZN(_2388_));
 XNOR2_X1 _7377_ (.A(_3550_),
    .B(_2388_),
    .ZN(_3415_));
 NAND3_X1 _7378_ (.A1(_0340_),
    .A2(_0621_),
    .A3(_1180_),
    .ZN(_2389_));
 NAND2_X1 _7379_ (.A1(net224),
    .A2(_2389_),
    .ZN(_2390_));
 XNOR2_X1 _7380_ (.A(_3352_),
    .B(_2390_),
    .ZN(_3419_));
 NAND2_X1 _7381_ (.A1(net224),
    .A2(_2383_),
    .ZN(_2391_));
 XNOR2_X1 _7382_ (.A(_3356_),
    .B(_2391_),
    .ZN(_3423_));
 NOR2_X1 _7383_ (.A1(net17),
    .A2(_1180_),
    .ZN(_2392_));
 XNOR2_X1 _7384_ (.A(_0340_),
    .B(_2392_),
    .ZN(_3427_));
 INV_X1 _7385_ (.A(_3258_),
    .ZN(_2393_));
 INV_X1 _7386_ (.A(_3265_),
    .ZN(_2394_));
 INV_X1 _7387_ (.A(_3271_),
    .ZN(_2395_));
 INV_X1 _7388_ (.A(_3277_),
    .ZN(_2396_));
 OAI21_X1 _7389_ (.A(_0495_),
    .B1(_0497_),
    .B2(_2943_),
    .ZN(_2397_));
 AOI21_X1 _7390_ (.A(_3285_),
    .B1(_2397_),
    .B2(_3286_),
    .ZN(_2398_));
 OAI21_X1 _7391_ (.A(_0494_),
    .B1(_2398_),
    .B2(_0500_),
    .ZN(_2399_));
 AOI21_X2 _7392_ (.A(_3280_),
    .B1(_2399_),
    .B2(_3281_),
    .ZN(_2400_));
 OAI21_X1 _7393_ (.A(_2396_),
    .B1(_2400_),
    .B2(_0503_),
    .ZN(_2401_));
 AOI21_X1 _7394_ (.A(_3274_),
    .B1(_2401_),
    .B2(_3275_),
    .ZN(_2402_));
 INV_X1 _7395_ (.A(_3272_),
    .ZN(_2403_));
 OAI21_X1 _7396_ (.A(_2395_),
    .B1(_2402_),
    .B2(_2403_),
    .ZN(_2404_));
 AOI21_X2 _7397_ (.A(_3268_),
    .B1(_2404_),
    .B2(_3269_),
    .ZN(_2405_));
 INV_X1 _7398_ (.A(_3266_),
    .ZN(_2406_));
 OAI21_X1 _7399_ (.A(_2394_),
    .B1(_2405_),
    .B2(_2406_),
    .ZN(_2407_));
 AOI21_X1 _7400_ (.A(_3262_),
    .B1(_2407_),
    .B2(_0508_),
    .ZN(_2408_));
 INV_X1 _7401_ (.A(_0509_),
    .ZN(_2409_));
 OAI21_X1 _7402_ (.A(_2393_),
    .B1(_2408_),
    .B2(_2409_),
    .ZN(_2410_));
 AOI21_X1 _7403_ (.A(_3255_),
    .B1(_2410_),
    .B2(_3256_),
    .ZN(_2411_));
 XNOR2_X1 _7404_ (.A(_3253_),
    .B(_2411_),
    .ZN(_3469_));
 NOR2_X1 _7405_ (.A1(_0505_),
    .A2(_0507_),
    .ZN(_2412_));
 AOI21_X1 _7406_ (.A(_3262_),
    .B1(_2412_),
    .B2(_0508_),
    .ZN(_2413_));
 OAI21_X1 _7407_ (.A(_2393_),
    .B1(_2413_),
    .B2(_2409_),
    .ZN(_2414_));
 XNOR2_X1 _7408_ (.A(_0514_),
    .B(_2414_),
    .ZN(_3473_));
 XNOR2_X1 _7409_ (.A(_0509_),
    .B(_2408_),
    .ZN(_3476_));
 XOR2_X2 _7410_ (.A(_0508_),
    .B(_2412_),
    .Z(_3479_));
 XNOR2_X1 _7411_ (.A(_3266_),
    .B(_2405_),
    .ZN(_3482_));
 AOI21_X1 _7412_ (.A(_3271_),
    .B1(_0504_),
    .B2(_0492_),
    .ZN(_2415_));
 XNOR2_X1 _7413_ (.A(_3269_),
    .B(_2415_),
    .ZN(_3486_));
 XNOR2_X1 _7414_ (.A(_3272_),
    .B(_2402_),
    .ZN(_3489_));
 NOR2_X1 _7415_ (.A1(_0503_),
    .A2(_0502_),
    .ZN(_2416_));
 NOR2_X1 _7416_ (.A1(_3277_),
    .A2(_2416_),
    .ZN(_2417_));
 XNOR2_X1 _7417_ (.A(_3275_),
    .B(_2417_),
    .ZN(_3492_));
 XNOR2_X1 _7418_ (.A(_3278_),
    .B(_2400_),
    .ZN(_3495_));
 XOR2_X2 _7419_ (.A(_3281_),
    .B(_0501_),
    .Z(_3498_));
 XNOR2_X1 _7420_ (.A(_3284_),
    .B(_2398_),
    .ZN(_3501_));
 XOR2_X2 _7421_ (.A(_3286_),
    .B(_0498_),
    .Z(_3504_));
 XNOR2_X1 _7422_ (.A(_2943_),
    .B(_3288_),
    .ZN(_3507_));
 INV_X1 _7423_ (.A(_2944_),
    .ZN(_3510_));
 OR2_X1 _7424_ (.A1(_3444_),
    .A2(_1197_),
    .ZN(_2418_));
 AND2_X1 _7425_ (.A1(net9),
    .A2(_2418_),
    .ZN(_2419_));
 XNOR2_X1 _7426_ (.A(_0905_),
    .B(_2419_),
    .ZN(_3513_));
 AND3_X1 _7427_ (.A1(_3534_),
    .A2(_0916_),
    .A3(_0917_),
    .ZN(_2420_));
 NOR2_X1 _7428_ (.A1(_3686_),
    .A2(_2420_),
    .ZN(_2421_));
 XNOR2_X1 _7429_ (.A(_1322_),
    .B(_2421_),
    .ZN(_3521_));
 XNOR2_X1 _7430_ (.A(_0526_),
    .B(_0910_),
    .ZN(_3524_));
 XOR2_X2 _7431_ (.A(_2947_),
    .B(_3309_),
    .Z(_3528_));
 OR2_X2 _7432_ (.A1(_3380_),
    .A2(_1055_),
    .ZN(_2422_));
 OAI21_X2 _7433_ (.A(_0191_),
    .B1(_2422_),
    .B2(_1052_),
    .ZN(_2423_));
 XNOR2_X1 _7434_ (.A(_3376_),
    .B(_2423_),
    .ZN(_3541_));
 NOR3_X4 _7435_ (.A1(_3376_),
    .A2(_2422_),
    .A3(_2379_),
    .ZN(_2424_));
 NOR2_X2 _7436_ (.A1(net227),
    .A2(_2424_),
    .ZN(_2425_));
 XNOR2_X2 _7437_ (.A(_1040_),
    .B(_2425_),
    .ZN(_3553_));
 XNOR2_X1 _7438_ (.A(_1185_),
    .B(_1184_),
    .ZN(_3561_));
 NOR2_X4 _7439_ (.A1(_3746_),
    .A2(_3762_),
    .ZN(_2426_));
 AND3_X1 _7440_ (.A1(_3312_),
    .A2(_0476_),
    .A3(_1195_),
    .ZN(_2427_));
 NAND3_X1 _7441_ (.A1(_0488_),
    .A2(_0905_),
    .A3(_2427_),
    .ZN(_2428_));
 OR3_X1 _7442_ (.A1(_3432_),
    .A2(_3570_),
    .A3(_2428_),
    .ZN(_2429_));
 NOR3_X2 _7443_ (.A1(_3566_),
    .A2(_3750_),
    .A3(_2429_),
    .ZN(_2430_));
 AOI21_X2 _7444_ (.A(_0519_),
    .B1(_2426_),
    .B2(_2430_),
    .ZN(_2431_));
 NAND2_X1 _7445_ (.A1(_1239_),
    .A2(_2431_),
    .ZN(_2432_));
 NAND2_X1 _7446_ (.A1(_1367_),
    .A2(_2432_),
    .ZN(_3585_));
 XNOR2_X2 _7447_ (.A(_2431_),
    .B(_1239_),
    .ZN(_3589_));
 NOR2_X1 _7448_ (.A1(_0519_),
    .A2(_2430_),
    .ZN(_2433_));
 XOR2_X2 _7449_ (.A(_3746_),
    .B(_2433_),
    .Z(_3595_));
 NAND2_X1 _7450_ (.A1(_0947_),
    .A2(_1199_),
    .ZN(_2434_));
 NAND2_X1 _7451_ (.A1(net9),
    .A2(_2434_),
    .ZN(_2435_));
 XNOR2_X1 _7452_ (.A(_3750_),
    .B(_2435_),
    .ZN(_3599_));
 NAND2_X1 _7453_ (.A1(net9),
    .A2(_2429_),
    .ZN(_2436_));
 XNOR2_X1 _7454_ (.A(_3566_),
    .B(_2436_),
    .ZN(_3603_));
 OAI21_X1 _7455_ (.A(net9),
    .B1(_2418_),
    .B2(_1198_),
    .ZN(_2437_));
 XNOR2_X1 _7456_ (.A(_3570_),
    .B(_2437_),
    .ZN(_3607_));
 NAND2_X1 _7457_ (.A1(net9),
    .A2(_2428_),
    .ZN(_2438_));
 XNOR2_X1 _7458_ (.A(_3432_),
    .B(_2438_),
    .ZN(_3611_));
 NAND2_X1 _7459_ (.A1(_1231_),
    .A2(_1367_),
    .ZN(_3615_));
 OAI21_X1 _7460_ (.A(net9),
    .B1(_3746_),
    .B2(_1200_),
    .ZN(_2439_));
 XNOR2_X1 _7461_ (.A(_3762_),
    .B(_2439_),
    .ZN(_3619_));
 INV_X1 _7462_ (.A(_3477_),
    .ZN(_2440_));
 INV_X1 _7463_ (.A(_3481_),
    .ZN(_2441_));
 INV_X1 _7464_ (.A(_3488_),
    .ZN(_2442_));
 INV_X1 _7465_ (.A(_3490_),
    .ZN(_2443_));
 INV_X1 _7466_ (.A(_3497_),
    .ZN(_2444_));
 INV_X1 _7467_ (.A(_3502_),
    .ZN(_2445_));
 INV_X1 _7468_ (.A(_3508_),
    .ZN(_2446_));
 MUX2_X1 _7469_ (.A(_0519_),
    .B(_1769_),
    .S(_3294_),
    .Z(_2447_));
 INV_X1 _7470_ (.A(_3509_),
    .ZN(_2448_));
 OAI21_X1 _7471_ (.A(_2446_),
    .B1(_2447_),
    .B2(_2448_),
    .ZN(_2449_));
 AOI21_X2 _7472_ (.A(_3505_),
    .B1(_2449_),
    .B2(_0886_),
    .ZN(_2450_));
 INV_X1 _7473_ (.A(_3503_),
    .ZN(_2451_));
 OAI21_X1 _7474_ (.A(_2445_),
    .B1(_2450_),
    .B2(_2451_),
    .ZN(_2452_));
 NAND2_X1 _7475_ (.A1(_0890_),
    .A2(_2452_),
    .ZN(_2453_));
 AOI21_X1 _7476_ (.A(_2444_),
    .B1(_0880_),
    .B2(_2453_),
    .ZN(_2454_));
 OAI21_X1 _7477_ (.A(_3494_),
    .B1(_3496_),
    .B2(_2454_),
    .ZN(_2455_));
 INV_X1 _7478_ (.A(_2455_),
    .ZN(_2456_));
 OAI21_X1 _7479_ (.A(_0877_),
    .B1(_3493_),
    .B2(_2456_),
    .ZN(_2457_));
 AOI21_X1 _7480_ (.A(_2442_),
    .B1(_2443_),
    .B2(_2457_),
    .ZN(_2458_));
 OAI21_X1 _7481_ (.A(_3485_),
    .B1(_3487_),
    .B2(_2458_),
    .ZN(_2459_));
 AOI21_X1 _7482_ (.A(_2441_),
    .B1(_0876_),
    .B2(_2459_),
    .ZN(_2460_));
 OAI21_X1 _7483_ (.A(_3478_),
    .B1(_3480_),
    .B2(_2460_),
    .ZN(_2461_));
 NAND2_X1 _7484_ (.A1(_2440_),
    .A2(_2461_),
    .ZN(_2462_));
 AOI21_X1 _7485_ (.A(_3474_),
    .B1(_2462_),
    .B2(_3475_),
    .ZN(_2463_));
 XNOR2_X1 _7486_ (.A(_3472_),
    .B(_2463_),
    .ZN(_3669_));
 INV_X1 _7487_ (.A(_3480_),
    .ZN(_2464_));
 INV_X1 _7488_ (.A(_3487_),
    .ZN(_2465_));
 INV_X1 _7489_ (.A(_0878_),
    .ZN(_2466_));
 AND2_X1 _7490_ (.A1(_0877_),
    .A2(_3494_),
    .ZN(_2467_));
 INV_X1 _7491_ (.A(_3496_),
    .ZN(_2468_));
 AOI21_X1 _7492_ (.A(_3511_),
    .B1(_3512_),
    .B2(_2940_),
    .ZN(_2469_));
 OAI21_X1 _7493_ (.A(_2446_),
    .B1(_2469_),
    .B2(_2448_),
    .ZN(_2470_));
 AOI21_X1 _7494_ (.A(_3505_),
    .B1(_2470_),
    .B2(_0886_),
    .ZN(_2471_));
 OAI21_X1 _7495_ (.A(_2445_),
    .B1(_2471_),
    .B2(_2451_),
    .ZN(_2472_));
 AOI21_X1 _7496_ (.A(_3499_),
    .B1(_2472_),
    .B2(_0890_),
    .ZN(_2473_));
 OAI21_X1 _7497_ (.A(_2468_),
    .B1(_2473_),
    .B2(_2444_),
    .ZN(_2474_));
 AOI21_X2 _7498_ (.A(_2466_),
    .B1(_2467_),
    .B2(_2474_),
    .ZN(_2475_));
 OAI21_X1 _7499_ (.A(_2465_),
    .B1(_2475_),
    .B2(_2442_),
    .ZN(_2476_));
 AOI21_X2 _7500_ (.A(_3484_),
    .B1(_2476_),
    .B2(_3485_),
    .ZN(_2477_));
 OAI21_X1 _7501_ (.A(_2464_),
    .B1(_2477_),
    .B2(_2441_),
    .ZN(_2478_));
 AOI21_X1 _7502_ (.A(_3477_),
    .B1(_2478_),
    .B2(_3478_),
    .ZN(_2479_));
 XNOR2_X1 _7503_ (.A(_3475_),
    .B(_2479_),
    .ZN(_3673_));
 OR3_X1 _7504_ (.A1(_3478_),
    .A2(_3480_),
    .A3(_2460_),
    .ZN(_2480_));
 AND2_X1 _7505_ (.A1(_2461_),
    .A2(_2480_),
    .ZN(_3676_));
 XNOR2_X1 _7506_ (.A(_3481_),
    .B(_2477_),
    .ZN(_3679_));
 OR3_X1 _7507_ (.A1(_3485_),
    .A2(_3487_),
    .A3(_2458_),
    .ZN(_2481_));
 AND2_X1 _7508_ (.A1(_2459_),
    .A2(_2481_),
    .ZN(_3682_));
 XNOR2_X1 _7509_ (.A(_3488_),
    .B(_2475_),
    .ZN(_3685_));
 OR3_X1 _7510_ (.A1(_0877_),
    .A2(_3493_),
    .A3(_2456_),
    .ZN(_2482_));
 AND2_X1 _7511_ (.A1(_2457_),
    .A2(_2482_),
    .ZN(_3689_));
 XNOR2_X1 _7512_ (.A(_3494_),
    .B(_0893_),
    .ZN(_3692_));
 NAND2_X1 _7513_ (.A1(_0880_),
    .A2(_2453_),
    .ZN(_2483_));
 XNOR2_X1 _7514_ (.A(_2444_),
    .B(_2483_),
    .ZN(_3695_));
 XNOR2_X1 _7515_ (.A(_0890_),
    .B(_0889_),
    .ZN(_3698_));
 XNOR2_X1 _7516_ (.A(_3503_),
    .B(_2450_),
    .ZN(_3701_));
 XNOR2_X1 _7517_ (.A(_0886_),
    .B(_0885_),
    .ZN(_3704_));
 XNOR2_X1 _7518_ (.A(_3509_),
    .B(_2447_),
    .ZN(_3707_));
 XNOR2_X1 _7519_ (.A(_1769_),
    .B(_3512_),
    .ZN(_3710_));
 INV_X1 _7520_ (.A(_3666_),
    .ZN(_2484_));
 NAND3_X1 _7521_ (.A1(_2484_),
    .A2(_1322_),
    .A3(_2420_),
    .ZN(_2485_));
 NAND2_X1 _7522_ (.A1(_3670_),
    .A2(_2485_),
    .ZN(_2486_));
 XNOR2_X1 _7523_ (.A(_3628_),
    .B(_2486_),
    .ZN(_3713_));
 NOR2_X1 _7524_ (.A1(_3810_),
    .A2(_3814_),
    .ZN(_2487_));
 AOI21_X1 _7525_ (.A(net226),
    .B1(_1679_),
    .B2(_2487_),
    .ZN(_2488_));
 XOR2_X2 _7526_ (.A(_3804_),
    .B(_2488_),
    .Z(_3721_));
 XNOR2_X1 _7527_ (.A(_0924_),
    .B(_1328_),
    .ZN(_3724_));
 XNOR2_X1 _7528_ (.A(_1327_),
    .B(_0922_),
    .ZN(_3728_));
 XOR2_X2 _7529_ (.A(_3531_),
    .B(_2956_),
    .Z(_3732_));
 NAND2_X2 _7530_ (.A1(_1460_),
    .A2(_1461_),
    .ZN(_2489_));
 NOR3_X1 _7531_ (.A1(_3624_),
    .A2(_3628_),
    .A3(_2485_),
    .ZN(_2490_));
 INV_X1 _7532_ (.A(_2490_),
    .ZN(_2491_));
 NOR3_X1 _7533_ (.A1(_3754_),
    .A2(_3758_),
    .A3(_2491_),
    .ZN(_2492_));
 AOI21_X1 _7534_ (.A(net219),
    .B1(_1466_),
    .B2(_2492_),
    .ZN(_2493_));
 NAND2_X1 _7535_ (.A1(_2489_),
    .A2(_2493_),
    .ZN(_2494_));
 NAND2_X1 _7536_ (.A1(_1476_),
    .A2(_2494_),
    .ZN(_3765_));
 NAND2_X1 _7537_ (.A1(_1476_),
    .A2(_2494_),
    .ZN(_3769_));
 NOR2_X1 _7538_ (.A1(net228),
    .A2(_2492_),
    .ZN(_2495_));
 XNOR2_X1 _7539_ (.A(_1466_),
    .B(_2495_),
    .ZN(_3775_));
 NOR3_X1 _7540_ (.A1(_3624_),
    .A2(_3758_),
    .A3(_1464_),
    .ZN(_2496_));
 NOR2_X1 _7541_ (.A1(net219),
    .A2(_2496_),
    .ZN(_2497_));
 XOR2_X2 _7542_ (.A(_3754_),
    .B(_2497_),
    .Z(_3779_));
 NOR2_X1 _7543_ (.A1(_0901_),
    .A2(_2490_),
    .ZN(_2498_));
 XOR2_X2 _7544_ (.A(_3758_),
    .B(_2498_),
    .Z(_3783_));
 NAND2_X1 _7545_ (.A1(_3670_),
    .A2(_1464_),
    .ZN(_2499_));
 XNOR2_X1 _7546_ (.A(_3624_),
    .B(_2499_),
    .ZN(_3787_));
 NAND2_X1 _7547_ (.A1(_1476_),
    .A2(_1478_),
    .ZN(_3791_));
 XNOR2_X1 _7548_ (.A(_2489_),
    .B(_1477_),
    .ZN(_3795_));
 INV_X1 _7549_ (.A(_2962_),
    .ZN(_2972_));
 INV_X1 _7550_ (.A(_3680_),
    .ZN(_2500_));
 INV_X1 _7551_ (.A(_3687_),
    .ZN(_2501_));
 INV_X1 _7552_ (.A(_3693_),
    .ZN(_2502_));
 INV_X1 _7553_ (.A(_3699_),
    .ZN(_2503_));
 INV_X1 _7554_ (.A(_3705_),
    .ZN(_2504_));
 MUX2_X1 _7555_ (.A(_1769_),
    .B(net219),
    .S(_0883_),
    .Z(_2505_));
 AOI21_X1 _7556_ (.A(_3708_),
    .B1(_2505_),
    .B2(_3709_),
    .ZN(_2506_));
 INV_X1 _7557_ (.A(_3706_),
    .ZN(_2507_));
 OAI21_X1 _7558_ (.A(_2504_),
    .B1(_2506_),
    .B2(_2507_),
    .ZN(_2508_));
 AOI21_X1 _7559_ (.A(_3702_),
    .B1(_2508_),
    .B2(_3703_),
    .ZN(_2509_));
 INV_X1 _7560_ (.A(_3700_),
    .ZN(_2510_));
 OAI21_X1 _7561_ (.A(_2503_),
    .B1(_2509_),
    .B2(_2510_),
    .ZN(_2511_));
 AOI21_X1 _7562_ (.A(_3696_),
    .B1(_2511_),
    .B2(_3697_),
    .ZN(_2512_));
 INV_X1 _7563_ (.A(_3694_),
    .ZN(_2513_));
 OAI21_X1 _7564_ (.A(_2502_),
    .B1(_2512_),
    .B2(_2513_),
    .ZN(_2514_));
 AOI21_X1 _7565_ (.A(_3690_),
    .B1(_2514_),
    .B2(_3691_),
    .ZN(_2515_));
 INV_X1 _7566_ (.A(_3688_),
    .ZN(_2516_));
 OAI21_X1 _7567_ (.A(_2501_),
    .B1(_2515_),
    .B2(_2516_),
    .ZN(_2517_));
 AOI21_X1 _7568_ (.A(_3683_),
    .B1(_2517_),
    .B2(_3684_),
    .ZN(_2518_));
 INV_X1 _7569_ (.A(_3681_),
    .ZN(_2519_));
 OAI21_X1 _7570_ (.A(_2500_),
    .B1(_2518_),
    .B2(_2519_),
    .ZN(_2520_));
 NAND2_X1 _7571_ (.A1(_3678_),
    .A2(_2520_),
    .ZN(_2521_));
 NAND2_X1 _7572_ (.A1(_1293_),
    .A2(_2521_),
    .ZN(_2522_));
 AOI21_X1 _7573_ (.A(_3674_),
    .B1(_2522_),
    .B2(_3675_),
    .ZN(_2523_));
 XNOR2_X1 _7574_ (.A(_3672_),
    .B(_2523_),
    .ZN(_3855_));
 XOR2_X2 _7575_ (.A(_3675_),
    .B(_1316_),
    .Z(_3859_));
 XNOR2_X1 _7576_ (.A(_1315_),
    .B(_2520_),
    .ZN(_3862_));
 XNOR2_X1 _7577_ (.A(_2519_),
    .B(_1313_),
    .ZN(_3865_));
 XNOR2_X1 _7578_ (.A(_1312_),
    .B(_2517_),
    .ZN(_3868_));
 XNOR2_X1 _7579_ (.A(_2516_),
    .B(_1310_),
    .ZN(_3871_));
 XNOR2_X1 _7580_ (.A(_1309_),
    .B(_2514_),
    .ZN(_3874_));
 XNOR2_X1 _7581_ (.A(_2513_),
    .B(_1307_),
    .ZN(_3878_));
 XNOR2_X1 _7582_ (.A(_1306_),
    .B(_2511_),
    .ZN(_3881_));
 XNOR2_X1 _7583_ (.A(_2510_),
    .B(_1304_),
    .ZN(_3884_));
 XNOR2_X1 _7584_ (.A(_1303_),
    .B(_2508_),
    .ZN(_3887_));
 XNOR2_X1 _7585_ (.A(_2507_),
    .B(_1301_),
    .ZN(_3890_));
 XNOR2_X1 _7586_ (.A(_1300_),
    .B(_2505_),
    .ZN(_3893_));
 XOR2_X2 _7587_ (.A(_1769_),
    .B(_3712_),
    .Z(_3896_));
 NAND2_X1 _7588_ (.A1(net1),
    .A2(_1682_),
    .ZN(_2524_));
 XNOR2_X1 _7589_ (.A(_3847_),
    .B(_2524_),
    .ZN(_3899_));
 OAI21_X1 _7590_ (.A(net4),
    .B1(_1866_),
    .B2(_1869_),
    .ZN(_2525_));
 XNOR2_X1 _7591_ (.A(_4015_),
    .B(_2525_),
    .ZN(_3903_));
 NAND2_X1 _7592_ (.A1(_3928_),
    .A2(_1865_),
    .ZN(_2526_));
 OAI21_X1 _7593_ (.A(_1657_),
    .B1(_1868_),
    .B2(_2526_),
    .ZN(_2527_));
 XNOR2_X1 _7594_ (.A(_4019_),
    .B(_2527_),
    .ZN(_3907_));
 XNOR2_X2 _7595_ (.A(_1346_),
    .B(_1600_),
    .ZN(_3910_));
 XNOR2_X2 _7596_ (.A(_1599_),
    .B(_1344_),
    .ZN(_3914_));
 XNOR2_X2 _7597_ (.A(_1343_),
    .B(_1597_),
    .ZN(_3918_));
 XOR2_X2 _7598_ (.A(_2966_),
    .B(_3735_),
    .Z(_3922_));
 NOR2_X4 _7599_ (.A1(_1697_),
    .A2(_1698_),
    .ZN(_2528_));
 INV_X1 _7600_ (.A(_3738_),
    .ZN(_2529_));
 NOR2_X1 _7601_ (.A1(_2529_),
    .A2(_3818_),
    .ZN(_2530_));
 NAND2_X1 _7602_ (.A1(_1680_),
    .A2(_2530_),
    .ZN(_2531_));
 NOR3_X1 _7603_ (.A1(_3852_),
    .A2(_3847_),
    .A3(_2531_),
    .ZN(_2532_));
 NOR2_X1 _7604_ (.A1(_3799_),
    .A2(_3939_),
    .ZN(_2533_));
 AOI21_X1 _7605_ (.A(net226),
    .B1(_2532_),
    .B2(_2533_),
    .ZN(_2534_));
 NAND2_X1 _7606_ (.A1(_2528_),
    .A2(_2534_),
    .ZN(_2535_));
 NAND2_X1 _7607_ (.A1(_1699_),
    .A2(_2535_),
    .ZN(_3943_));
 NAND2_X1 _7608_ (.A1(_1695_),
    .A2(_1699_),
    .ZN(_3947_));
 XNOR2_X2 _7609_ (.A(_2528_),
    .B(_2534_),
    .ZN(_3955_));
 NOR2_X1 _7610_ (.A1(net229),
    .A2(_1683_),
    .ZN(_2536_));
 XNOR2_X1 _7611_ (.A(_1621_),
    .B(_2536_),
    .ZN(_3959_));
 NOR2_X1 _7612_ (.A1(net226),
    .A2(_2532_),
    .ZN(_2537_));
 XOR2_X2 _7613_ (.A(_3799_),
    .B(_2537_),
    .Z(_3963_));
 NAND2_X1 _7614_ (.A1(_1699_),
    .A2(_2535_),
    .ZN(_3951_));
 NAND2_X2 _7615_ (.A1(_1695_),
    .A2(_1699_),
    .ZN(_3969_));
 XNOR2_X1 _7616_ (.A(_3836_),
    .B(_1522_),
    .ZN(_4001_));
 INV_X1 _7617_ (.A(_2971_),
    .ZN(_2978_));
 INV_X1 _7618_ (.A(_3885_),
    .ZN(_2538_));
 INV_X1 _7619_ (.A(_3891_),
    .ZN(_2539_));
 MUX2_X1 _7620_ (.A(_1320_),
    .B(_1769_),
    .S(_3712_),
    .Z(_2540_));
 OAI21_X1 _7621_ (.A(_1568_),
    .B1(_2540_),
    .B2(_1571_),
    .ZN(_2541_));
 NAND2_X1 _7622_ (.A1(_3892_),
    .A2(_2541_),
    .ZN(_2542_));
 AOI21_X1 _7623_ (.A(_1574_),
    .B1(_2539_),
    .B2(_2542_),
    .ZN(_2543_));
 OAI21_X1 _7624_ (.A(_3886_),
    .B1(_3888_),
    .B2(_2543_),
    .ZN(_2544_));
 NAND2_X1 _7625_ (.A1(_2538_),
    .A2(_2544_),
    .ZN(_2545_));
 XNOR2_X1 _7626_ (.A(_1577_),
    .B(_2545_),
    .ZN(_4057_));
 XNOR2_X1 _7627_ (.A(_1769_),
    .B(_1569_),
    .ZN(_4072_));
 XNOR2_X1 _7628_ (.A(_1614_),
    .B(_1800_),
    .ZN(_4083_));
 OAI21_X1 _7629_ (.A(_1791_),
    .B1(_2172_),
    .B2(_4186_),
    .ZN(_2546_));
 XNOR2_X1 _7630_ (.A(_4183_),
    .B(_2546_),
    .ZN(_4087_));
 NOR2_X1 _7631_ (.A1(_4142_),
    .A2(_4190_),
    .ZN(_2547_));
 NAND2_X1 _7632_ (.A1(_4105_),
    .A2(_2547_),
    .ZN(_2548_));
 NAND2_X1 _7633_ (.A1(_4198_),
    .A2(_2548_),
    .ZN(_2549_));
 XNOR2_X1 _7634_ (.A(_4186_),
    .B(_2549_),
    .ZN(_4091_));
 NAND2_X1 _7635_ (.A1(_1791_),
    .A2(_2171_),
    .ZN(_2550_));
 XNOR2_X1 _7636_ (.A(_4142_),
    .B(_2550_),
    .ZN(_4095_));
 NOR2_X2 _7637_ (.A1(_4105_),
    .A2(_4223_),
    .ZN(_2551_));
 XNOR2_X1 _7638_ (.A(_2170_),
    .B(_2551_),
    .ZN(_4099_));
 MUX2_X1 _7639_ (.A(_4146_),
    .B(_4106_),
    .S(_4198_),
    .Z(_2985_));
 XOR2_X2 _7640_ (.A(_3992_),
    .B(_1733_),
    .Z(_4150_));
 XNOR2_X1 _7641_ (.A(_3996_),
    .B(_1752_),
    .ZN(_4156_));
 XNOR2_X1 _7642_ (.A(_4004_),
    .B(_1750_),
    .ZN(_4164_));
 XOR2_X2 _7643_ (.A(_2981_),
    .B(net127),
    .Z(_4168_));
 NOR2_X4 _7644_ (.A1(_2002_),
    .A2(_2001_),
    .ZN(_2552_));
 OR2_X1 _7645_ (.A1(_2173_),
    .A2(_2548_),
    .ZN(_2553_));
 NOR3_X1 _7646_ (.A1(_4139_),
    .A2(_4179_),
    .A3(_2553_),
    .ZN(_2554_));
 NOR2_X1 _7647_ (.A1(_4223_),
    .A2(_2554_),
    .ZN(_2555_));
 XNOR2_X2 _7648_ (.A(_2555_),
    .B(_2552_),
    .ZN(_4079_));
 NAND2_X1 _7649_ (.A1(net3),
    .A2(_2174_),
    .ZN(_2556_));
 XNOR2_X1 _7650_ (.A(_4139_),
    .B(_2556_),
    .ZN(_4248_));
 NOR2_X1 _7651_ (.A1(_4335_),
    .A2(_2056_),
    .ZN(_2557_));
 XNOR2_X1 _7652_ (.A(_1951_),
    .B(_2557_),
    .ZN(_4262_));
 XNOR2_X2 _7653_ (.A(_1808_),
    .B(_2020_),
    .ZN(_4266_));
 NOR2_X2 _7654_ (.A1(_4335_),
    .A2(_2054_),
    .ZN(_2558_));
 XNOR2_X1 _7655_ (.A(_1953_),
    .B(_2558_),
    .ZN(_4270_));
 XNOR2_X2 _7656_ (.A(_1814_),
    .B(_2026_),
    .ZN(_4291_));
 NOR2_X1 _7657_ (.A1(_4335_),
    .A2(_2058_),
    .ZN(_2559_));
 XNOR2_X1 _7658_ (.A(_1929_),
    .B(_2559_),
    .ZN(_4295_));
 NAND2_X1 _7659_ (.A1(_4307_),
    .A2(_2057_),
    .ZN(_2560_));
 XNOR2_X1 _7660_ (.A(_4475_),
    .B(_2560_),
    .ZN(_4299_));
 INV_X1 _7661_ (.A(_4215_),
    .ZN(_2561_));
 INV_X1 _7662_ (.A(_4221_),
    .ZN(_2562_));
 INV_X1 _7663_ (.A(_4228_),
    .ZN(_2563_));
 INV_X1 _7664_ (.A(_4234_),
    .ZN(_2564_));
 INV_X1 _7665_ (.A(net142),
    .ZN(_2565_));
 OAI211_X2 _7666_ (.A(_1761_),
    .B(_2565_),
    .C1(_1788_),
    .C2(_1789_),
    .ZN(_2566_));
 AOI21_X1 _7667_ (.A(_1966_),
    .B1(net141),
    .B2(_1769_),
    .ZN(_2567_));
 AOI21_X1 _7668_ (.A(_4237_),
    .B1(_2566_),
    .B2(_2567_),
    .ZN(_2568_));
 OAI21_X1 _7669_ (.A(_2564_),
    .B1(_2568_),
    .B2(_2093_),
    .ZN(_2569_));
 AOI21_X1 _7670_ (.A(_4231_),
    .B1(_2569_),
    .B2(_4232_),
    .ZN(_2570_));
 INV_X1 _7671_ (.A(_4229_),
    .ZN(_2571_));
 OAI21_X2 _7672_ (.A(_2563_),
    .B1(_2570_),
    .B2(_2571_),
    .ZN(_2572_));
 AOI21_X1 _7673_ (.A(_4225_),
    .B1(_2572_),
    .B2(_4226_),
    .ZN(_2573_));
 OAI21_X2 _7674_ (.A(_2562_),
    .B1(_2573_),
    .B2(_1961_),
    .ZN(_2574_));
 AOI21_X1 _7675_ (.A(_4218_),
    .B1(_2574_),
    .B2(_4219_),
    .ZN(_2575_));
 OAI21_X2 _7676_ (.A(_2561_),
    .B1(_2575_),
    .B2(_1959_),
    .ZN(_2576_));
 AOI21_X1 _7677_ (.A(_4212_),
    .B1(_2576_),
    .B2(_4213_),
    .ZN(_2577_));
 INV_X1 _7678_ (.A(_2577_),
    .ZN(_2578_));
 AOI21_X2 _7679_ (.A(_4209_),
    .B1(_2578_),
    .B2(_4210_),
    .ZN(_2579_));
 XNOR2_X1 _7680_ (.A(_4207_),
    .B(_2579_),
    .ZN(_4314_));
 AND3_X1 _7681_ (.A1(_1957_),
    .A2(_1958_),
    .A3(_1976_),
    .ZN(_2580_));
 NOR2_X1 _7682_ (.A1(_1977_),
    .A2(_2580_),
    .ZN(_4317_));
 XNOR2_X1 _7683_ (.A(_1969_),
    .B(_2569_),
    .ZN(_4339_));
 INV_X1 _7684_ (.A(_2997_),
    .ZN(_3003_));
 NOR2_X2 _7685_ (.A1(_4279_),
    .A2(_4335_),
    .ZN(_2581_));
 XNOR2_X1 _7686_ (.A(_2581_),
    .B(_4287_),
    .ZN(_4347_));
 CLKBUF_X3 _7687_ (.A(_2108_),
    .Z(_2582_));
 NOR2_X1 _7688_ (.A1(_4305_),
    .A2(_2582_),
    .ZN(_2583_));
 XNOR2_X1 _7689_ (.A(net193),
    .B(_2583_),
    .ZN(_4359_));
 NOR2_X1 _7690_ (.A1(_4335_),
    .A2(_2202_),
    .ZN(_2584_));
 XNOR2_X1 _7691_ (.A(_4355_),
    .B(_2584_),
    .ZN(_4363_));
 NAND2_X2 _7692_ (.A1(_4335_),
    .A2(_2013_),
    .ZN(_2585_));
 OAI21_X1 _7693_ (.A(_2585_),
    .B1(_2075_),
    .B2(net276),
    .ZN(_4371_));
 XNOR2_X1 _7694_ (.A(_4366_),
    .B(_2212_),
    .ZN(_4375_));
 NOR2_X1 _7695_ (.A1(_4335_),
    .A2(_2189_),
    .ZN(_2586_));
 XNOR2_X1 _7696_ (.A(_4372_),
    .B(_2586_),
    .ZN(_4379_));
 XNOR2_X1 _7697_ (.A(_4382_),
    .B(net149),
    .ZN(_4391_));
 XNOR2_X2 _7698_ (.A(_4159_),
    .B(_1940_),
    .ZN(_4395_));
 XNOR2_X1 _7699_ (.A(_4398_),
    .B(_2215_),
    .ZN(_4407_));
 XOR2_X2 _7700_ (.A(_4153_),
    .B(_1916_),
    .Z(_4411_));
 XNOR2_X2 _7701_ (.A(_4414_),
    .B(_2243_),
    .ZN(_4419_));
 INV_X1 _7702_ (.A(_4426_),
    .ZN(_2587_));
 AOI21_X2 _7703_ (.A(_2186_),
    .B1(_2587_),
    .B2(_4307_),
    .ZN(_4427_));
 NAND4_X2 _7704_ (.A1(net111),
    .A2(_4416_),
    .A3(net264),
    .A4(_2230_),
    .ZN(_4431_));
 INV_X1 _7705_ (.A(_4433_),
    .ZN(_2588_));
 AOI21_X2 _7706_ (.A(_2228_),
    .B1(_2588_),
    .B2(_2227_),
    .ZN(_4434_));
 XNOR2_X2 _7707_ (.A(_4441_),
    .B(net223),
    .ZN(_4442_));
 MUX2_X1 _7708_ (.A(_4493_),
    .B(_4454_),
    .S(_2582_),
    .Z(_3010_));
 XOR2_X2 _7709_ (.A(net192),
    .B(net185),
    .Z(_4507_));
 XNOR2_X2 _7710_ (.A(_2064_),
    .B(_2036_),
    .ZN(_4511_));
 AND2_X1 _7711_ (.A1(_4492_),
    .A2(net168),
    .ZN(_2589_));
 AOI21_X1 _7712_ (.A(_2582_),
    .B1(_2271_),
    .B2(_2589_),
    .ZN(_2590_));
 XNOR2_X1 _7713_ (.A(_2279_),
    .B(_2590_),
    .ZN(_4515_));
 NOR4_X4 _7714_ (.A1(net102),
    .A2(_4454_),
    .A3(_4463_),
    .A4(_4471_),
    .ZN(_2591_));
 AOI21_X2 _7715_ (.A(_2108_),
    .B1(net120),
    .B2(_2591_),
    .ZN(_2592_));
 XOR2_X2 _7716_ (.A(net158),
    .B(_2592_),
    .Z(_4519_));
 XNOR2_X2 _7717_ (.A(_2041_),
    .B(net275),
    .ZN(_4527_));
 OR2_X1 _7718_ (.A1(_2227_),
    .A2(_4523_),
    .ZN(_2593_));
 BUF_X4 _7719_ (.A(_2593_),
    .Z(_2594_));
 OAI21_X2 _7720_ (.A(_2594_),
    .B1(_4533_),
    .B2(_2582_),
    .ZN(_4534_));
 XNOR2_X2 _7721_ (.A(_2044_),
    .B(net262),
    .ZN(_4538_));
 NAND3_X2 _7722_ (.A1(_4491_),
    .A2(_4490_),
    .A3(_2258_),
    .ZN(_2595_));
 NOR4_X4 _7723_ (.A1(net156),
    .A2(_4479_),
    .A3(_4471_),
    .A4(_2595_),
    .ZN(_2596_));
 NAND2_X2 _7724_ (.A1(_2227_),
    .A2(_4523_),
    .ZN(_2597_));
 OAI21_X1 _7725_ (.A(_2594_),
    .B1(net273),
    .B2(_2597_),
    .ZN(_4557_));
 INV_X1 _7726_ (.A(net25),
    .ZN(_3015_));
 INV_X1 _7727_ (.A(net32),
    .ZN(_2900_));
 INV_X1 _7728_ (.A(net35),
    .ZN(_3030_));
 INV_X1 _7729_ (.A(net33),
    .ZN(_3038_));
 NAND2_X1 _7730_ (.A1(_2332_),
    .A2(_0191_),
    .ZN(_2598_));
 XNOR2_X1 _7731_ (.A(_3090_),
    .B(_2598_),
    .ZN(_3046_));
 INV_X1 _7732_ (.A(net37),
    .ZN(_3060_));
 INV_X1 _7733_ (.A(net36),
    .ZN(_3068_));
 INV_X1 _7734_ (.A(net38),
    .ZN(_3076_));
 NAND2_X1 _7735_ (.A1(_2942_),
    .A2(_1179_),
    .ZN(_2599_));
 XNOR2_X1 _7736_ (.A(_3230_),
    .B(_2599_),
    .ZN(_3139_));
 MUX2_X1 _7737_ (.A(_3148_),
    .B(_3238_),
    .S(_3261_),
    .Z(_2931_));
 INV_X1 _7738_ (.A(_3014_),
    .ZN(_3152_));
 INV_X1 _7739_ (.A(net39),
    .ZN(_3160_));
 INV_X1 _7740_ (.A(net40),
    .ZN(_3168_));
 INV_X1 _7741_ (.A(net26),
    .ZN(_3184_));
 INV_X1 _7742_ (.A(net41),
    .ZN(_3192_));
 OAI21_X1 _7743_ (.A(_0179_),
    .B1(_2376_),
    .B2(_1052_),
    .ZN(_2600_));
 XNOR2_X1 _7744_ (.A(_3388_),
    .B(_2600_),
    .ZN(_3198_));
 INV_X1 _7745_ (.A(_1178_),
    .ZN(_3234_));
 NOR2_X1 _7746_ (.A1(_3483_),
    .A2(_2427_),
    .ZN(_2601_));
 XNOR2_X1 _7747_ (.A(_0488_),
    .B(_2601_),
    .ZN(_3300_));
 NOR2_X1 _7748_ (.A1(_3312_),
    .A2(_3483_),
    .ZN(_2602_));
 XNOR2_X1 _7749_ (.A(_0476_),
    .B(_2602_),
    .ZN(_3307_));
 MUX2_X1 _7750_ (.A(_3313_),
    .B(_3452_),
    .S(_3483_),
    .Z(_2946_));
 INV_X1 _7751_ (.A(net28),
    .ZN(_3330_));
 INV_X1 _7752_ (.A(net27),
    .ZN(_3338_));
 OAI21_X1 _7753_ (.A(_0179_),
    .B1(_1049_),
    .B2(_1052_),
    .ZN(_2603_));
 XNOR2_X1 _7754_ (.A(_3384_),
    .B(_2603_),
    .ZN(_3344_));
 INV_X1 _7755_ (.A(net30),
    .ZN(_3362_));
 INV_X1 _7756_ (.A(net29),
    .ZN(_3370_));
 AND4_X1 _7757_ (.A1(_1177_),
    .A2(_0774_),
    .A3(_2382_),
    .A4(_2385_),
    .ZN(_2604_));
 NOR2_X1 _7758_ (.A1(net17),
    .A2(_2604_),
    .ZN(_2605_));
 XNOR2_X1 _7759_ (.A(_0763_),
    .B(_2605_),
    .ZN(_3400_));
 XNOR2_X1 _7760_ (.A(_2937_),
    .B(_3244_),
    .ZN(_3460_));
 INV_X1 _7761_ (.A(_2938_),
    .ZN(_2951_));
 NAND2_X1 _7762_ (.A1(_3670_),
    .A2(_1463_),
    .ZN(_2606_));
 XNOR2_X1 _7763_ (.A(_3666_),
    .B(_2606_),
    .ZN(_3518_));
 INV_X1 _7764_ (.A(_3660_),
    .ZN(_3317_));
 NOR2_X1 _7765_ (.A1(_3686_),
    .A2(_1462_),
    .ZN(_2607_));
 XNOR2_X1 _7766_ (.A(_0917_),
    .B(_2607_),
    .ZN(_3525_));
 NOR2_X1 _7767_ (.A1(_3534_),
    .A2(_0901_),
    .ZN(_2608_));
 XNOR2_X1 _7768_ (.A(_0916_),
    .B(_2608_),
    .ZN(_3529_));
 MUX2_X1 _7769_ (.A(_3535_),
    .B(_3644_),
    .S(_3686_),
    .Z(_2955_));
 AOI21_X1 _7770_ (.A(net67),
    .B1(_0763_),
    .B2(_2604_),
    .ZN(_2609_));
 MUX2_X1 _7771_ (.A(net17),
    .B(_2609_),
    .S(_1185_),
    .Z(_3558_));
 XNOR2_X1 _7772_ (.A(_3458_),
    .B(_0857_),
    .ZN(_3652_));
 XOR2_X2 _7773_ (.A(_2952_),
    .B(_0856_),
    .Z(_3656_));
 AOI21_X1 _7774_ (.A(net226),
    .B1(_1680_),
    .B2(_2530_),
    .ZN(_2610_));
 XOR2_X2 _7775_ (.A(_3852_),
    .B(_2610_),
    .Z(_3718_));
 INV_X1 _7776_ (.A(_3814_),
    .ZN(_2611_));
 AOI21_X1 _7777_ (.A(_1321_),
    .B1(_2611_),
    .B2(_2530_),
    .ZN(_2612_));
 XOR2_X2 _7778_ (.A(_3810_),
    .B(_2612_),
    .Z(_3725_));
 NOR2_X1 _7779_ (.A1(_3875_),
    .A2(_1679_),
    .ZN(_2613_));
 XNOR2_X1 _7780_ (.A(_2611_),
    .B(_2613_),
    .ZN(_3729_));
 NOR2_X2 _7781_ (.A1(_3738_),
    .A2(_1321_),
    .ZN(_2614_));
 XOR2_X2 _7782_ (.A(_3818_),
    .B(_2614_),
    .Z(_3733_));
 MUX2_X1 _7783_ (.A(_3739_),
    .B(_3822_),
    .S(_3875_),
    .Z(_2965_));
 XNOR2_X1 _7784_ (.A(_3650_),
    .B(_1289_),
    .ZN(_3830_));
 XNOR2_X1 _7785_ (.A(_1269_),
    .B(_1268_),
    .ZN(_3834_));
 XNOR2_X1 _7786_ (.A(_3658_),
    .B(_2961_),
    .ZN(_3838_));
 INV_X1 _7787_ (.A(_4009_),
    .ZN(_3904_));
 INV_X1 _7788_ (.A(_4010_),
    .ZN(_3743_));
 NOR3_X1 _7789_ (.A1(_3977_),
    .A2(_4027_),
    .A3(_1866_),
    .ZN(_2615_));
 NOR2_X1 _7790_ (.A1(_4053_),
    .A2(_2615_),
    .ZN(_2616_));
 XOR2_X2 _7791_ (.A(_4023_),
    .B(_2616_),
    .Z(_3911_));
 OAI21_X1 _7792_ (.A(_1657_),
    .B1(_2526_),
    .B2(_4027_),
    .ZN(_2617_));
 XNOR2_X1 _7793_ (.A(_3977_),
    .B(_2617_),
    .ZN(_3915_));
 NAND2_X1 _7794_ (.A1(net225),
    .A2(_1866_),
    .ZN(_2618_));
 XNOR2_X1 _7795_ (.A(_4027_),
    .B(_2618_),
    .ZN(_3919_));
 NOR2_X2 _7796_ (.A1(_3928_),
    .A2(_4053_),
    .ZN(_2619_));
 XNOR2_X1 _7797_ (.A(_1865_),
    .B(_2619_),
    .ZN(_3923_));
 MUX2_X1 _7798_ (.A(_3985_),
    .B(_3929_),
    .S(_4031_),
    .Z(_2975_));
 XNOR2_X1 _7799_ (.A(_3828_),
    .B(_1525_),
    .ZN(_3994_));
 XNOR2_X1 _7800_ (.A(_3832_),
    .B(_1543_),
    .ZN(_3998_));
 XNOR2_X1 _7801_ (.A(_2970_),
    .B(_3840_),
    .ZN(_4006_));
 INV_X1 _7802_ (.A(_3860_),
    .ZN(_2620_));
 INV_X1 _7803_ (.A(_3866_),
    .ZN(_2621_));
 INV_X1 _7804_ (.A(_3872_),
    .ZN(_2622_));
 INV_X1 _7805_ (.A(_3879_),
    .ZN(_2623_));
 AOI21_X1 _7806_ (.A(_1577_),
    .B1(_2538_),
    .B2(_2544_),
    .ZN(_2624_));
 OAI21_X1 _7807_ (.A(_3880_),
    .B1(_3882_),
    .B2(_2624_),
    .ZN(_2625_));
 AOI21_X1 _7808_ (.A(_1580_),
    .B1(_2623_),
    .B2(_2625_),
    .ZN(_2626_));
 OAI21_X1 _7809_ (.A(_3873_),
    .B1(_3876_),
    .B2(_2626_),
    .ZN(_2627_));
 AOI21_X1 _7810_ (.A(_1583_),
    .B1(_2622_),
    .B2(_2627_),
    .ZN(_2628_));
 OAI21_X1 _7811_ (.A(_3867_),
    .B1(_3869_),
    .B2(_2628_),
    .ZN(_2629_));
 AOI21_X1 _7812_ (.A(_1586_),
    .B1(_2621_),
    .B2(_2629_),
    .ZN(_2630_));
 OAI21_X1 _7813_ (.A(_3861_),
    .B1(_3863_),
    .B2(_2630_),
    .ZN(_2631_));
 NAND2_X1 _7814_ (.A1(_2620_),
    .A2(_2631_),
    .ZN(_2632_));
 XNOR2_X2 _7815_ (.A(_1589_),
    .B(_2632_),
    .ZN(_4032_));
 XOR2_X2 _7816_ (.A(_3861_),
    .B(_1587_),
    .Z(_4035_));
 NAND2_X1 _7817_ (.A1(_2621_),
    .A2(_2629_),
    .ZN(_2633_));
 XNOR2_X2 _7818_ (.A(_1586_),
    .B(_2633_),
    .ZN(_4038_));
 XOR2_X2 _7819_ (.A(_3867_),
    .B(_1584_),
    .Z(_4041_));
 NAND2_X1 _7820_ (.A1(_2622_),
    .A2(_2627_),
    .ZN(_2634_));
 XNOR2_X1 _7821_ (.A(_1583_),
    .B(_2634_),
    .ZN(_4044_));
 XOR2_X2 _7822_ (.A(_3873_),
    .B(_1581_),
    .Z(_4047_));
 NAND2_X1 _7823_ (.A1(_2623_),
    .A2(_2625_),
    .ZN(_2635_));
 XNOR2_X1 _7824_ (.A(_1580_),
    .B(_2635_),
    .ZN(_4050_));
 XOR2_X2 _7825_ (.A(_3880_),
    .B(_1578_),
    .Z(_4054_));
 XOR2_X2 _7826_ (.A(_3886_),
    .B(_1575_),
    .Z(_4060_));
 NAND2_X1 _7827_ (.A1(_2539_),
    .A2(_2542_),
    .ZN(_2636_));
 XNOR2_X1 _7828_ (.A(_1574_),
    .B(_2636_),
    .ZN(_4063_));
 XOR2_X2 _7829_ (.A(_3892_),
    .B(_1572_),
    .Z(_4066_));
 XNOR2_X1 _7830_ (.A(_3895_),
    .B(_2540_),
    .ZN(_4069_));
 INV_X1 _7831_ (.A(_3974_),
    .ZN(_2637_));
 NOR2_X2 _7832_ (.A1(_1870_),
    .A2(_2526_),
    .ZN(_2638_));
 NOR2_X1 _7833_ (.A1(net220),
    .A2(_2638_),
    .ZN(_2639_));
 XNOR2_X1 _7834_ (.A(_2639_),
    .B(_2637_),
    .ZN(_4076_));
 NAND2_X1 _7835_ (.A1(net3),
    .A2(_2553_),
    .ZN(_2640_));
 XNOR2_X1 _7836_ (.A(_4179_),
    .B(_2640_),
    .ZN(_4084_));
 XNOR2_X1 _7837_ (.A(_1799_),
    .B(_1612_),
    .ZN(_4088_));
 XNOR2_X1 _7838_ (.A(_1611_),
    .B(_1797_),
    .ZN(_4092_));
 XNOR2_X1 _7839_ (.A(_1796_),
    .B(_1609_),
    .ZN(_4096_));
 XOR2_X2 _7840_ (.A(_3925_),
    .B(_2976_),
    .Z(_4100_));
 NAND2_X2 _7841_ (.A1(_1873_),
    .A2(_1872_),
    .ZN(_2641_));
 AOI21_X1 _7842_ (.A(net220),
    .B1(_2637_),
    .B2(_2638_),
    .ZN(_2642_));
 NAND2_X1 _7843_ (.A1(_2641_),
    .A2(_2642_),
    .ZN(_2643_));
 NAND2_X1 _7844_ (.A1(_1883_),
    .A2(_2643_),
    .ZN(_4113_));
 NAND2_X1 _7845_ (.A1(_1883_),
    .A2(_2643_),
    .ZN(_4121_));
 XNOR2_X2 _7846_ (.A(_2641_),
    .B(_1884_),
    .ZN(_4125_));
 NAND2_X1 _7847_ (.A1(_1883_),
    .A2(_1885_),
    .ZN(_4129_));
 NAND2_X1 _7848_ (.A1(_1883_),
    .A2(_2643_),
    .ZN(_4117_));
 NAND2_X1 _7849_ (.A1(_1883_),
    .A2(_1885_),
    .ZN(_4135_));
 XOR2_X2 _7850_ (.A(_4000_),
    .B(_1730_),
    .Z(_4161_));
 INV_X1 _7851_ (.A(_4048_),
    .ZN(_2644_));
 INV_X1 _7852_ (.A(_4055_),
    .ZN(_2645_));
 INV_X1 _7853_ (.A(_4061_),
    .ZN(_2646_));
 INV_X1 _7854_ (.A(_4067_),
    .ZN(_2647_));
 NAND2_X1 _7855_ (.A1(_1769_),
    .A2(_1569_),
    .ZN(_2648_));
 INV_X1 _7856_ (.A(_1569_),
    .ZN(_2649_));
 OAI211_X2 _7857_ (.A(_1562_),
    .B(_2649_),
    .C1(_1588_),
    .C2(_1589_),
    .ZN(_2650_));
 AOI21_X1 _7858_ (.A(_1771_),
    .B1(_2648_),
    .B2(_2650_),
    .ZN(_2651_));
 OAI21_X1 _7859_ (.A(_4068_),
    .B1(_4070_),
    .B2(_2651_),
    .ZN(_2652_));
 AOI21_X1 _7860_ (.A(_1774_),
    .B1(_2647_),
    .B2(_2652_),
    .ZN(_2653_));
 OAI21_X1 _7861_ (.A(_4062_),
    .B1(_4064_),
    .B2(_2653_),
    .ZN(_2654_));
 AOI21_X1 _7862_ (.A(_1777_),
    .B1(_2646_),
    .B2(_2654_),
    .ZN(_2655_));
 OAI21_X1 _7863_ (.A(_4056_),
    .B1(_4058_),
    .B2(_2655_),
    .ZN(_2656_));
 AOI21_X1 _7864_ (.A(_1780_),
    .B1(_2645_),
    .B2(_2656_),
    .ZN(_2657_));
 OAI21_X1 _7865_ (.A(_4049_),
    .B1(_4051_),
    .B2(_2657_),
    .ZN(_2658_));
 NAND2_X1 _7866_ (.A1(_2644_),
    .A2(_2658_),
    .ZN(_2659_));
 AND2_X1 _7867_ (.A1(_4043_),
    .A2(_4046_),
    .ZN(_2660_));
 AOI221_X2 _7868_ (.A(_4042_),
    .B1(_2659_),
    .B2(_2660_),
    .C1(_4045_),
    .C2(_4043_),
    .ZN(_2661_));
 OAI21_X1 _7869_ (.A(_1762_),
    .B1(_2661_),
    .B2(_1786_),
    .ZN(_2662_));
 AOI21_X1 _7870_ (.A(_4036_),
    .B1(_2662_),
    .B2(_4037_),
    .ZN(_2663_));
 XNOR2_X1 _7871_ (.A(_4034_),
    .B(_2663_),
    .ZN(_4199_));
 XOR2_X2 _7872_ (.A(_4037_),
    .B(_1787_),
    .Z(_4202_));
 XNOR2_X1 _7873_ (.A(_4040_),
    .B(_2661_),
    .ZN(_4205_));
 XOR2_X2 _7874_ (.A(_4043_),
    .B(_1784_),
    .Z(_4208_));
 XNOR2_X1 _7875_ (.A(_1783_),
    .B(_2659_),
    .ZN(_4211_));
 XOR2_X2 _7876_ (.A(_4049_),
    .B(_1781_),
    .Z(_4214_));
 AND3_X1 _7877_ (.A1(_1780_),
    .A2(_2645_),
    .A3(_2656_),
    .ZN(_2664_));
 NOR2_X1 _7878_ (.A1(_2657_),
    .A2(_2664_),
    .ZN(_4217_));
 XOR2_X2 _7879_ (.A(_4056_),
    .B(_1778_),
    .Z(_4220_));
 AND3_X1 _7880_ (.A1(_1777_),
    .A2(_2646_),
    .A3(_2654_),
    .ZN(_2665_));
 NOR2_X1 _7881_ (.A1(_2655_),
    .A2(_2665_),
    .ZN(_4224_));
 XOR2_X2 _7882_ (.A(_4062_),
    .B(_1775_),
    .Z(_4227_));
 NAND2_X1 _7883_ (.A1(_2647_),
    .A2(_2652_),
    .ZN(_2666_));
 XNOR2_X1 _7884_ (.A(_1774_),
    .B(_2666_),
    .ZN(_4230_));
 XOR2_X2 _7885_ (.A(net234),
    .B(_1772_),
    .Z(_4233_));
 NAND2_X1 _7886_ (.A1(_2648_),
    .A2(_2650_),
    .ZN(_2667_));
 XNOR2_X1 _7887_ (.A(_1771_),
    .B(_2667_),
    .ZN(_4236_));
 XOR2_X2 _7888_ (.A(_1769_),
    .B(net141),
    .Z(_4239_));
 NAND2_X1 _7889_ (.A1(_2176_),
    .A2(_2177_),
    .ZN(_4243_));
 OAI21_X1 _7890_ (.A(_2585_),
    .B1(_2075_),
    .B2(net276),
    .ZN(_4252_));
 OAI21_X1 _7891_ (.A(_2585_),
    .B1(_2075_),
    .B2(_2013_),
    .ZN(_4255_));
 XNOR2_X1 _7892_ (.A(_2022_),
    .B(_1809_),
    .ZN(_4263_));
 NAND2_X1 _7893_ (.A1(_4307_),
    .A2(_2055_),
    .ZN(_2668_));
 XNOR2_X1 _7894_ (.A(_4459_),
    .B(_2668_),
    .ZN(_4267_));
 XOR2_X2 _7895_ (.A(_2986_),
    .B(net116),
    .Z(_4271_));
 NAND2_X1 _7896_ (.A1(_4438_),
    .A2(_4307_),
    .ZN(_2669_));
 XNOR2_X2 _7897_ (.A(_2053_),
    .B(_2669_),
    .ZN(_3006_));
 NAND2_X1 _7898_ (.A1(_2552_),
    .A2(_2555_),
    .ZN(_2670_));
 NAND2_X1 _7899_ (.A1(_2177_),
    .A2(_2670_),
    .ZN(_4284_));
 OAI21_X1 _7900_ (.A(_2585_),
    .B1(_2075_),
    .B2(_2013_),
    .ZN(_4288_));
 OAI21_X2 _7901_ (.A(_2585_),
    .B1(_4261_),
    .B2(_4335_),
    .ZN(_4292_));
 XNOR2_X1 _7902_ (.A(_2025_),
    .B(_1812_),
    .ZN(_4296_));
 XNOR2_X2 _7903_ (.A(_1811_),
    .B(_2023_),
    .ZN(_4300_));
 INV_X1 _7904_ (.A(_4207_),
    .ZN(_2671_));
 OAI21_X1 _7905_ (.A(_1956_),
    .B1(_2579_),
    .B2(_2671_),
    .ZN(_2672_));
 AOI21_X1 _7906_ (.A(_4203_),
    .B1(_2672_),
    .B2(_4204_),
    .ZN(_2673_));
 XNOR2_X1 _7907_ (.A(_4201_),
    .B(_2673_),
    .ZN(_4308_));
 AND3_X1 _7908_ (.A1(_1955_),
    .A2(_1956_),
    .A3(_1978_),
    .ZN(_2674_));
 NOR2_X1 _7909_ (.A1(_1979_),
    .A2(_2674_),
    .ZN(_4311_));
 XOR2_X2 _7910_ (.A(_4213_),
    .B(_2576_),
    .Z(_4320_));
 AND3_X1 _7911_ (.A1(_1959_),
    .A2(_1960_),
    .A3(_1974_),
    .ZN(_2675_));
 NOR2_X1 _7912_ (.A1(_1975_),
    .A2(_2675_),
    .ZN(_4323_));
 XOR2_X2 _7913_ (.A(_4219_),
    .B(_2574_),
    .Z(_4326_));
 AND3_X1 _7914_ (.A1(_1961_),
    .A2(_1962_),
    .A3(_1972_),
    .ZN(_2676_));
 NOR2_X1 _7915_ (.A1(_1973_),
    .A2(_2676_),
    .ZN(_4329_));
 XOR2_X2 _7916_ (.A(_4226_),
    .B(_2572_),
    .Z(_4332_));
 XNOR2_X1 _7917_ (.A(_2571_),
    .B(_1970_),
    .ZN(_4336_));
 INV_X2 _7918_ (.A(net303),
    .ZN(_3004_));
 XOR2_X2 _7919_ (.A(_2990_),
    .B(net91),
    .Z(_4348_));
 NAND2_X1 _7920_ (.A1(_2176_),
    .A2(_2177_),
    .ZN(_4352_));
 OAI21_X1 _7921_ (.A(_2585_),
    .B1(_2075_),
    .B2(_2013_),
    .ZN(_4356_));
 XNOR2_X1 _7922_ (.A(_2996_),
    .B(net97),
    .ZN(_4360_));
 XNOR2_X2 _7923_ (.A(net278),
    .B(_1938_),
    .ZN(_4364_));
 NAND2_X1 _7924_ (.A1(_2177_),
    .A2(_2670_),
    .ZN(_4368_));
 NOR2_X2 _7925_ (.A1(_2582_),
    .A2(_2229_),
    .ZN(_2677_));
 XNOR2_X2 _7926_ (.A(_2677_),
    .B(net190),
    .ZN(_4376_));
 XOR2_X2 _7927_ (.A(_4163_),
    .B(_1913_),
    .Z(_4380_));
 NAND2_X1 _7928_ (.A1(_2176_),
    .A2(_2177_),
    .ZN(_4384_));
 OAI21_X1 _7929_ (.A(_2585_),
    .B1(_2075_),
    .B2(net276),
    .ZN(_4388_));
 AOI21_X1 _7930_ (.A(_2582_),
    .B1(_2252_),
    .B2(net119),
    .ZN(_2678_));
 XNOR2_X1 _7931_ (.A(_4558_),
    .B(_2678_),
    .ZN(_4392_));
 NAND2_X1 _7932_ (.A1(_4307_),
    .A2(_2203_),
    .ZN(_2679_));
 XOR2_X2 _7933_ (.A(_4387_),
    .B(_2679_),
    .Z(_4396_));
 NAND2_X1 _7934_ (.A1(_2177_),
    .A2(_2670_),
    .ZN(_4400_));
 OAI21_X1 _7935_ (.A(_2585_),
    .B1(_2075_),
    .B2(net276),
    .ZN(_4404_));
 AOI21_X1 _7936_ (.A(_2108_),
    .B1(net263),
    .B2(_2230_),
    .ZN(_2680_));
 XNOR2_X1 _7937_ (.A(_4561_),
    .B(_2680_),
    .ZN(_4408_));
 XNOR2_X1 _7938_ (.A(_2187_),
    .B(_2191_),
    .ZN(_4412_));
 INV_X1 _7939_ (.A(_4418_),
    .ZN(_2681_));
 AOI21_X2 _7940_ (.A(_2228_),
    .B1(_2227_),
    .B2(_2681_),
    .ZN(_4420_));
 XNOR2_X2 _7941_ (.A(_1918_),
    .B(_1941_),
    .ZN(_4428_));
 XNOR2_X2 _7942_ (.A(net94),
    .B(_2218_),
    .ZN(_4435_));
 AOI21_X1 _7943_ (.A(_2228_),
    .B1(_2232_),
    .B2(_4415_),
    .ZN(_4443_));
 NOR2_X1 _7944_ (.A1(_4492_),
    .A2(_2582_),
    .ZN(_2682_));
 XNOR2_X1 _7945_ (.A(net106),
    .B(_2682_),
    .ZN(_4508_));
 NAND2_X1 _7946_ (.A1(_2227_),
    .A2(_2595_),
    .ZN(_2683_));
 XNOR2_X1 _7947_ (.A(_4471_),
    .B(_2683_),
    .ZN(_4512_));
 XNOR2_X2 _7948_ (.A(_2038_),
    .B(_2065_),
    .ZN(_4516_));
 XNOR2_X2 _7949_ (.A(_2067_),
    .B(net237),
    .ZN(_4520_));
 NAND2_X2 _7950_ (.A1(_4492_),
    .A2(net217),
    .ZN(_2684_));
 NOR4_X4 _7951_ (.A1(_4479_),
    .A2(_4487_),
    .A3(_4471_),
    .A4(_2684_),
    .ZN(_2685_));
 INV_X1 _7952_ (.A(_2685_),
    .ZN(_4524_));
 OAI21_X2 _7953_ (.A(_2594_),
    .B1(_4526_),
    .B2(_2582_),
    .ZN(_4528_));
 NAND2_X1 _7954_ (.A1(_4523_),
    .A2(_2596_),
    .ZN(_4531_));
 XNOR2_X2 _7955_ (.A(net236),
    .B(net189),
    .ZN(_4535_));
 OAI21_X2 _7956_ (.A(_2594_),
    .B1(_2597_),
    .B2(net122),
    .ZN(_4539_));
 OAI21_X1 _7957_ (.A(_2594_),
    .B1(net271),
    .B2(_2597_),
    .ZN(_4543_));
 OAI21_X1 _7958_ (.A(_2594_),
    .B1(_2597_),
    .B2(net123),
    .ZN(_4547_));
 OAI21_X1 _7959_ (.A(_2594_),
    .B1(net272),
    .B2(_2597_),
    .ZN(_4551_));
 INV_X1 _7960_ (.A(_4525_),
    .ZN(_2686_));
 OAI21_X1 _7961_ (.A(_2594_),
    .B1(_2582_),
    .B2(_2686_),
    .ZN(_4562_));
 INV_X1 _7962_ (.A(net315),
    .ZN(net75));
 INV_X1 _7963_ (.A(_4544_),
    .ZN(_2687_));
 INV_X1 _7964_ (.A(_4536_),
    .ZN(_2688_));
 INV_X1 _7965_ (.A(_4521_),
    .ZN(_2689_));
 INV_X1 _7966_ (.A(_4513_),
    .ZN(_2690_));
 AOI21_X1 _7967_ (.A(_4509_),
    .B1(_3011_),
    .B2(_4510_),
    .ZN(_2691_));
 INV_X1 _7968_ (.A(_4514_),
    .ZN(_2692_));
 OAI21_X2 _7969_ (.A(_2690_),
    .B1(_2691_),
    .B2(_2692_),
    .ZN(_2693_));
 AOI21_X1 _7970_ (.A(_4517_),
    .B1(_2693_),
    .B2(_4518_),
    .ZN(_2694_));
 INV_X1 _7971_ (.A(_4522_),
    .ZN(_2695_));
 OAI21_X2 _7972_ (.A(_2689_),
    .B1(_2694_),
    .B2(_2695_),
    .ZN(_2696_));
 AOI21_X2 _7973_ (.A(_4529_),
    .B1(_4530_),
    .B2(_2696_),
    .ZN(_2697_));
 INV_X1 _7974_ (.A(_4537_),
    .ZN(_2698_));
 OAI21_X2 _7975_ (.A(_2688_),
    .B1(_2698_),
    .B2(_2697_),
    .ZN(_2699_));
 AOI21_X2 _7976_ (.A(_4540_),
    .B1(_2699_),
    .B2(_4541_),
    .ZN(_2700_));
 INV_X1 _7977_ (.A(_4545_),
    .ZN(_2701_));
 OAI21_X2 _7978_ (.A(_2687_),
    .B1(_2700_),
    .B2(_2701_),
    .ZN(_2702_));
 XNOR2_X2 _7979_ (.A(net129),
    .B(_4549_),
    .ZN(_2703_));
 CLKBUF_X3 _7980_ (.A(_4504_),
    .Z(_2704_));
 INV_X1 _7981_ (.A(_2704_),
    .ZN(_2705_));
 INV_X1 _7982_ (.A(_4540_),
    .ZN(_2706_));
 INV_X1 _7983_ (.A(_4529_),
    .ZN(_2707_));
 INV_X1 _7984_ (.A(_4517_),
    .ZN(_2708_));
 INV_X1 _7985_ (.A(_4509_),
    .ZN(_2709_));
 AOI21_X1 _7986_ (.A(_4494_),
    .B1(_4495_),
    .B2(_3009_),
    .ZN(_2710_));
 INV_X1 _7987_ (.A(_4510_),
    .ZN(_2711_));
 OAI21_X2 _7988_ (.A(_2709_),
    .B1(_2710_),
    .B2(_2711_),
    .ZN(_2712_));
 AOI21_X1 _7989_ (.A(_4513_),
    .B1(_2712_),
    .B2(net110),
    .ZN(_2713_));
 INV_X1 _7990_ (.A(_4518_),
    .ZN(_2714_));
 OAI21_X2 _7991_ (.A(_2708_),
    .B1(_2713_),
    .B2(_2714_),
    .ZN(_2715_));
 AOI21_X2 _7992_ (.A(_4521_),
    .B1(_2715_),
    .B2(net104),
    .ZN(_2716_));
 INV_X2 _7993_ (.A(_4530_),
    .ZN(_2717_));
 OAI21_X4 _7994_ (.A(_2707_),
    .B1(_2717_),
    .B2(_2716_),
    .ZN(_2718_));
 AOI21_X4 _7995_ (.A(_4536_),
    .B1(_2718_),
    .B2(net99),
    .ZN(_2719_));
 INV_X1 _7996_ (.A(_4541_),
    .ZN(_2720_));
 OAI21_X4 _7997_ (.A(_2706_),
    .B1(_2720_),
    .B2(_2719_),
    .ZN(_2721_));
 XNOR2_X2 _7998_ (.A(net162),
    .B(_4545_),
    .ZN(_2722_));
 XNOR2_X2 _7999_ (.A(net128),
    .B(_4541_),
    .ZN(_2723_));
 XNOR2_X2 _8000_ (.A(net100),
    .B(net173),
    .ZN(_2724_));
 XNOR2_X2 _8001_ (.A(net92),
    .B(_2696_),
    .ZN(_2725_));
 XNOR2_X2 _8002_ (.A(_2715_),
    .B(net105),
    .ZN(_2726_));
 INV_X1 _8003_ (.A(_2726_),
    .ZN(_2727_));
 XNOR2_X2 _8004_ (.A(_4518_),
    .B(_2693_),
    .ZN(_2728_));
 XNOR2_X2 _8005_ (.A(_4514_),
    .B(_2712_),
    .ZN(_2729_));
 NAND2_X2 _8006_ (.A1(_2728_),
    .A2(_2729_),
    .ZN(_2730_));
 XNOR2_X2 _8007_ (.A(net161),
    .B(net284),
    .ZN(_2731_));
 NAND2_X2 _8008_ (.A1(_4499_),
    .A2(_2731_),
    .ZN(_2732_));
 NOR3_X4 _8009_ (.A1(_2727_),
    .A2(_2730_),
    .A3(_2732_),
    .ZN(_2733_));
 NAND3_X2 _8010_ (.A1(_2724_),
    .A2(_2725_),
    .A3(_2733_),
    .ZN(_2734_));
 INV_X1 _8011_ (.A(_2734_),
    .ZN(_2735_));
 AND3_X4 _8012_ (.A1(_2735_),
    .A2(_2723_),
    .A3(_2722_),
    .ZN(_2736_));
 NOR2_X1 _8013_ (.A1(_2705_),
    .A2(_2736_),
    .ZN(_2737_));
 XNOR2_X1 _8014_ (.A(net180),
    .B(_2737_),
    .ZN(net57));
 INV_X1 _8015_ (.A(_4548_),
    .ZN(_2738_));
 AOI21_X4 _8016_ (.A(_4544_),
    .B1(_4545_),
    .B2(_2721_),
    .ZN(_2739_));
 INV_X1 _8017_ (.A(_4549_),
    .ZN(_2740_));
 OAI21_X4 _8018_ (.A(_2738_),
    .B1(_2740_),
    .B2(_2739_),
    .ZN(_2741_));
 XNOR2_X2 _8019_ (.A(_4553_),
    .B(net143),
    .ZN(_2742_));
 NAND3_X2 _8020_ (.A1(_4498_),
    .A2(_4497_),
    .A3(_2731_),
    .ZN(_2743_));
 NOR2_X4 _8021_ (.A1(_2730_),
    .A2(_2743_),
    .ZN(_2744_));
 NAND3_X4 _8022_ (.A1(_2725_),
    .A2(_2726_),
    .A3(_2744_),
    .ZN(_2745_));
 NAND2_X2 _8023_ (.A1(_2724_),
    .A2(_2723_),
    .ZN(_2746_));
 NOR2_X4 _8024_ (.A1(_2746_),
    .A2(_2745_),
    .ZN(_2747_));
 NAND3_X4 _8025_ (.A1(_2747_),
    .A2(_2722_),
    .A3(_2703_),
    .ZN(_2748_));
 NAND2_X2 _8026_ (.A1(_2704_),
    .A2(_2748_),
    .ZN(_2749_));
 XOR2_X1 _8027_ (.A(_2742_),
    .B(_2749_),
    .Z(net58));
 INV_X1 _8028_ (.A(_4552_),
    .ZN(_2750_));
 AOI21_X1 _8029_ (.A(_4548_),
    .B1(_2702_),
    .B2(_4549_),
    .ZN(_2751_));
 INV_X1 _8030_ (.A(_4553_),
    .ZN(_2752_));
 OAI21_X2 _8031_ (.A(_2750_),
    .B1(_2751_),
    .B2(_2752_),
    .ZN(_2753_));
 XNOR2_X2 _8032_ (.A(_2753_),
    .B(_4556_),
    .ZN(_2754_));
 NAND3_X1 _8033_ (.A1(net180),
    .A2(_2736_),
    .A3(_2742_),
    .ZN(_2755_));
 NAND2_X1 _8034_ (.A1(_2704_),
    .A2(_2755_),
    .ZN(_2756_));
 XOR2_X1 _8035_ (.A(_2756_),
    .B(_2754_),
    .Z(net59));
 INV_X1 _8036_ (.A(_4555_),
    .ZN(_2757_));
 AOI21_X1 _8037_ (.A(_4552_),
    .B1(_2741_),
    .B2(_4553_),
    .ZN(_2758_));
 INV_X1 _8038_ (.A(_4556_),
    .ZN(_2759_));
 OAI21_X2 _8039_ (.A(_2757_),
    .B1(_2758_),
    .B2(_2759_),
    .ZN(_2760_));
 XOR2_X2 _8040_ (.A(_4560_),
    .B(_2760_),
    .Z(_2761_));
 NAND2_X2 _8041_ (.A1(_2742_),
    .A2(_2754_),
    .ZN(_2762_));
 OAI21_X4 _8042_ (.A(_4504_),
    .B1(_2748_),
    .B2(_2762_),
    .ZN(_2763_));
 XNOR2_X1 _8043_ (.A(_2761_),
    .B(_2763_),
    .ZN(net60));
 AOI21_X1 _8044_ (.A(_4555_),
    .B1(_2753_),
    .B2(_4556_),
    .ZN(_2764_));
 INV_X1 _8045_ (.A(_2764_),
    .ZN(_2765_));
 AOI21_X1 _8046_ (.A(_4559_),
    .B1(_2765_),
    .B2(_4560_),
    .ZN(_2766_));
 XNOR2_X1 _8047_ (.A(_4564_),
    .B(_2766_),
    .ZN(_2767_));
 NAND4_X2 _8048_ (.A1(_2703_),
    .A2(_2736_),
    .A3(net172),
    .A4(_2754_),
    .ZN(_2768_));
 OAI21_X2 _8049_ (.A(_2704_),
    .B1(_2768_),
    .B2(_2761_),
    .ZN(_2769_));
 XNOR2_X1 _8050_ (.A(_2767_),
    .B(_2769_),
    .ZN(net61));
 OAI21_X1 _8051_ (.A(_4504_),
    .B1(_2761_),
    .B2(_2767_),
    .ZN(_2770_));
 NAND2_X1 _8052_ (.A1(_2763_),
    .A2(_2770_),
    .ZN(_2771_));
 AOI21_X1 _8053_ (.A(_4559_),
    .B1(net159),
    .B2(_4560_),
    .ZN(_2772_));
 INV_X1 _8054_ (.A(_2772_),
    .ZN(_2773_));
 AOI21_X1 _8055_ (.A(_4563_),
    .B1(_2773_),
    .B2(_4564_),
    .ZN(_2774_));
 XOR2_X1 _8056_ (.A(_2771_),
    .B(_2774_),
    .Z(_2775_));
 XNOR2_X1 _8057_ (.A(net114),
    .B(_2775_),
    .ZN(_2776_));
 NOR2_X1 _8058_ (.A1(_4532_),
    .A2(_2108_),
    .ZN(_2777_));
 AOI21_X1 _8059_ (.A(_2777_),
    .B1(_4523_),
    .B2(_2582_),
    .ZN(_2778_));
 XNOR2_X1 _8060_ (.A(_2776_),
    .B(_2778_),
    .ZN(net62));
 MUX2_X1 _8061_ (.A(_3012_),
    .B(_4500_),
    .S(_2704_),
    .Z(net63));
 NOR2_X2 _8062_ (.A1(net297),
    .A2(_2705_),
    .ZN(_2779_));
 XNOR2_X1 _8063_ (.A(_2731_),
    .B(_2779_),
    .ZN(net64));
 NAND2_X1 _8064_ (.A1(_2704_),
    .A2(_2743_),
    .ZN(_2780_));
 XOR2_X1 _8065_ (.A(_2729_),
    .B(_2780_),
    .Z(net65));
 INV_X1 _8066_ (.A(_2729_),
    .ZN(_2781_));
 OAI21_X2 _8067_ (.A(_2704_),
    .B1(_2781_),
    .B2(_2732_),
    .ZN(_2782_));
 XOR2_X1 _8068_ (.A(_2728_),
    .B(_2782_),
    .Z(net66));
 NOR2_X1 _8069_ (.A1(_2705_),
    .A2(_2744_),
    .ZN(_2783_));
 XNOR2_X1 _8070_ (.A(_2783_),
    .B(_2726_),
    .ZN(net70));
 NOR2_X1 _8071_ (.A1(_2705_),
    .A2(_2733_),
    .ZN(_2784_));
 XNOR2_X1 _8072_ (.A(_2725_),
    .B(_2784_),
    .ZN(net71));
 NAND2_X1 _8073_ (.A1(_2704_),
    .A2(_2745_),
    .ZN(_2785_));
 XOR2_X1 _8074_ (.A(_2724_),
    .B(_2785_),
    .Z(net72));
 NAND2_X1 _8075_ (.A1(_2704_),
    .A2(_2734_),
    .ZN(_2786_));
 XOR2_X1 _8076_ (.A(_2723_),
    .B(_2786_),
    .Z(net73));
 OAI21_X2 _8077_ (.A(_2704_),
    .B1(_2746_),
    .B2(_2745_),
    .ZN(_2787_));
 XOR2_X1 _8078_ (.A(_2787_),
    .B(_2722_),
    .Z(net74));
 INV_X1 _8079_ (.A(_4444_),
    .ZN(_2788_));
 INV_X1 _8080_ (.A(_4421_),
    .ZN(_2789_));
 INV_X1 _8081_ (.A(_4393_),
    .ZN(_2790_));
 INV_X1 _8082_ (.A(_4361_),
    .ZN(_2791_));
 INV_X1 _8083_ (.A(_4362_),
    .ZN(_2792_));
 OAI21_X4 _8084_ (.A(_2791_),
    .B1(_2792_),
    .B2(_3001_),
    .ZN(_2793_));
 AOI21_X4 _8085_ (.A(_4377_),
    .B1(net289),
    .B2(_2793_),
    .ZN(_2794_));
 INV_X1 _8086_ (.A(_4394_),
    .ZN(_2795_));
 OAI21_X4 _8087_ (.A(_2790_),
    .B1(_2794_),
    .B2(_2795_),
    .ZN(_2796_));
 AOI21_X2 _8088_ (.A(_4409_),
    .B1(_2796_),
    .B2(_4410_),
    .ZN(_2797_));
 INV_X1 _8089_ (.A(_4422_),
    .ZN(_2798_));
 OAI21_X4 _8090_ (.A(_2789_),
    .B1(_2798_),
    .B2(_2797_),
    .ZN(_2799_));
 AOI21_X4 _8091_ (.A(_4436_),
    .B1(_2799_),
    .B2(_4437_),
    .ZN(_2800_));
 INV_X1 _8092_ (.A(_4445_),
    .ZN(_2801_));
 OAI21_X4 _8093_ (.A(_2788_),
    .B1(_2800_),
    .B2(_2801_),
    .ZN(_2802_));
 AOI21_X4 _8094_ (.A(_4448_),
    .B1(_4449_),
    .B2(_2802_),
    .ZN(_2803_));
 XNOR2_X2 _8095_ (.A(_2803_),
    .B(_4457_),
    .ZN(_2804_));
 NOR2_X4 _8096_ (.A1(_4502_),
    .A2(_4503_),
    .ZN(_2805_));
 INV_X1 _8097_ (.A(_4436_),
    .ZN(_2806_));
 INV_X1 _8098_ (.A(_4409_),
    .ZN(_2807_));
 INV_X1 _8099_ (.A(_4377_),
    .ZN(_2808_));
 INV_X1 _8100_ (.A(_4342_),
    .ZN(_2809_));
 INV_X1 _8101_ (.A(_4343_),
    .ZN(_2810_));
 OAI21_X4 _8102_ (.A(_2809_),
    .B1(_2810_),
    .B2(_2999_),
    .ZN(_2811_));
 AOI21_X4 _8103_ (.A(_4361_),
    .B1(_2811_),
    .B2(net115),
    .ZN(_2812_));
 INV_X2 _8104_ (.A(net289),
    .ZN(_2813_));
 OAI21_X2 _8105_ (.A(_2808_),
    .B1(_2812_),
    .B2(_2813_),
    .ZN(_2814_));
 AOI21_X2 _8106_ (.A(_4393_),
    .B1(net108),
    .B2(_2814_),
    .ZN(_2815_));
 INV_X2 _8107_ (.A(_4410_),
    .ZN(_2816_));
 OAI21_X2 _8108_ (.A(_2807_),
    .B1(_2815_),
    .B2(_2816_),
    .ZN(_2817_));
 AOI21_X4 _8109_ (.A(_4421_),
    .B1(_2817_),
    .B2(net95),
    .ZN(_2818_));
 INV_X1 _8110_ (.A(_4437_),
    .ZN(_2819_));
 OAI21_X4 _8111_ (.A(_2806_),
    .B1(_2818_),
    .B2(_2819_),
    .ZN(_2820_));
 AOI21_X4 _8112_ (.A(_4444_),
    .B1(_2820_),
    .B2(_4445_),
    .ZN(_2821_));
 XNOR2_X2 _8113_ (.A(_4449_),
    .B(_2821_),
    .ZN(_2822_));
 INV_X1 _8114_ (.A(_2822_),
    .ZN(_2823_));
 XNOR2_X2 _8115_ (.A(_2801_),
    .B(net137),
    .ZN(_2824_));
 XNOR2_X2 _8116_ (.A(_2818_),
    .B(net246),
    .ZN(_2825_));
 XNOR2_X2 _8117_ (.A(net248),
    .B(net153),
    .ZN(_2826_));
 XNOR2_X2 _8118_ (.A(net231),
    .B(_2816_),
    .ZN(_2827_));
 INV_X2 _8119_ (.A(_2827_),
    .ZN(_2828_));
 XNOR2_X2 _8120_ (.A(_2794_),
    .B(net107),
    .ZN(_2829_));
 XNOR2_X2 _8121_ (.A(net261),
    .B(net184),
    .ZN(_2830_));
 XOR2_X2 _8122_ (.A(_3001_),
    .B(net109),
    .Z(_2831_));
 NAND2_X1 _8123_ (.A1(_4345_),
    .A2(_2831_),
    .ZN(_2832_));
 OR4_X4 _8124_ (.A1(_2828_),
    .A2(_2829_),
    .A3(net290),
    .A4(_2832_),
    .ZN(_2833_));
 NOR3_X4 _8125_ (.A1(net287),
    .A2(_2833_),
    .A3(_2825_),
    .ZN(_2834_));
 NAND3_X4 _8126_ (.A1(_2823_),
    .A2(net202),
    .A3(_2834_),
    .ZN(_2835_));
 NAND2_X2 _8127_ (.A1(_2805_),
    .A2(_2835_),
    .ZN(_2836_));
 XNOR2_X1 _8128_ (.A(_2804_),
    .B(_2836_),
    .ZN(net76));
 INV_X1 _8129_ (.A(_4448_),
    .ZN(_2837_));
 INV_X1 _8130_ (.A(_4449_),
    .ZN(_2838_));
 OAI21_X2 _8131_ (.A(_2837_),
    .B1(_2821_),
    .B2(_2838_),
    .ZN(_2839_));
 AOI21_X2 _8132_ (.A(_4456_),
    .B1(_2839_),
    .B2(_4457_),
    .ZN(_2840_));
 XNOR2_X2 _8133_ (.A(_2840_),
    .B(_4465_),
    .ZN(_2841_));
 NAND2_X2 _8134_ (.A1(_0000_),
    .A2(_0002_),
    .ZN(_2842_));
 INV_X1 _8135_ (.A(_2825_),
    .ZN(_2843_));
 NAND3_X1 _8136_ (.A1(_3002_),
    .A2(_4344_),
    .A3(_2831_),
    .ZN(_2844_));
 OR3_X4 _8137_ (.A1(_2829_),
    .A2(_2830_),
    .A3(_2844_),
    .ZN(_2845_));
 NOR3_X4 _8138_ (.A1(_2826_),
    .A2(_2828_),
    .A3(_2845_),
    .ZN(_2846_));
 NAND3_X2 _8139_ (.A1(_2843_),
    .A2(_2824_),
    .A3(_2846_),
    .ZN(_2847_));
 NOR3_X4 _8140_ (.A1(_2847_),
    .A2(_2822_),
    .A3(_2804_),
    .ZN(_2848_));
 NOR2_X1 _8141_ (.A1(_2842_),
    .A2(_2848_),
    .ZN(_2849_));
 XOR2_X1 _8142_ (.A(_2841_),
    .B(_2849_),
    .Z(net77));
 INV_X1 _8143_ (.A(_4456_),
    .ZN(_2850_));
 INV_X1 _8144_ (.A(_4457_),
    .ZN(_2851_));
 OAI21_X4 _8145_ (.A(_2850_),
    .B1(_2851_),
    .B2(_2803_),
    .ZN(_2852_));
 AOI21_X4 _8146_ (.A(_4464_),
    .B1(_4465_),
    .B2(_2852_),
    .ZN(_2853_));
 XNOR2_X2 _8147_ (.A(_2853_),
    .B(_4473_),
    .ZN(_2854_));
 INV_X2 _8148_ (.A(_2854_),
    .ZN(_2855_));
 NOR3_X4 _8149_ (.A1(_2835_),
    .A2(_2804_),
    .A3(_2841_),
    .ZN(_2856_));
 NOR2_X2 _8150_ (.A1(_2842_),
    .A2(_2856_),
    .ZN(_2857_));
 XNOR2_X1 _8151_ (.A(_2855_),
    .B(_2857_),
    .ZN(net78));
 INV_X1 _8152_ (.A(_4464_),
    .ZN(_2858_));
 INV_X1 _8153_ (.A(_4465_),
    .ZN(_2859_));
 OAI21_X2 _8154_ (.A(_2858_),
    .B1(_2840_),
    .B2(_2859_),
    .ZN(_2860_));
 AOI21_X2 _8155_ (.A(_4472_),
    .B1(_2860_),
    .B2(_4473_),
    .ZN(_2861_));
 XNOR2_X2 _8156_ (.A(_4481_),
    .B(_2861_),
    .ZN(_2862_));
 NAND2_X4 _8157_ (.A1(_2848_),
    .A2(_2855_),
    .ZN(_2863_));
 OAI21_X4 _8158_ (.A(_2805_),
    .B1(_2841_),
    .B2(_2863_),
    .ZN(_2864_));
 XNOR2_X1 _8159_ (.A(_2862_),
    .B(_2864_),
    .ZN(net79));
 INV_X1 _8160_ (.A(_4472_),
    .ZN(_2865_));
 INV_X1 _8161_ (.A(_4473_),
    .ZN(_2866_));
 OAI21_X1 _8162_ (.A(_2865_),
    .B1(_2853_),
    .B2(_2866_),
    .ZN(_2867_));
 AOI21_X2 _8163_ (.A(_4480_),
    .B1(_2867_),
    .B2(_4481_),
    .ZN(_2868_));
 XNOR2_X1 _8164_ (.A(_4489_),
    .B(_2868_),
    .ZN(_2869_));
 NAND2_X2 _8165_ (.A1(_2855_),
    .A2(_2856_),
    .ZN(_2870_));
 OAI21_X2 _8166_ (.A(_2805_),
    .B1(_2862_),
    .B2(_2870_),
    .ZN(_2871_));
 XNOR2_X1 _8167_ (.A(_2869_),
    .B(_2871_),
    .ZN(net80));
 INV_X1 _8168_ (.A(_4480_),
    .ZN(_2872_));
 INV_X1 _8169_ (.A(_4481_),
    .ZN(_2873_));
 OAI21_X1 _8170_ (.A(_2872_),
    .B1(_2861_),
    .B2(_2873_),
    .ZN(_2874_));
 AOI21_X1 _8171_ (.A(_4488_),
    .B1(_2874_),
    .B2(_4489_),
    .ZN(_2875_));
 OAI21_X1 _8172_ (.A(_2805_),
    .B1(_2862_),
    .B2(_2869_),
    .ZN(_2876_));
 NAND2_X1 _8173_ (.A1(_2876_),
    .A2(_2864_),
    .ZN(_2877_));
 XOR2_X1 _8174_ (.A(_2877_),
    .B(_2875_),
    .Z(_2878_));
 AND2_X1 _8175_ (.A1(_4432_),
    .A2(_2227_),
    .ZN(_2879_));
 NOR4_X2 _8176_ (.A1(_4405_),
    .A2(_2227_),
    .A3(_2194_),
    .A4(_2200_),
    .ZN(_2880_));
 AND4_X1 _8177_ (.A1(_2158_),
    .A2(_2108_),
    .A3(_2194_),
    .A4(_2200_),
    .ZN(_2881_));
 NOR3_X1 _8178_ (.A1(_2158_),
    .A2(_4405_),
    .A3(_2226_),
    .ZN(_2882_));
 AND2_X1 _8179_ (.A1(_4405_),
    .A2(_2108_),
    .ZN(_2883_));
 MUX2_X1 _8180_ (.A(_2882_),
    .B(_2883_),
    .S(_2194_),
    .Z(_2884_));
 NOR4_X2 _8181_ (.A1(_2879_),
    .A2(_2880_),
    .A3(_2881_),
    .A4(_2884_),
    .ZN(_2885_));
 XNOR2_X1 _8182_ (.A(_2885_),
    .B(_2878_),
    .ZN(_2886_));
 XNOR2_X1 _8183_ (.A(_4523_),
    .B(_2886_),
    .ZN(net81));
 NOR2_X1 _8184_ (.A1(_4346_),
    .A2(_2842_),
    .ZN(_2887_));
 AOI21_X1 _8185_ (.A(_2887_),
    .B1(_2842_),
    .B2(_3002_),
    .ZN(net82));
 NOR2_X1 _8186_ (.A1(_4345_),
    .A2(_2842_),
    .ZN(_2888_));
 XNOR2_X1 _8187_ (.A(_2831_),
    .B(_2888_),
    .ZN(net83));
 NAND2_X1 _8188_ (.A1(_2805_),
    .A2(_2844_),
    .ZN(_2889_));
 XNOR2_X1 _8189_ (.A(_2830_),
    .B(_2889_),
    .ZN(net84));
 OAI21_X2 _8190_ (.A(_2805_),
    .B1(net290),
    .B2(_2832_),
    .ZN(_2890_));
 XNOR2_X1 _8191_ (.A(_2829_),
    .B(_2890_),
    .ZN(net85));
 NAND2_X2 _8192_ (.A1(_2845_),
    .A2(_2805_),
    .ZN(_2891_));
 XOR2_X1 _8193_ (.A(_2891_),
    .B(_2827_),
    .Z(net86));
 NAND2_X4 _8194_ (.A1(_2805_),
    .A2(_2833_),
    .ZN(_2892_));
 XNOR2_X1 _8195_ (.A(net288),
    .B(_2892_),
    .ZN(net87));
 NOR2_X1 _8196_ (.A1(_2842_),
    .A2(_2846_),
    .ZN(_2893_));
 XNOR2_X1 _8197_ (.A(_2843_),
    .B(_2893_),
    .ZN(net88));
 NOR2_X2 _8198_ (.A1(_2842_),
    .A2(_2834_),
    .ZN(_2894_));
 XNOR2_X1 _8199_ (.A(net203),
    .B(_2894_),
    .ZN(net89));
 NAND2_X2 _8200_ (.A1(_2847_),
    .A2(_2805_),
    .ZN(_2895_));
 XNOR2_X1 _8201_ (.A(_2822_),
    .B(_2895_),
    .ZN(net90));
 FA_X1 _8202_ (.A(_2896_),
    .B(net32),
    .CI(_2897_),
    .CO(_2898_),
    .S(_2899_));
 FA_X1 _8203_ (.A(_2896_),
    .B(_2900_),
    .CI(_2901_),
    .CO(_2902_),
    .S(_2903_));
 FA_X1 _8204_ (.A(net14),
    .B(_2900_),
    .CI(_2904_),
    .CO(_2905_),
    .S(_2906_));
 FA_X1 _8205_ (.A(_2908_),
    .B(_2907_),
    .CI(_2909_),
    .CO(_2910_),
    .S(_2911_));
 FA_X1 _8206_ (.A(_2912_),
    .B(_2913_),
    .CI(_2914_),
    .CO(_2915_),
    .S(_2916_));
 FA_X1 _8207_ (.A(_2917_),
    .B(_2918_),
    .CI(_2919_),
    .CO(_2920_),
    .S(_2921_));
 FA_X1 _8208_ (.A(_2924_),
    .B(_2925_),
    .CI(_2910_),
    .CO(_2926_),
    .S(_2927_));
 FA_X1 _8209_ (.A(_2930_),
    .B(_2916_),
    .CI(_2931_),
    .CO(_2932_),
    .S(_2933_));
 FA_X1 _8210_ (.A(_2934_),
    .B(_2935_),
    .CI(_2936_),
    .CO(_2937_),
    .S(_2938_));
 FA_X1 _8211_ (.A(_2940_),
    .B(_2941_),
    .CI(_2942_),
    .CO(_2943_),
    .S(_2944_));
 FA_X1 _8212_ (.A(_2945_),
    .B(_2933_),
    .CI(_2946_),
    .CO(_2947_),
    .S(_2948_));
 FA_X1 _8213_ (.A(_2949_),
    .B(_2950_),
    .CI(_2951_),
    .CO(_2952_),
    .S(_2953_));
 FA_X1 _8214_ (.A(_2954_),
    .B(_2948_),
    .CI(_2955_),
    .CO(_2956_),
    .S(_2957_));
 FA_X1 _8215_ (.A(_2958_),
    .B(_2959_),
    .CI(_2960_),
    .CO(_2961_),
    .S(_2962_));
 FA_X1 _8216_ (.A(_2964_),
    .B(_2957_),
    .CI(_2965_),
    .CO(_2966_),
    .S(_2967_));
 FA_X1 _8217_ (.A(_2962_),
    .B(_2968_),
    .CI(_2969_),
    .CO(_2970_),
    .S(_2971_));
 FA_X1 _8218_ (.A(_2974_),
    .B(_2967_),
    .CI(_2975_),
    .CO(_2976_),
    .S(_2977_));
 FA_X1 _8219_ (.A(_2978_),
    .B(_2980_),
    .CI(net139),
    .CO(_2981_),
    .S(_2982_));
 FA_X1 _8220_ (.A(_2984_),
    .B(_2985_),
    .CI(_2977_),
    .CO(_2986_),
    .S(_2987_));
 FA_X1 _8221_ (.A(_2982_),
    .B(_2988_),
    .CI(_2989_),
    .CO(_2990_),
    .S(_2991_));
 FA_X1 _8222_ (.A(_2993_),
    .B(_2994_),
    .CI(_2995_),
    .CO(_2996_),
    .S(_2997_));
 FA_X1 _8223_ (.A(_2997_),
    .B(_2999_),
    .CI(_3000_),
    .CO(_3001_),
    .S(_3002_));
 FA_X1 _8224_ (.A(_2987_),
    .B(_3005_),
    .CI(_3006_),
    .CO(_3007_),
    .S(_3008_));
 FA_X1 _8225_ (.A(_3010_),
    .B(_3009_),
    .CI(_3008_),
    .CO(_3011_),
    .S(_3012_));
 HA_X1 _8226_ (.A(_3013_),
    .B(net25),
    .CO(_2897_),
    .S(_3014_));
 HA_X1 _8227_ (.A(net5),
    .B(_3015_),
    .CO(_2904_),
    .S(_3016_));
 HA_X1 _8228_ (.A(net5),
    .B(net25),
    .CO(_3017_),
    .S(_3018_));
 HA_X1 _8229_ (.A(_2896_),
    .B(net32),
    .CO(_3020_),
    .S(_3019_));
 HA_X1 _8230_ (.A(net14),
    .B(_2900_),
    .CO(_3021_),
    .S(_3022_));
 HA_X1 _8231_ (.A(net14),
    .B(net32),
    .CO(_3023_),
    .S(_3024_));
 HA_X1 _8232_ (.A(_3025_),
    .B(_3014_),
    .CO(_2922_),
    .S(_3026_));
 HA_X1 _8233_ (.A(_3027_),
    .B(net35),
    .CO(_3028_),
    .S(_3029_));
 HA_X1 _8234_ (.A(net16),
    .B(_3030_),
    .CO(_3031_),
    .S(_3032_));
 HA_X1 _8235_ (.A(net16),
    .B(net35),
    .CO(_3033_),
    .S(_3034_));
 HA_X1 _8236_ (.A(net33),
    .B(_3035_),
    .CO(_3036_),
    .S(_3037_));
 HA_X1 _8237_ (.A(net15),
    .B(_3038_),
    .CO(_3039_),
    .S(_3040_));
 HA_X1 _8238_ (.A(net15),
    .B(net33),
    .CO(_3041_),
    .S(_3042_));
 HA_X1 _8239_ (.A(_2908_),
    .B(_2909_),
    .CO(_3043_),
    .S(_3044_));
 HA_X1 _8240_ (.A(_3045_),
    .B(_3046_),
    .CO(_3047_),
    .S(_3048_));
 HA_X1 _8241_ (.A(_2923_),
    .B(_3049_),
    .CO(_3050_),
    .S(_3051_));
 HA_X1 _8242_ (.A(_3052_),
    .B(_3025_),
    .CO(_3053_),
    .S(_3054_));
 HA_X1 _8243_ (.A(_3055_),
    .B(_3026_),
    .CO(_2934_),
    .S(_3056_));
 HA_X1 _8244_ (.A(net37),
    .B(_3057_),
    .CO(_3058_),
    .S(_3059_));
 HA_X1 _8245_ (.A(net20),
    .B(_3060_),
    .CO(_3061_),
    .S(_3062_));
 HA_X1 _8246_ (.A(net20),
    .B(net37),
    .CO(_3063_),
    .S(_3064_));
 HA_X1 _8247_ (.A(_3065_),
    .B(net36),
    .CO(_3066_),
    .S(_3067_));
 HA_X1 _8248_ (.A(net19),
    .B(_3068_),
    .CO(_3069_),
    .S(_3070_));
 HA_X1 _8249_ (.A(net19),
    .B(net36),
    .CO(_3071_),
    .S(_3072_));
 HA_X1 _8250_ (.A(_3073_),
    .B(net38),
    .CO(_3074_),
    .S(_3075_));
 HA_X1 _8251_ (.A(net21),
    .B(_3076_),
    .CO(_3077_),
    .S(_3078_));
 HA_X1 _8252_ (.A(net21),
    .B(net38),
    .CO(_3079_),
    .S(_3080_));
 HA_X1 _8253_ (.A(_3081_),
    .B(_3082_),
    .CO(_3083_),
    .S(_3084_));
 HA_X1 _8254_ (.A(_3085_),
    .B(_3086_),
    .CO(_3087_),
    .S(_3088_));
 HA_X1 _8255_ (.A(_3089_),
    .B(_3090_),
    .CO(_3091_),
    .S(_3092_));
 HA_X1 _8256_ (.A(_3093_),
    .B(_3094_),
    .CO(_3095_),
    .S(_3096_));
 HA_X1 _8257_ (.A(_3097_),
    .B(_2914_),
    .CO(_3098_),
    .S(_3099_));
 HA_X1 _8258_ (.A(_2919_),
    .B(_2918_),
    .CO(_3100_),
    .S(_3101_));
 HA_X1 _8259_ (.A(_2910_),
    .B(_3102_),
    .CO(_3103_),
    .S(_3104_));
 HA_X1 _8260_ (.A(_3105_),
    .B(_2929_),
    .CO(_3106_),
    .S(_3107_));
 HA_X1 _8261_ (.A(_3108_),
    .B(_2910_),
    .CO(_3109_),
    .S(_3110_));
 HA_X1 _8262_ (.A(_3111_),
    .B(_2910_),
    .CO(_3112_),
    .S(_3113_));
 HA_X1 _8263_ (.A(_3114_),
    .B(_2929_),
    .CO(_3115_),
    .S(_3116_));
 HA_X1 _8264_ (.A(_3117_),
    .B(_2910_),
    .CO(_3118_),
    .S(_3119_));
 HA_X1 _8265_ (.A(_3120_),
    .B(_2929_),
    .CO(_3121_),
    .S(_3122_));
 HA_X1 _8266_ (.A(_3123_),
    .B(_2929_),
    .CO(_3124_),
    .S(_3125_));
 HA_X1 _8267_ (.A(_3126_),
    .B(_2929_),
    .CO(_3127_),
    .S(_3128_));
 HA_X1 _8268_ (.A(_3129_),
    .B(_2910_),
    .CO(_3130_),
    .S(_3131_));
 HA_X1 _8269_ (.A(_2925_),
    .B(_2910_),
    .CO(_3132_),
    .S(_3133_));
 HA_X1 _8270_ (.A(_3134_),
    .B(_3135_),
    .CO(_3136_),
    .S(_3137_));
 HA_X1 _8271_ (.A(_3138_),
    .B(_3139_),
    .CO(_3140_),
    .S(_3141_));
 HA_X1 _8272_ (.A(_3142_),
    .B(_3055_),
    .CO(_3143_),
    .S(_3144_));
 HA_X1 _8273_ (.A(_3145_),
    .B(_3146_),
    .CO(_3147_),
    .S(_3148_));
 HA_X1 _8274_ (.A(_2916_),
    .B(_2931_),
    .CO(_3150_),
    .S(_3151_));
 HA_X1 _8275_ (.A(_2919_),
    .B(_3152_),
    .CO(_3149_),
    .S(_3153_));
 HA_X1 _8276_ (.A(_3154_),
    .B(_3056_),
    .CO(_3155_),
    .S(_3156_));
 HA_X1 _8277_ (.A(_3157_),
    .B(net39),
    .CO(_3158_),
    .S(_3159_));
 HA_X1 _8278_ (.A(net22),
    .B(_3160_),
    .CO(_3161_),
    .S(_3162_));
 HA_X1 _8279_ (.A(net22),
    .B(net39),
    .CO(_3163_),
    .S(_3164_));
 HA_X1 _8280_ (.A(_3165_),
    .B(net40),
    .CO(_3166_),
    .S(_3167_));
 HA_X1 _8281_ (.A(net23),
    .B(_3168_),
    .CO(_3169_),
    .S(_3170_));
 HA_X1 _8282_ (.A(net23),
    .B(net40),
    .CO(_3171_),
    .S(_3172_));
 HA_X1 _8283_ (.A(_3173_),
    .B(_3174_),
    .CO(_3175_),
    .S(_3176_));
 HA_X1 _8284_ (.A(_3177_),
    .B(_3178_),
    .CO(_3179_),
    .S(_3180_));
 HA_X1 _8285_ (.A(_3181_),
    .B(net26),
    .CO(_3182_),
    .S(_3183_));
 HA_X1 _8286_ (.A(net6),
    .B(_3184_),
    .CO(_3185_),
    .S(_3186_));
 HA_X1 _8287_ (.A(net6),
    .B(net26),
    .CO(_3187_),
    .S(_3188_));
 HA_X1 _8288_ (.A(_3189_),
    .B(net41),
    .CO(_3190_),
    .S(_3191_));
 HA_X1 _8289_ (.A(net24),
    .B(_3192_),
    .CO(_3193_),
    .S(_3194_));
 HA_X1 _8290_ (.A(net24),
    .B(net41),
    .CO(_3195_),
    .S(_3196_));
 HA_X1 _8291_ (.A(_3197_),
    .B(_3198_),
    .CO(_3199_),
    .S(_3200_));
 HA_X1 _8292_ (.A(_3201_),
    .B(_3202_),
    .CO(_3203_),
    .S(_3204_));
 HA_X1 _8293_ (.A(_3205_),
    .B(_3206_),
    .CO(_3207_),
    .S(_3208_));
 HA_X1 _8294_ (.A(_3209_),
    .B(_3210_),
    .CO(_3211_),
    .S(_3212_));
 HA_X1 _8295_ (.A(_3213_),
    .B(_3214_),
    .CO(_3215_),
    .S(_3216_));
 HA_X1 _8296_ (.A(_3217_),
    .B(_3218_),
    .CO(_3219_),
    .S(_3220_));
 HA_X1 _8297_ (.A(_3221_),
    .B(_3222_),
    .CO(_3223_),
    .S(_3224_));
 HA_X1 _8298_ (.A(_3225_),
    .B(_3226_),
    .CO(_3227_),
    .S(_3228_));
 HA_X1 _8299_ (.A(_3229_),
    .B(_3230_),
    .CO(_3231_),
    .S(_3232_));
 HA_X1 _8300_ (.A(_3233_),
    .B(_3234_),
    .CO(_3235_),
    .S(_3236_));
 HA_X1 _8301_ (.A(_3237_),
    .B(_3238_),
    .CO(_3239_),
    .S(_3240_));
 HA_X1 _8302_ (.A(_3241_),
    .B(_3242_),
    .CO(_3243_),
    .S(_3244_));
 HA_X1 _8303_ (.A(_3245_),
    .B(_3246_),
    .CO(_3247_),
    .S(_3248_));
 HA_X1 _8304_ (.A(_2939_),
    .B(_2921_),
    .CO(_3249_),
    .S(_3250_));
 HA_X1 _8305_ (.A(_2942_),
    .B(_3251_),
    .CO(_3252_),
    .S(_3253_));
 HA_X1 _8306_ (.A(_3254_),
    .B(_2942_),
    .CO(_3255_),
    .S(_3256_));
 HA_X1 _8307_ (.A(_3257_),
    .B(_2942_),
    .CO(_3258_),
    .S(_3259_));
 HA_X1 _8308_ (.A(_3260_),
    .B(_3261_),
    .CO(_3262_),
    .S(_3263_));
 HA_X1 _8309_ (.A(_3264_),
    .B(_2942_),
    .CO(_3265_),
    .S(_3266_));
 HA_X1 _8310_ (.A(_3267_),
    .B(_2942_),
    .CO(_3268_),
    .S(_3269_));
 HA_X1 _8311_ (.A(_3270_),
    .B(net17),
    .CO(_3271_),
    .S(_3272_));
 HA_X1 _8312_ (.A(_3273_),
    .B(net17),
    .CO(_3274_),
    .S(_3275_));
 HA_X1 _8313_ (.A(_3276_),
    .B(_3261_),
    .CO(_3277_),
    .S(_3278_));
 HA_X1 _8314_ (.A(_3279_),
    .B(_3261_),
    .CO(_3280_),
    .S(_3281_));
 HA_X1 _8315_ (.A(_3282_),
    .B(_3261_),
    .CO(_3283_),
    .S(_3284_));
 HA_X1 _8316_ (.A(_2927_),
    .B(_3261_),
    .CO(_3285_),
    .S(_3286_));
 HA_X1 _8317_ (.A(_2928_),
    .B(_2942_),
    .CO(_3287_),
    .S(_3288_));
 HA_X1 _8318_ (.A(_2940_),
    .B(_3289_),
    .CO(_3290_),
    .S(_3291_));
 HA_X1 _8319_ (.A(_3261_),
    .B(_3292_),
    .CO(_3293_),
    .S(_3294_));
 HA_X1 _8320_ (.A(_3295_),
    .B(_3296_),
    .CO(_3297_),
    .S(_3298_));
 HA_X1 _8321_ (.A(_3299_),
    .B(_3300_),
    .CO(_3301_),
    .S(_3302_));
 HA_X1 _8322_ (.A(_3303_),
    .B(_3154_),
    .CO(_3304_),
    .S(_3305_));
 HA_X1 _8323_ (.A(_3306_),
    .B(_3307_),
    .CO(_3308_),
    .S(_3309_));
 HA_X1 _8324_ (.A(_3310_),
    .B(_3311_),
    .CO(_3312_),
    .S(_3313_));
 HA_X1 _8325_ (.A(_2933_),
    .B(_2946_),
    .CO(_3314_),
    .S(_3315_));
 HA_X1 _8326_ (.A(_3153_),
    .B(_3242_),
    .CO(_2930_),
    .S(_3316_));
 HA_X1 _8327_ (.A(_3317_),
    .B(_3156_),
    .CO(_2958_),
    .S(_3318_));
 HA_X1 _8328_ (.A(_3319_),
    .B(_3320_),
    .CO(_3321_),
    .S(_3322_));
 HA_X1 _8329_ (.A(_3323_),
    .B(_3324_),
    .CO(_3325_),
    .S(_3326_));
 HA_X1 _8330_ (.A(_3327_),
    .B(net28),
    .CO(_3328_),
    .S(_3329_));
 HA_X1 _8331_ (.A(net8),
    .B(_3330_),
    .CO(_3331_),
    .S(_3332_));
 HA_X1 _8332_ (.A(net8),
    .B(net28),
    .CO(_3333_),
    .S(_3334_));
 HA_X1 _8333_ (.A(_3335_),
    .B(net27),
    .CO(_3336_),
    .S(_3337_));
 HA_X1 _8334_ (.A(net7),
    .B(_3338_),
    .CO(_3339_),
    .S(_3340_));
 HA_X1 _8335_ (.A(net7),
    .B(net27),
    .CO(_3341_),
    .S(_3342_));
 HA_X1 _8336_ (.A(_3343_),
    .B(_3344_),
    .CO(_3345_),
    .S(_3346_));
 HA_X1 _8337_ (.A(_3347_),
    .B(_3348_),
    .CO(_3349_),
    .S(_3350_));
 HA_X1 _8338_ (.A(_3351_),
    .B(_3352_),
    .CO(_3353_),
    .S(_3354_));
 HA_X1 _8339_ (.A(_3356_),
    .B(_3355_),
    .CO(_3357_),
    .S(_3358_));
 HA_X1 _8340_ (.A(_3359_),
    .B(net30),
    .CO(_3360_),
    .S(_3361_));
 HA_X1 _8341_ (.A(net12),
    .B(_3362_),
    .CO(_3363_),
    .S(_3364_));
 HA_X1 _8342_ (.A(net12),
    .B(net30),
    .CO(_3365_),
    .S(_3366_));
 HA_X1 _8343_ (.A(_3367_),
    .B(net29),
    .CO(_3368_),
    .S(_3369_));
 HA_X1 _8344_ (.A(net11),
    .B(_3370_),
    .CO(_3371_),
    .S(_3372_));
 HA_X1 _8345_ (.A(net11),
    .B(net29),
    .CO(_3373_),
    .S(_3374_));
 HA_X1 _8346_ (.A(_3375_),
    .B(_3376_),
    .CO(_3377_),
    .S(_3378_));
 HA_X1 _8347_ (.A(_3379_),
    .B(_3380_),
    .CO(_3381_),
    .S(_3382_));
 HA_X1 _8348_ (.A(_3383_),
    .B(_3384_),
    .CO(_3385_),
    .S(_3386_));
 HA_X1 _8349_ (.A(_3387_),
    .B(_3388_),
    .CO(_3389_),
    .S(_3390_));
 HA_X1 _8350_ (.A(_3391_),
    .B(_3392_),
    .CO(_3393_),
    .S(_3394_));
 HA_X1 _8351_ (.A(_3395_),
    .B(_3396_),
    .CO(_3397_),
    .S(_3398_));
 HA_X1 _8352_ (.A(_3399_),
    .B(_3400_),
    .CO(_3401_),
    .S(_3402_));
 HA_X1 _8353_ (.A(_3403_),
    .B(_3404_),
    .CO(_3405_),
    .S(_3406_));
 HA_X1 _8354_ (.A(_3407_),
    .B(_3408_),
    .CO(_3409_),
    .S(_3410_));
 HA_X1 _8355_ (.A(_3411_),
    .B(_3412_),
    .CO(_3413_),
    .S(_3414_));
 HA_X1 _8356_ (.A(_3415_),
    .B(_3416_),
    .CO(_3417_),
    .S(_3418_));
 HA_X1 _8357_ (.A(_3419_),
    .B(_3420_),
    .CO(_3421_),
    .S(_3422_));
 HA_X1 _8358_ (.A(_3423_),
    .B(_3424_),
    .CO(_3425_),
    .S(_3426_));
 HA_X1 _8359_ (.A(_3427_),
    .B(_3428_),
    .CO(_3429_),
    .S(_3430_));
 HA_X1 _8360_ (.A(_3431_),
    .B(_3432_),
    .CO(_3433_),
    .S(_3434_));
 HA_X1 _8361_ (.A(_3435_),
    .B(_3436_),
    .CO(_3437_),
    .S(_3438_));
 HA_X1 _8362_ (.A(_3439_),
    .B(_3440_),
    .CO(_3441_),
    .S(_3442_));
 HA_X1 _8363_ (.A(_3443_),
    .B(_3444_),
    .CO(_3445_),
    .S(_3446_));
 HA_X1 _8364_ (.A(_3447_),
    .B(_3448_),
    .CO(_3449_),
    .S(_3450_));
 HA_X1 _8365_ (.A(_3451_),
    .B(_3452_),
    .CO(_3453_),
    .S(_3454_));
 HA_X1 _8366_ (.A(_3455_),
    .B(_3456_),
    .CO(_3457_),
    .S(_3458_));
 HA_X1 _8367_ (.A(_3459_),
    .B(_3460_),
    .CO(_3461_),
    .S(_3462_));
 HA_X1 _8368_ (.A(_3463_),
    .B(_3464_),
    .CO(_3465_),
    .S(_3466_));
 HA_X1 _8369_ (.A(_2950_),
    .B(_2951_),
    .CO(_3467_),
    .S(_3468_));
 HA_X1 _8370_ (.A(_3469_),
    .B(net218),
    .CO(_3471_),
    .S(_3472_));
 HA_X1 _8371_ (.A(_3473_),
    .B(net218),
    .CO(_3474_),
    .S(_3475_));
 HA_X1 _8372_ (.A(_3476_),
    .B(net9),
    .CO(_3477_),
    .S(_3478_));
 HA_X1 _8373_ (.A(_3479_),
    .B(net9),
    .CO(_3480_),
    .S(_3481_));
 HA_X1 _8374_ (.A(_3482_),
    .B(_3483_),
    .CO(_3484_),
    .S(_3485_));
 HA_X1 _8375_ (.A(_3486_),
    .B(net218),
    .CO(_3487_),
    .S(_3488_));
 HA_X1 _8376_ (.A(_3489_),
    .B(_3483_),
    .CO(_3490_),
    .S(_3491_));
 HA_X1 _8377_ (.A(_3492_),
    .B(_3470_),
    .CO(_3493_),
    .S(_3494_));
 HA_X1 _8378_ (.A(_3495_),
    .B(net218),
    .CO(_3496_),
    .S(_3497_));
 HA_X1 _8379_ (.A(_3498_),
    .B(_3470_),
    .CO(_3499_),
    .S(_3500_));
 HA_X1 _8380_ (.A(_3501_),
    .B(_3483_),
    .CO(_3502_),
    .S(_3503_));
 HA_X1 _8381_ (.A(_3504_),
    .B(_3470_),
    .CO(_3505_),
    .S(_3506_));
 HA_X1 _8382_ (.A(_3507_),
    .B(_3470_),
    .CO(_3508_),
    .S(_3509_));
 HA_X1 _8383_ (.A(_3510_),
    .B(_3470_),
    .CO(_3511_),
    .S(_3512_));
 HA_X1 _8384_ (.A(_3513_),
    .B(_3514_),
    .CO(_3515_),
    .S(_3516_));
 HA_X1 _8385_ (.A(_3517_),
    .B(_3518_),
    .CO(_3519_),
    .S(_3520_));
 HA_X1 _8386_ (.A(_3521_),
    .B(_3317_),
    .CO(_3522_),
    .S(_3523_));
 HA_X1 _8387_ (.A(_3524_),
    .B(_3525_),
    .CO(_3526_),
    .S(_3527_));
 HA_X1 _8388_ (.A(_3528_),
    .B(_3529_),
    .CO(_3530_),
    .S(_3531_));
 HA_X1 _8389_ (.A(_3532_),
    .B(_3533_),
    .CO(_3534_),
    .S(_3535_));
 HA_X1 _8390_ (.A(_2948_),
    .B(_2955_),
    .CO(_3536_),
    .S(_3537_));
 HA_X1 _8391_ (.A(_3316_),
    .B(_3456_),
    .CO(_2945_),
    .S(_3538_));
 HA_X1 _8392_ (.A(_3539_),
    .B(_3318_),
    .CO(_2968_),
    .S(_3540_));
 HA_X1 _8393_ (.A(_3542_),
    .B(_3541_),
    .CO(_3543_),
    .S(_3544_));
 HA_X1 _8394_ (.A(_3545_),
    .B(_3546_),
    .CO(_3547_),
    .S(_3548_));
 HA_X1 _8395_ (.A(_3549_),
    .B(_3550_),
    .CO(_3551_),
    .S(_3552_));
 HA_X1 _8396_ (.A(_3553_),
    .B(_3554_),
    .CO(_3555_),
    .S(_3556_));
 HA_X1 _8397_ (.A(_3557_),
    .B(_3558_),
    .CO(_3559_),
    .S(_3560_));
 HA_X1 _8398_ (.A(_3561_),
    .B(_3562_),
    .CO(_3563_),
    .S(_3564_));
 HA_X1 _8399_ (.A(_3565_),
    .B(_3566_),
    .CO(_3567_),
    .S(_3568_));
 HA_X1 _8400_ (.A(_3569_),
    .B(_3570_),
    .CO(_3571_),
    .S(_3572_));
 HA_X1 _8401_ (.A(_3574_),
    .B(_3573_),
    .CO(_3575_),
    .S(_3576_));
 HA_X1 _8402_ (.A(_3577_),
    .B(_3578_),
    .CO(_3579_),
    .S(_3580_));
 HA_X1 _8403_ (.A(_3582_),
    .B(_3581_),
    .CO(_3583_),
    .S(_3584_));
 HA_X1 _8404_ (.A(_3585_),
    .B(_3586_),
    .CO(_3587_),
    .S(_3588_));
 HA_X1 _8405_ (.A(_3589_),
    .B(_3590_),
    .CO(_3591_),
    .S(_3592_));
 HA_X1 _8406_ (.A(_3590_),
    .B(_3589_),
    .CO(_3593_),
    .S(_3594_));
 HA_X1 _8407_ (.A(_3595_),
    .B(_3596_),
    .CO(_3597_),
    .S(_3598_));
 HA_X1 _8408_ (.A(_3599_),
    .B(_3600_),
    .CO(_3601_),
    .S(_3602_));
 HA_X1 _8409_ (.A(_3603_),
    .B(_3604_),
    .CO(_3605_),
    .S(_3606_));
 HA_X1 _8410_ (.A(_3607_),
    .B(_3608_),
    .CO(_3609_),
    .S(_3610_));
 HA_X1 _8411_ (.A(_3611_),
    .B(_3612_),
    .CO(_3613_),
    .S(_3614_));
 HA_X1 _8412_ (.A(_3615_),
    .B(_3616_),
    .CO(_3617_),
    .S(_3618_));
 HA_X1 _8413_ (.A(_3619_),
    .B(_3620_),
    .CO(_3621_),
    .S(_3622_));
 HA_X1 _8414_ (.A(_3623_),
    .B(_3624_),
    .CO(_3625_),
    .S(_3626_));
 HA_X1 _8415_ (.A(_3627_),
    .B(_3628_),
    .CO(_3629_),
    .S(_3630_));
 HA_X1 _8416_ (.A(_3631_),
    .B(_3632_),
    .CO(_3633_),
    .S(_3634_));
 HA_X1 _8417_ (.A(_3635_),
    .B(_3636_),
    .CO(_3637_),
    .S(_3638_));
 HA_X1 _8418_ (.A(_3639_),
    .B(_3640_),
    .CO(_3641_),
    .S(_3642_));
 HA_X1 _8419_ (.A(_3643_),
    .B(_3644_),
    .CO(_3645_),
    .S(_3646_));
 HA_X1 _8420_ (.A(_3647_),
    .B(_3648_),
    .CO(_3649_),
    .S(_3650_));
 HA_X1 _8421_ (.A(_3651_),
    .B(_3652_),
    .CO(_3653_),
    .S(_3654_));
 HA_X1 _8422_ (.A(_3655_),
    .B(_3656_),
    .CO(_3657_),
    .S(_3658_));
 HA_X1 _8423_ (.A(_3659_),
    .B(_3660_),
    .CO(_3661_),
    .S(_3662_));
 HA_X1 _8424_ (.A(_2963_),
    .B(_2953_),
    .CO(_3663_),
    .S(_3664_));
 HA_X1 _8425_ (.A(_3665_),
    .B(_3666_),
    .CO(_3667_),
    .S(_3668_));
 HA_X1 _8426_ (.A(_3669_),
    .B(_3670_),
    .CO(_3671_),
    .S(_3672_));
 HA_X1 _8427_ (.A(_3673_),
    .B(_3670_),
    .CO(_3674_),
    .S(_3675_));
 HA_X1 _8428_ (.A(_3676_),
    .B(_3670_),
    .CO(_3677_),
    .S(_3678_));
 HA_X1 _8429_ (.A(_3679_),
    .B(_3670_),
    .CO(_3680_),
    .S(_3681_));
 HA_X1 _8430_ (.A(_3682_),
    .B(_3670_),
    .CO(_3683_),
    .S(_3684_));
 HA_X1 _8431_ (.A(_3685_),
    .B(net228),
    .CO(_3687_),
    .S(_3688_));
 HA_X1 _8432_ (.A(_3689_),
    .B(_3670_),
    .CO(_3690_),
    .S(_3691_));
 HA_X1 _8433_ (.A(_3692_),
    .B(net228),
    .CO(_3693_),
    .S(_3694_));
 HA_X1 _8434_ (.A(_3695_),
    .B(_3670_),
    .CO(_3696_),
    .S(_3697_));
 HA_X1 _8435_ (.A(_3698_),
    .B(_3670_),
    .CO(_3699_),
    .S(_3700_));
 HA_X1 _8436_ (.A(_3701_),
    .B(_3670_),
    .CO(_3702_),
    .S(_3703_));
 HA_X1 _8437_ (.A(_3704_),
    .B(_3686_),
    .CO(_3705_),
    .S(_3706_));
 HA_X1 _8438_ (.A(_3707_),
    .B(_3670_),
    .CO(_3708_),
    .S(_3709_));
 HA_X1 _8439_ (.A(_3710_),
    .B(_3686_),
    .CO(_3711_),
    .S(_3712_));
 HA_X1 _8440_ (.A(_3713_),
    .B(_3714_),
    .CO(_3715_),
    .S(_3716_));
 HA_X1 _8441_ (.A(_3717_),
    .B(_3718_),
    .CO(_3719_),
    .S(_3720_));
 HA_X1 _8442_ (.A(_3721_),
    .B(_3539_),
    .CO(_3722_),
    .S(_3723_));
 HA_X1 _8443_ (.A(_3724_),
    .B(_3725_),
    .CO(_3726_),
    .S(_3727_));
 HA_X1 _8444_ (.A(_3728_),
    .B(_3729_),
    .CO(_3730_),
    .S(_3731_));
 HA_X1 _8445_ (.A(_3732_),
    .B(_3733_),
    .CO(_3734_),
    .S(_3735_));
 HA_X1 _8446_ (.A(_3736_),
    .B(_3737_),
    .CO(_3738_),
    .S(_3739_));
 HA_X1 _8447_ (.A(_2957_),
    .B(_2965_),
    .CO(_3740_),
    .S(_3741_));
 HA_X1 _8448_ (.A(_3538_),
    .B(_3648_),
    .CO(_2954_),
    .S(_3742_));
 HA_X1 _8449_ (.A(_3743_),
    .B(_3540_),
    .CO(_2983_),
    .S(_3744_));
 HA_X1 _8450_ (.A(_3745_),
    .B(_3746_),
    .CO(_3747_),
    .S(_3748_));
 HA_X1 _8451_ (.A(_3749_),
    .B(_3750_),
    .CO(_3751_),
    .S(_3752_));
 HA_X1 _8452_ (.A(_3753_),
    .B(_3754_),
    .CO(_3755_),
    .S(_3756_));
 HA_X1 _8453_ (.A(_3757_),
    .B(_3758_),
    .CO(_3759_),
    .S(_3760_));
 HA_X1 _8454_ (.A(_3762_),
    .B(_3761_),
    .CO(_3763_),
    .S(_3764_));
 HA_X1 _8455_ (.A(_3765_),
    .B(_3766_),
    .CO(_3767_),
    .S(_3768_));
 HA_X1 _8456_ (.A(_3769_),
    .B(_3770_),
    .CO(_3771_),
    .S(_3772_));
 HA_X1 _8457_ (.A(_3769_),
    .B(_3770_),
    .CO(_3773_),
    .S(_3774_));
 HA_X1 _8458_ (.A(_3775_),
    .B(_3776_),
    .CO(_3777_),
    .S(_3778_));
 HA_X1 _8459_ (.A(_3779_),
    .B(_3780_),
    .CO(_3781_),
    .S(_3782_));
 HA_X1 _8460_ (.A(_3783_),
    .B(_3784_),
    .CO(_3785_),
    .S(_3786_));
 HA_X1 _8461_ (.A(_3787_),
    .B(_3788_),
    .CO(_3789_),
    .S(_3790_));
 HA_X1 _8462_ (.A(_3791_),
    .B(_3792_),
    .CO(_3793_),
    .S(_3794_));
 HA_X1 _8463_ (.A(_3795_),
    .B(_3796_),
    .CO(_3797_),
    .S(_3798_));
 HA_X1 _8464_ (.A(_3799_),
    .B(_3800_),
    .CO(_3801_),
    .S(_3802_));
 HA_X1 _8465_ (.A(_3803_),
    .B(_3804_),
    .CO(_3805_),
    .S(_3806_));
 HA_X1 _8466_ (.A(_3803_),
    .B(_3804_),
    .CO(_3807_),
    .S(_3808_));
 HA_X1 _8467_ (.A(_3809_),
    .B(_3810_),
    .CO(_3811_),
    .S(_3812_));
 HA_X1 _8468_ (.A(_3813_),
    .B(_3814_),
    .CO(_3815_),
    .S(_3816_));
 HA_X1 _8469_ (.A(_3817_),
    .B(_3818_),
    .CO(_3819_),
    .S(_3820_));
 HA_X1 _8470_ (.A(_3821_),
    .B(_3822_),
    .CO(_3823_),
    .S(_3824_));
 HA_X1 _8471_ (.A(_3825_),
    .B(_3826_),
    .CO(_3827_),
    .S(_3828_));
 HA_X1 _8472_ (.A(_3829_),
    .B(_3830_),
    .CO(_3831_),
    .S(_3832_));
 HA_X1 _8473_ (.A(_3833_),
    .B(_3834_),
    .CO(_3835_),
    .S(_3836_));
 HA_X1 _8474_ (.A(_3837_),
    .B(_3838_),
    .CO(_3839_),
    .S(_3840_));
 HA_X1 _8475_ (.A(_3841_),
    .B(_3842_),
    .CO(_3843_),
    .S(_3844_));
 HA_X1 _8476_ (.A(_2972_),
    .B(_2973_),
    .CO(_3845_),
    .S(_3846_));
 HA_X1 _8477_ (.A(_3847_),
    .B(_3848_),
    .CO(_3849_),
    .S(_3850_));
 HA_X1 _8478_ (.A(_3851_),
    .B(_3852_),
    .CO(_3853_),
    .S(_3854_));
 HA_X1 _8479_ (.A(_3855_),
    .B(net1),
    .CO(_3857_),
    .S(_3858_));
 HA_X1 _8480_ (.A(_3859_),
    .B(net1),
    .CO(_3860_),
    .S(_3861_));
 HA_X1 _8481_ (.A(_3862_),
    .B(net1),
    .CO(_3863_),
    .S(_3864_));
 HA_X1 _8482_ (.A(_3865_),
    .B(net2),
    .CO(_3866_),
    .S(_3867_));
 HA_X1 _8483_ (.A(_3868_),
    .B(net2),
    .CO(_3869_),
    .S(_3870_));
 HA_X1 _8484_ (.A(_3871_),
    .B(net2),
    .CO(_3872_),
    .S(_3873_));
 HA_X1 _8485_ (.A(_3874_),
    .B(net229),
    .CO(_3876_),
    .S(_3877_));
 HA_X1 _8486_ (.A(_3878_),
    .B(net2),
    .CO(_3879_),
    .S(_3880_));
 HA_X1 _8487_ (.A(_3881_),
    .B(_3875_),
    .CO(_3882_),
    .S(_3883_));
 HA_X1 _8488_ (.A(_3884_),
    .B(_3856_),
    .CO(_3885_),
    .S(_3886_));
 HA_X1 _8489_ (.A(_3887_),
    .B(_3856_),
    .CO(_3888_),
    .S(_3889_));
 HA_X1 _8490_ (.A(_3890_),
    .B(_3856_),
    .CO(_3891_),
    .S(_3892_));
 HA_X1 _8491_ (.A(_3893_),
    .B(_3875_),
    .CO(_3894_),
    .S(_3895_));
 HA_X1 _8492_ (.A(_3896_),
    .B(_3856_),
    .CO(_3897_),
    .S(_3898_));
 HA_X1 _8493_ (.A(_3899_),
    .B(_3900_),
    .CO(_3901_),
    .S(_3902_));
 HA_X1 _8494_ (.A(_3903_),
    .B(_3904_),
    .CO(_3905_),
    .S(_3906_));
 HA_X1 _8495_ (.A(_3907_),
    .B(_3743_),
    .CO(_3908_),
    .S(_3909_));
 HA_X1 _8496_ (.A(_3910_),
    .B(_3911_),
    .CO(_3912_),
    .S(_3913_));
 HA_X1 _8497_ (.A(_3914_),
    .B(_3915_),
    .CO(_3916_),
    .S(_3917_));
 HA_X1 _8498_ (.A(_3918_),
    .B(_3919_),
    .CO(_3920_),
    .S(_3921_));
 HA_X1 _8499_ (.A(_3922_),
    .B(_3923_),
    .CO(_3924_),
    .S(_3925_));
 HA_X1 _8500_ (.A(_3926_),
    .B(_3927_),
    .CO(_3928_),
    .S(_3929_));
 HA_X1 _8501_ (.A(_2967_),
    .B(_2975_),
    .CO(_3930_),
    .S(_3931_));
 HA_X1 _8502_ (.A(_3742_),
    .B(_3826_),
    .CO(_2964_),
    .S(_3932_));
 HA_X1 _8503_ (.A(_3933_),
    .B(_3744_),
    .CO(_2992_),
    .S(_3934_));
 HA_X1 _8504_ (.A(_3935_),
    .B(_3936_),
    .CO(_3937_),
    .S(_3938_));
 HA_X1 _8505_ (.A(_3939_),
    .B(_3940_),
    .CO(_3941_),
    .S(_3942_));
 HA_X1 _8506_ (.A(_3943_),
    .B(_3944_),
    .CO(_3945_),
    .S(_3946_));
 HA_X1 _8507_ (.A(_3947_),
    .B(_3948_),
    .CO(_3949_),
    .S(_3950_));
 HA_X1 _8508_ (.A(_3951_),
    .B(_3952_),
    .CO(_3953_),
    .S(_3954_));
 HA_X1 _8509_ (.A(_3955_),
    .B(_3956_),
    .CO(_3957_),
    .S(_3958_));
 HA_X1 _8510_ (.A(_3959_),
    .B(_3960_),
    .CO(_3961_),
    .S(_3962_));
 HA_X1 _8511_ (.A(_3964_),
    .B(_3963_),
    .CO(_3965_),
    .S(_3966_));
 HA_X1 _8512_ (.A(_3951_),
    .B(_3952_),
    .CO(_3967_),
    .S(_3968_));
 HA_X1 _8513_ (.A(_3969_),
    .B(_3970_),
    .CO(_3971_),
    .S(_3972_));
 HA_X1 _8514_ (.A(_3973_),
    .B(_3974_),
    .CO(_3975_),
    .S(_3976_));
 HA_X1 _8515_ (.A(_3977_),
    .B(_3978_),
    .CO(_3979_),
    .S(_3980_));
 HA_X1 _8516_ (.A(_3981_),
    .B(_3982_),
    .CO(_3983_),
    .S(_3984_));
 HA_X1 _8517_ (.A(_3985_),
    .B(_3986_),
    .CO(_3987_),
    .S(_3988_));
 HA_X1 _8518_ (.A(_3989_),
    .B(_3990_),
    .CO(_3991_),
    .S(_3992_));
 HA_X1 _8519_ (.A(_3993_),
    .B(_3994_),
    .CO(_3995_),
    .S(_3996_));
 HA_X1 _8520_ (.A(_3997_),
    .B(_3998_),
    .CO(_3999_),
    .S(_4000_));
 HA_X1 _8521_ (.A(_4001_),
    .B(_4002_),
    .CO(_4003_),
    .S(_4004_));
 HA_X1 _8522_ (.A(_4006_),
    .B(_4005_),
    .CO(_4007_),
    .S(_4008_));
 HA_X1 _8523_ (.A(_4009_),
    .B(_4010_),
    .CO(_4011_),
    .S(_4012_));
 HA_X1 _8524_ (.A(_2978_),
    .B(_2979_),
    .CO(_4013_),
    .S(_4014_));
 HA_X1 _8525_ (.A(_4015_),
    .B(_4016_),
    .CO(_4017_),
    .S(_4018_));
 HA_X1 _8526_ (.A(_4019_),
    .B(_4020_),
    .CO(_4021_),
    .S(_4022_));
 HA_X1 _8527_ (.A(_4023_),
    .B(_4024_),
    .CO(_4025_),
    .S(_4026_));
 HA_X1 _8528_ (.A(_4027_),
    .B(_4028_),
    .CO(_4029_),
    .S(_4030_));
 HA_X1 _8529_ (.A(net221),
    .B(_4032_),
    .CO(_4033_),
    .S(_4034_));
 HA_X1 _8530_ (.A(net221),
    .B(_4035_),
    .CO(_4036_),
    .S(_4037_));
 HA_X1 _8531_ (.A(net221),
    .B(_4038_),
    .CO(_4039_),
    .S(_4040_));
 HA_X1 _8532_ (.A(net221),
    .B(_4041_),
    .CO(_4042_),
    .S(_4043_));
 HA_X1 _8533_ (.A(net221),
    .B(_4044_),
    .CO(_4045_),
    .S(_4046_));
 HA_X1 _8534_ (.A(net221),
    .B(_4047_),
    .CO(_4048_),
    .S(_4049_));
 HA_X1 _8535_ (.A(net221),
    .B(_4050_),
    .CO(_4051_),
    .S(_4052_));
 HA_X1 _8536_ (.A(net220),
    .B(_4054_),
    .CO(_4055_),
    .S(_4056_));
 HA_X1 _8537_ (.A(_4057_),
    .B(net225),
    .CO(_4058_),
    .S(_4059_));
 HA_X1 _8538_ (.A(net220),
    .B(_4060_),
    .CO(_4061_),
    .S(_4062_));
 HA_X1 _8539_ (.A(net225),
    .B(_4063_),
    .CO(_4064_),
    .S(_4065_));
 HA_X1 _8540_ (.A(_4031_),
    .B(_4066_),
    .CO(_4067_),
    .S(_4068_));
 HA_X1 _8541_ (.A(_4031_),
    .B(_4069_),
    .CO(_4070_),
    .S(_4071_));
 HA_X1 _8542_ (.A(_4072_),
    .B(_4053_),
    .CO(_4073_),
    .S(_4074_));
 HA_X1 _8543_ (.A(_4075_),
    .B(_4076_),
    .CO(_4077_),
    .S(_4078_));
 HA_X1 _8544_ (.A(_4080_),
    .B(_4079_),
    .CO(_4081_),
    .S(_4082_));
 HA_X1 _8545_ (.A(_4083_),
    .B(_4084_),
    .CO(_4085_),
    .S(_4086_));
 HA_X1 _8546_ (.A(_4087_),
    .B(_4088_),
    .CO(_4089_),
    .S(_4090_));
 HA_X1 _8547_ (.A(_4091_),
    .B(_4092_),
    .CO(_4093_),
    .S(_4094_));
 HA_X1 _8548_ (.A(_4095_),
    .B(_4096_),
    .CO(_4097_),
    .S(_4098_));
 HA_X1 _8549_ (.A(_4100_),
    .B(_4099_),
    .CO(_4101_),
    .S(_4102_));
 HA_X1 _8550_ (.A(_4103_),
    .B(_4104_),
    .CO(_4105_),
    .S(_4106_));
 HA_X1 _8551_ (.A(_2985_),
    .B(_2977_),
    .CO(_4107_),
    .S(_4108_));
 HA_X1 _8552_ (.A(_3932_),
    .B(_3990_),
    .CO(_2974_),
    .S(_4109_));
 HA_X1 _8553_ (.A(_4110_),
    .B(_3934_),
    .CO(_2994_),
    .S(_4111_));
 HA_X1 _8554_ (.A(_4112_),
    .B(_4113_),
    .CO(_4114_),
    .S(_4115_));
 HA_X1 _8555_ (.A(_4116_),
    .B(_4117_),
    .CO(_4118_),
    .S(_4119_));
 HA_X1 _8556_ (.A(_4120_),
    .B(_4121_),
    .CO(_4122_),
    .S(_4123_));
 HA_X1 _8557_ (.A(_4124_),
    .B(_4125_),
    .CO(_4126_),
    .S(_4127_));
 HA_X1 _8558_ (.A(_4128_),
    .B(_4129_),
    .CO(_4130_),
    .S(_4131_));
 HA_X1 _8559_ (.A(_4116_),
    .B(_4117_),
    .CO(_4132_),
    .S(_4133_));
 HA_X1 _8560_ (.A(_4134_),
    .B(_4135_),
    .CO(_4136_),
    .S(_4137_));
 HA_X1 _8561_ (.A(_4138_),
    .B(_4139_),
    .CO(_4140_),
    .S(_4141_));
 HA_X1 _8562_ (.A(_4142_),
    .B(_4143_),
    .CO(_4144_),
    .S(_4145_));
 HA_X1 _8563_ (.A(_4146_),
    .B(_4147_),
    .CO(_4148_),
    .S(_4149_));
 HA_X1 _8564_ (.A(_4150_),
    .B(_4151_),
    .CO(_4152_),
    .S(_4153_));
 HA_X1 _8565_ (.A(_4151_),
    .B(_4150_),
    .CO(_4154_),
    .S(_4155_));
 HA_X1 _8566_ (.A(_4156_),
    .B(_4157_),
    .CO(_4158_),
    .S(_4159_));
 HA_X1 _8567_ (.A(_4160_),
    .B(_4161_),
    .CO(_4162_),
    .S(_4163_));
 HA_X1 _8568_ (.A(_4164_),
    .B(_4165_),
    .CO(_4166_),
    .S(_4167_));
 HA_X1 _8569_ (.A(_4169_),
    .B(_4168_),
    .CO(_4170_),
    .S(_4171_));
 HA_X1 _8570_ (.A(_4172_),
    .B(_4173_),
    .CO(_4174_),
    .S(_4175_));
 HA_X1 _8571_ (.A(_2989_),
    .B(_2982_),
    .CO(_4176_),
    .S(_4177_));
 HA_X1 _8572_ (.A(_4178_),
    .B(_4179_),
    .CO(_4180_),
    .S(_4181_));
 HA_X1 _8573_ (.A(_4182_),
    .B(_4183_),
    .CO(_4184_),
    .S(_4185_));
 HA_X1 _8574_ (.A(_4186_),
    .B(_4187_),
    .CO(_4188_),
    .S(_4189_));
 HA_X1 _8575_ (.A(_4190_),
    .B(_4191_),
    .CO(_4192_),
    .S(_4193_));
 HA_X1 _8576_ (.A(_4194_),
    .B(_4195_),
    .CO(_4196_),
    .S(_4197_));
 HA_X1 _8577_ (.A(net69),
    .B(_4199_),
    .CO(_4200_),
    .S(_4201_));
 HA_X1 _8578_ (.A(net69),
    .B(_4202_),
    .CO(_4203_),
    .S(_4204_));
 HA_X1 _8579_ (.A(net69),
    .B(_4205_),
    .CO(_4206_),
    .S(_4207_));
 HA_X1 _8580_ (.A(net69),
    .B(_4208_),
    .CO(_4209_),
    .S(_4210_));
 HA_X1 _8581_ (.A(net69),
    .B(_4211_),
    .CO(_4212_),
    .S(_4213_));
 HA_X1 _8582_ (.A(net69),
    .B(_4214_),
    .CO(_4215_),
    .S(_4216_));
 HA_X1 _8583_ (.A(net69),
    .B(_4217_),
    .CO(_4218_),
    .S(_4219_));
 HA_X1 _8584_ (.A(net277),
    .B(_4220_),
    .CO(_4221_),
    .S(_4222_));
 HA_X1 _8585_ (.A(_4223_),
    .B(_4224_),
    .CO(_4225_),
    .S(_4226_));
 HA_X1 _8586_ (.A(net277),
    .B(_4227_),
    .CO(_4228_),
    .S(_4229_));
 HA_X1 _8587_ (.A(_4223_),
    .B(_4230_),
    .CO(_4231_),
    .S(_4232_));
 HA_X1 _8588_ (.A(_4198_),
    .B(_4233_),
    .CO(_4234_),
    .S(_4235_));
 HA_X1 _8589_ (.A(_4198_),
    .B(_4236_),
    .CO(_4237_),
    .S(_4238_));
 HA_X1 _8590_ (.A(_4198_),
    .B(_4239_),
    .CO(_4240_),
    .S(_4241_));
 HA_X1 _8591_ (.A(_4242_),
    .B(_4243_),
    .CO(_4244_),
    .S(_4245_));
 HA_X1 _8592_ (.A(_4079_),
    .B(_4080_),
    .CO(_4246_),
    .S(_4247_));
 HA_X1 _8593_ (.A(_4248_),
    .B(_3933_),
    .CO(_4249_),
    .S(_4250_));
 HA_X1 _8594_ (.A(_4251_),
    .B(_4252_),
    .CO(_4253_),
    .S(_4254_));
 HA_X1 _8595_ (.A(_4110_),
    .B(_4255_),
    .CO(_4256_),
    .S(_4257_));
 HA_X1 _8596_ (.A(_4259_),
    .B(_4258_),
    .CO(_4260_),
    .S(_4261_));
 HA_X1 _8597_ (.A(_4262_),
    .B(_4263_),
    .CO(_4264_),
    .S(_4265_));
 HA_X1 _8598_ (.A(_4266_),
    .B(_4267_),
    .CO(_4268_),
    .S(_4269_));
 HA_X1 _8599_ (.A(_4271_),
    .B(_4270_),
    .CO(_4272_),
    .S(_4273_));
 HA_X1 _8600_ (.A(_2987_),
    .B(_3006_),
    .CO(_4274_),
    .S(_4275_));
 HA_X1 _8601_ (.A(_4109_),
    .B(_4194_),
    .CO(_2984_),
    .S(_4276_));
 HA_X1 _8602_ (.A(_4277_),
    .B(_4278_),
    .CO(_4279_),
    .S(_4280_));
 HA_X1 _8603_ (.A(_2991_),
    .B(_2998_),
    .CO(_4281_),
    .S(_4282_));
 HA_X1 _8604_ (.A(_4283_),
    .B(_4284_),
    .CO(_4285_),
    .S(_4286_));
 HA_X1 _8605_ (.A(_4287_),
    .B(_4288_),
    .CO(_4289_),
    .S(_4290_));
 HA_X1 _8606_ (.A(_4291_),
    .B(_4292_),
    .CO(_4293_),
    .S(_4294_));
 HA_X1 _8607_ (.A(_4295_),
    .B(_4296_),
    .CO(_4297_),
    .S(_4298_));
 HA_X1 _8608_ (.A(_4299_),
    .B(_4300_),
    .CO(_4301_),
    .S(_4302_));
 HA_X1 _8609_ (.A(_4303_),
    .B(_4304_),
    .CO(_4305_),
    .S(_4306_));
 HA_X1 _8610_ (.A(_4307_),
    .B(_4308_),
    .CO(_4309_),
    .S(_4310_));
 HA_X1 _8611_ (.A(_4307_),
    .B(_4311_),
    .CO(_4312_),
    .S(_4313_));
 HA_X1 _8612_ (.A(_4314_),
    .B(_4307_),
    .CO(_4315_),
    .S(_4316_));
 HA_X1 _8613_ (.A(_4317_),
    .B(_4307_),
    .CO(_4318_),
    .S(_4319_));
 HA_X1 _8614_ (.A(_4307_),
    .B(_4320_),
    .CO(_4321_),
    .S(_4322_));
 HA_X1 _8615_ (.A(_4307_),
    .B(_4323_),
    .CO(_4324_),
    .S(_4325_));
 HA_X1 _8616_ (.A(_4307_),
    .B(_4326_),
    .CO(_4327_),
    .S(_4328_));
 HA_X1 _8617_ (.A(_4307_),
    .B(_4329_),
    .CO(_4330_),
    .S(_4331_));
 HA_X1 _8618_ (.A(_4307_),
    .B(_4332_),
    .CO(_4333_),
    .S(_4334_));
 HA_X1 _8619_ (.A(_4335_),
    .B(_4336_),
    .CO(_4337_),
    .S(_4338_));
 HA_X1 _8620_ (.A(_4339_),
    .B(_4307_),
    .CO(_4340_),
    .S(_4341_));
 HA_X1 _8621_ (.A(_3003_),
    .B(_3004_),
    .CO(_4342_),
    .S(_4343_));
 HA_X1 _8622_ (.A(net314),
    .B(_3002_),
    .CO(_4345_),
    .S(_4346_));
 HA_X1 _8623_ (.A(_4348_),
    .B(_4347_),
    .CO(_4349_),
    .S(_4350_));
 HA_X1 _8624_ (.A(_4351_),
    .B(_4352_),
    .CO(_4353_),
    .S(_4354_));
 HA_X1 _8625_ (.A(_4355_),
    .B(_4356_),
    .CO(_4357_),
    .S(_4358_));
 HA_X1 _8626_ (.A(_4360_),
    .B(_4359_),
    .CO(_4361_),
    .S(_4362_));
 HA_X1 _8627_ (.A(_4363_),
    .B(_4364_),
    .CO(_4365_),
    .S(_4366_));
 HA_X1 _8628_ (.A(net182),
    .B(_4368_),
    .CO(_4369_),
    .S(_4370_));
 HA_X1 _8629_ (.A(_4371_),
    .B(_4372_),
    .CO(_4373_),
    .S(_4374_));
 HA_X1 _8630_ (.A(_4375_),
    .B(_4376_),
    .CO(_4377_),
    .S(_4378_));
 HA_X1 _8631_ (.A(_4379_),
    .B(_4380_),
    .CO(_4381_),
    .S(_4382_));
 HA_X1 _8632_ (.A(_4383_),
    .B(_4384_),
    .CO(_4385_),
    .S(_4386_));
 HA_X1 _8633_ (.A(_4387_),
    .B(_4388_),
    .CO(_4389_),
    .S(_4390_));
 HA_X1 _8634_ (.A(_4391_),
    .B(_4392_),
    .CO(_4393_),
    .S(_4394_));
 HA_X1 _8635_ (.A(_4395_),
    .B(_4396_),
    .CO(_4397_),
    .S(_4398_));
 HA_X1 _8636_ (.A(_4399_),
    .B(_4400_),
    .CO(_4401_),
    .S(_4402_));
 HA_X1 _8637_ (.A(_4403_),
    .B(_4404_),
    .CO(_4405_),
    .S(_4406_));
 HA_X1 _8638_ (.A(_4407_),
    .B(_4408_),
    .CO(_4409_),
    .S(_4410_));
 HA_X1 _8639_ (.A(_4411_),
    .B(_4412_),
    .CO(_4413_),
    .S(_4414_));
 HA_X1 _8640_ (.A(_4415_),
    .B(_4416_),
    .CO(_4417_),
    .S(_4418_));
 HA_X1 _8641_ (.A(_4419_),
    .B(_4420_),
    .CO(_4421_),
    .S(_4422_));
 HA_X1 _8642_ (.A(_4424_),
    .B(_4423_),
    .CO(_4425_),
    .S(_4426_));
 HA_X1 _8643_ (.A(_4427_),
    .B(_4428_),
    .CO(_4429_),
    .S(_4430_));
 HA_X1 _8644_ (.A(net112),
    .B(_4431_),
    .CO(_4432_),
    .S(_4433_));
 HA_X1 _8645_ (.A(_4435_),
    .B(_4434_),
    .CO(_4436_),
    .S(_4437_));
 HA_X1 _8646_ (.A(_4438_),
    .B(_4439_),
    .CO(_4440_),
    .S(_4441_));
 HA_X1 _8647_ (.A(_4442_),
    .B(_4443_),
    .CO(_4444_),
    .S(_4445_));
 HA_X1 _8648_ (.A(_4446_),
    .B(net103),
    .CO(_4448_),
    .S(_4449_));
 HA_X1 _8649_ (.A(_4450_),
    .B(_4451_),
    .CO(_4452_),
    .S(_4453_));
 HA_X1 _8650_ (.A(_4454_),
    .B(_4455_),
    .CO(_4456_),
    .S(_4457_));
 HA_X1 _8651_ (.A(_4458_),
    .B(_4459_),
    .CO(_4460_),
    .S(_4461_));
 HA_X1 _8652_ (.A(_4462_),
    .B(_4463_),
    .CO(_4464_),
    .S(_4465_));
 HA_X1 _8653_ (.A(_4466_),
    .B(_4467_),
    .CO(_4468_),
    .S(_4469_));
 HA_X1 _8654_ (.A(_4470_),
    .B(_4471_),
    .CO(_4472_),
    .S(_4473_));
 HA_X1 _8655_ (.A(_4474_),
    .B(_4475_),
    .CO(_4476_),
    .S(_4477_));
 HA_X1 _8656_ (.A(_4478_),
    .B(_4479_),
    .CO(_4480_),
    .S(_4481_));
 HA_X1 _8657_ (.A(_4482_),
    .B(_4483_),
    .CO(_4484_),
    .S(_4485_));
 HA_X1 _8658_ (.A(_4486_),
    .B(net157),
    .CO(_4488_),
    .S(_4489_));
 HA_X1 _8659_ (.A(_4490_),
    .B(_4491_),
    .CO(_4492_),
    .S(_4493_));
 HA_X1 _8660_ (.A(_3010_),
    .B(_3008_),
    .CO(_4494_),
    .S(_4495_));
 HA_X1 _8661_ (.A(_4438_),
    .B(_4276_),
    .CO(_3005_),
    .S(_4496_));
 HA_X1 _8662_ (.A(net101),
    .B(_4496_),
    .CO(_3009_),
    .S(net56));
 HA_X1 _8663_ (.A(_4497_),
    .B(_4498_),
    .CO(_4499_),
    .S(_4500_));
 HA_X1 _8664_ (.A(_4502_),
    .B(_4501_),
    .CO(_4503_),
    .S(_4504_));
 HA_X1 _8665_ (.A(net46),
    .B(net47),
    .CO(_4505_),
    .S(_4506_));
 HA_X1 _8666_ (.A(_4507_),
    .B(_4508_),
    .CO(_4509_),
    .S(_4510_));
 HA_X1 _8667_ (.A(_4511_),
    .B(_4512_),
    .CO(_4513_),
    .S(_4514_));
 HA_X1 _8668_ (.A(_4515_),
    .B(_4516_),
    .CO(_4517_),
    .S(_4518_));
 HA_X1 _8669_ (.A(_4520_),
    .B(_4519_),
    .CO(_4521_),
    .S(_4522_));
 HA_X1 _8670_ (.A(_4524_),
    .B(_4523_),
    .CO(_4525_),
    .S(_4526_));
 HA_X1 _8671_ (.A(_4527_),
    .B(_4528_),
    .CO(_4529_),
    .S(_4530_));
 HA_X1 _8672_ (.A(_4523_),
    .B(_4531_),
    .CO(_4532_),
    .S(_4533_));
 HA_X1 _8673_ (.A(_4535_),
    .B(_4534_),
    .CO(_4536_),
    .S(_4537_));
 HA_X1 _8674_ (.A(_4538_),
    .B(_4539_),
    .CO(_4540_),
    .S(_4541_));
 HA_X1 _8675_ (.A(net316),
    .B(_4543_),
    .CO(_4544_),
    .S(_4545_));
 HA_X1 _8676_ (.A(_4546_),
    .B(_4547_),
    .CO(_4548_),
    .S(_4549_));
 HA_X1 _8677_ (.A(net194),
    .B(_4551_),
    .CO(_4552_),
    .S(_4553_));
 HA_X1 _8678_ (.A(net191),
    .B(_4539_),
    .CO(_4555_),
    .S(_4556_));
 HA_X1 _8679_ (.A(_4557_),
    .B(_4558_),
    .CO(_4559_),
    .S(_4560_));
 HA_X1 _8680_ (.A(_4561_),
    .B(_4562_),
    .CO(_4563_),
    .S(_4564_));
 HA_X1 _8681_ (.A(_4111_),
    .B(_4542_),
    .CO(_2999_),
    .S(_4344_));
 NAND2_X4 clone1 (.A1(_1318_),
    .A2(_1319_),
    .ZN(net1));
 NAND2_X2 clone2 (.A1(_1318_),
    .A2(_1319_),
    .ZN(net2));
 BUF_X4 clone18 (.A(_0234_),
    .Z(net18));
 XOR2_X2 clone34 (.A(net131),
    .B(_1152_),
    .Z(net34));
 INV_X4 clone67 (.A(_0234_),
    .ZN(net67));
 BUF_X4 clone68 (.A(_2185_),
    .Z(net68));
 BUF_X8 clone69 (.A(_1791_),
    .Z(net69));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Left_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Left_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Left_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Left_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Left_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Left_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Left_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Left_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Left_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Left_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Left_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Left_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Left_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Left_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Left_143 ();
 CLKBUF_X2 input1 (.A(x_in[0]),
    .Z(net5));
 BUF_X1 input2 (.A(x_in[10]),
    .Z(net6));
 BUF_X1 input3 (.A(x_in[11]),
    .Z(net7));
 BUF_X1 input4 (.A(x_in[12]),
    .Z(net8));
 BUF_X1 input5 (.A(x_in[13]),
    .Z(net11));
 BUF_X1 input6 (.A(x_in[14]),
    .Z(net12));
 BUF_X1 input7 (.A(x_in[15]),
    .Z(net13));
 BUF_X4 input8 (.A(x_in[1]),
    .Z(net14));
 BUF_X2 input9 (.A(x_in[2]),
    .Z(net15));
 BUF_X1 input10 (.A(x_in[3]),
    .Z(net16));
 BUF_X1 input11 (.A(x_in[4]),
    .Z(net19));
 BUF_X1 input12 (.A(x_in[5]),
    .Z(net20));
 BUF_X1 input13 (.A(x_in[6]),
    .Z(net21));
 BUF_X1 input14 (.A(x_in[7]),
    .Z(net22));
 BUF_X1 input15 (.A(x_in[8]),
    .Z(net23));
 BUF_X1 input16 (.A(x_in[9]),
    .Z(net24));
 CLKBUF_X2 input17 (.A(y_in[0]),
    .Z(net25));
 BUF_X1 input18 (.A(y_in[10]),
    .Z(net26));
 BUF_X1 input19 (.A(y_in[11]),
    .Z(net27));
 BUF_X1 input20 (.A(y_in[12]),
    .Z(net28));
 BUF_X1 input21 (.A(y_in[13]),
    .Z(net29));
 BUF_X1 input22 (.A(y_in[14]),
    .Z(net30));
 BUF_X1 input23 (.A(y_in[15]),
    .Z(net31));
 BUF_X2 input24 (.A(y_in[1]),
    .Z(net32));
 CLKBUF_X2 input25 (.A(y_in[2]),
    .Z(net33));
 BUF_X1 input26 (.A(y_in[3]),
    .Z(net35));
 BUF_X1 input27 (.A(y_in[4]),
    .Z(net36));
 BUF_X1 input28 (.A(y_in[5]),
    .Z(net37));
 BUF_X1 input29 (.A(y_in[6]),
    .Z(net38));
 BUF_X1 input30 (.A(y_in[7]),
    .Z(net39));
 BUF_X1 input31 (.A(y_in[8]),
    .Z(net40));
 BUF_X1 input32 (.A(y_in[9]),
    .Z(net41));
 CLKBUF_X2 input33 (.A(z_in[10]),
    .Z(net42));
 BUF_X1 input34 (.A(z_in[11]),
    .Z(net43));
 BUF_X1 input35 (.A(z_in[12]),
    .Z(net44));
 BUF_X1 input36 (.A(z_in[13]),
    .Z(net45));
 BUF_X1 input37 (.A(z_in[14]),
    .Z(net46));
 BUF_X4 input38 (.A(z_in[15]),
    .Z(net47));
 BUF_X8 input39 (.A(z_in[1]),
    .Z(net48));
 BUF_X1 input40 (.A(z_in[2]),
    .Z(net49));
 BUF_X1 input41 (.A(z_in[4]),
    .Z(net50));
 BUF_X1 input42 (.A(z_in[5]),
    .Z(net51));
 BUF_X1 input43 (.A(z_in[6]),
    .Z(net52));
 BUF_X1 input44 (.A(z_in[7]),
    .Z(net53));
 BUF_X2 input45 (.A(z_in[8]),
    .Z(net54));
 CLKBUF_X2 input46 (.A(z_in[9]),
    .Z(net55));
 BUF_X1 output47 (.A(net56),
    .Z(x_out[0]));
 BUF_X1 output48 (.A(net57),
    .Z(x_out[10]));
 BUF_X1 output49 (.A(net58),
    .Z(x_out[11]));
 BUF_X1 output50 (.A(net59),
    .Z(x_out[12]));
 BUF_X1 output51 (.A(net60),
    .Z(x_out[13]));
 BUF_X1 output52 (.A(net61),
    .Z(x_out[14]));
 BUF_X1 output53 (.A(net62),
    .Z(x_out[15]));
 BUF_X1 output54 (.A(net63),
    .Z(x_out[1]));
 BUF_X1 output55 (.A(net64),
    .Z(x_out[2]));
 BUF_X1 output56 (.A(net65),
    .Z(x_out[3]));
 BUF_X1 output57 (.A(net66),
    .Z(x_out[4]));
 BUF_X1 output58 (.A(net70),
    .Z(x_out[5]));
 BUF_X1 output59 (.A(net71),
    .Z(x_out[6]));
 BUF_X1 output60 (.A(net72),
    .Z(x_out[7]));
 BUF_X1 output61 (.A(net73),
    .Z(x_out[8]));
 BUF_X1 output62 (.A(net74),
    .Z(x_out[9]));
 BUF_X1 output63 (.A(net75),
    .Z(y_out[0]));
 BUF_X1 output64 (.A(net76),
    .Z(y_out[10]));
 BUF_X1 output65 (.A(net77),
    .Z(y_out[11]));
 BUF_X1 output66 (.A(net78),
    .Z(y_out[12]));
 BUF_X1 output67 (.A(net79),
    .Z(y_out[13]));
 BUF_X1 output68 (.A(net80),
    .Z(y_out[14]));
 BUF_X1 output69 (.A(net81),
    .Z(y_out[15]));
 BUF_X1 output70 (.A(net82),
    .Z(y_out[1]));
 BUF_X1 output71 (.A(net83),
    .Z(y_out[2]));
 BUF_X1 output72 (.A(net84),
    .Z(y_out[3]));
 BUF_X1 output73 (.A(net85),
    .Z(y_out[4]));
 BUF_X1 output74 (.A(net86),
    .Z(y_out[5]));
 BUF_X1 output75 (.A(net87),
    .Z(y_out[6]));
 BUF_X1 output76 (.A(net88),
    .Z(y_out[7]));
 BUF_X1 output77 (.A(net89),
    .Z(y_out[8]));
 BUF_X1 output78 (.A(net90),
    .Z(y_out[9]));
 BUF_X1 rebuffer1 (.A(_4171_),
    .Z(net91));
 BUF_X1 rebuffer2 (.A(_4530_),
    .Z(net92));
 BUF_X1 rebuffer3 (.A(_4430_),
    .Z(net93));
 BUF_X1 rebuffer4 (.A(_4430_),
    .Z(net94));
 BUF_X2 rebuffer5 (.A(_4422_),
    .Z(net95));
 BUF_X1 rebuffer6 (.A(_4350_),
    .Z(net96));
 BUF_X1 rebuffer7 (.A(_4350_),
    .Z(net97));
 BUF_X2 rebuffer8 (.A(_4294_),
    .Z(net98));
 BUF_X1 rebuffer9 (.A(_4537_),
    .Z(net99));
 BUF_X1 rebuffer10 (.A(net99),
    .Z(net100));
 BUF_X1 rebuffer11 (.A(_4447_),
    .Z(net101));
 BUF_X1 rebuffer12 (.A(_4447_),
    .Z(net102));
 BUF_X1 rebuffer13 (.A(net102),
    .Z(net103));
 BUF_X2 rebuffer14 (.A(_4522_),
    .Z(net104));
 BUF_X1 rebuffer15 (.A(net104),
    .Z(net105));
 BUF_X1 rebuffer16 (.A(_2258_),
    .Z(net106));
 BUF_X1 rebuffer17 (.A(_4394_),
    .Z(net107));
 BUF_X1 rebuffer18 (.A(_4394_),
    .Z(net108));
 BUF_X2 rebuffer19 (.A(_4362_),
    .Z(net109));
 BUF_X1 rebuffer20 (.A(_4514_),
    .Z(net110));
 BUF_X4 rebuffer21 (.A(_2169_),
    .Z(net111));
 BUF_X1 rebuffer22 (.A(_4416_),
    .Z(net112));
 BUF_X1 rebuffer23 (.A(_4416_),
    .Z(net113));
 BUF_X1 rebuffer24 (.A(net113),
    .Z(net114));
 BUF_X1 rebuffer25 (.A(_4362_),
    .Z(net115));
 BUF_X1 rebuffer26 (.A(_4102_),
    .Z(net116));
 BUF_X2 rebuffer27 (.A(_3059_),
    .Z(net117));
 BUF_X2 rebuffer28 (.A(_4416_),
    .Z(net118));
 BUF_X1 rebuffer29 (.A(_4305_),
    .Z(net119));
 BUF_X1 rebuffer30 (.A(_2279_),
    .Z(net120));
 BUF_X4 rebuffer31 (.A(_1369_),
    .Z(net121));
 BUF_X1 rebuffer32 (.A(_2685_),
    .Z(net122));
 BUF_X1 rebuffer33 (.A(net122),
    .Z(net123));
 BUF_X1 rebuffer34 (.A(_2004_),
    .Z(net124));
 BUF_X2 rebuffer35 (.A(_1698_),
    .Z(net125));
 BUF_X1 rebuffer36 (.A(net125),
    .Z(net126));
 BUF_X1 rebuffer37 (.A(_4008_),
    .Z(net127));
 BUF_X2 rebuffer38 (.A(_2699_),
    .Z(net128));
 BUF_X2 rebuffer39 (.A(_2702_),
    .Z(net129));
 BUF_X2 clone40 (.A(_3037_),
    .Z(net130));
 BUF_X2 clone41 (.A(_1058_),
    .Z(net131));
 BUF_X1 rebuffer42 (.A(_2137_),
    .Z(net132));
 BUF_X4 rebuffer43 (.A(_1240_),
    .Z(net133));
 BUF_X1 rebuffer44 (.A(_1705_),
    .Z(net134));
 BUF_X1 rebuffer45 (.A(_2248_),
    .Z(net135));
 BUF_X1 rebuffer46 (.A(_3748_),
    .Z(net136));
 BUF_X4 rebuffer47 (.A(_2800_),
    .Z(net137));
 BUF_X1 rebuffer48 (.A(_3808_),
    .Z(net138));
 BUF_X2 rebuffer49 (.A(_2979_),
    .Z(net139));
 BUF_X2 rebuffer50 (.A(_1432_),
    .Z(net140));
 BUF_X1 rebuffer51 (.A(_4074_),
    .Z(net141));
 BUF_X1 rebuffer52 (.A(net141),
    .Z(net142));
 BUF_X4 rebuffer53 (.A(_2741_),
    .Z(net143));
 BUF_X1 rebuffer54 (.A(_4078_),
    .Z(net144));
 BUF_X1 rebuffer55 (.A(_1489_),
    .Z(net145));
 BUF_X1 rebuffer56 (.A(_2184_),
    .Z(net146));
 BUF_X4 rebuffer57 (.A(_1986_),
    .Z(net147));
 BUF_X1 rebuffer58 (.A(_1882_),
    .Z(net148));
 BUF_X1 rebuffer59 (.A(_2240_),
    .Z(net149));
 BUF_X4 rebuffer66 (.A(_4487_),
    .Z(net156));
 BUF_X1 rebuffer67 (.A(net156),
    .Z(net157));
 BUF_X1 rebuffer68 (.A(_4487_),
    .Z(net158));
 BUF_X2 rebuffer69 (.A(_2760_),
    .Z(net159));
 BUF_X2 rebuffer70 (.A(_2221_),
    .Z(net160));
 BUF_X1 rebuffer71 (.A(_3011_),
    .Z(net161));
 BUF_X2 rebuffer72 (.A(_2721_),
    .Z(net162));
 BUF_X2 rebuffer73 (.A(_3980_),
    .Z(net163));
 BUF_X1 rebuffer74 (.A(net163),
    .Z(net164));
 BUF_X1 rebuffer83 (.A(_2718_),
    .Z(net173));
 BUF_X2 rebuffer91 (.A(_4367_),
    .Z(net181));
 BUF_X1 rebuffer92 (.A(net181),
    .Z(net182));
 BUF_X1 rebuffer93 (.A(_1891_),
    .Z(net183));
 BUF_X2 rebuffer94 (.A(net289),
    .Z(net184));
 BUF_X1 rebuffer95 (.A(_4273_),
    .Z(net185));
 BUF_X1 rebuffer96 (.A(_2005_),
    .Z(net186));
 BUF_X1 rebuffer97 (.A(net186),
    .Z(net187));
 BUF_X2 rebuffer98 (.A(net155),
    .Z(net188));
 BUF_X1 rebuffer99 (.A(_2042_),
    .Z(net189));
 BUF_X2 rebuffer100 (.A(_4554_),
    .Z(net190));
 BUF_X1 rebuffer101 (.A(net190),
    .Z(net191));
 BUF_X1 rebuffer102 (.A(_3007_),
    .Z(net192));
 BUF_X8 rebuffer103 (.A(_4550_),
    .Z(net193));
 BUF_X1 rebuffer104 (.A(net193),
    .Z(net194));
 BUF_X4 rebuffer105 (.A(net230),
    .Z(net195));
 BUF_X1 rebuffer106 (.A(_1897_),
    .Z(net196));
 BUF_X1 rebuffer107 (.A(net196),
    .Z(net197));
 BUF_X2 rebuffer119 (.A(_4430_),
    .Z(net209));
 INV_X4 clone123 (.A(_0052_),
    .ZN(net213));
 BUF_X1 rebuffer124 (.A(_2204_),
    .Z(net214));
 BUF_X4 rebuffer125 (.A(net214),
    .Z(net215));
 BUF_X2 rebuffer126 (.A(net215),
    .Z(net216));
 BUF_X4 rebuffer127 (.A(_2258_),
    .Z(net217));
 BUF_X8 clone128 (.A(_0517_),
    .Z(net218));
 BUF_X8 clone129 (.A(_0900_),
    .Z(net219));
 BUF_X8 clone130 (.A(_1591_),
    .Z(net220));
 BUF_X8 clone131 (.A(_1657_),
    .Z(net221));
 BUF_X1 rebuffer132 (.A(_2183_),
    .Z(net222));
 BUF_X1 rebuffer133 (.A(_2246_),
    .Z(net223));
 BUF_X8 clone134 (.A(_0435_),
    .Z(net224));
 BUF_X8 clone135 (.A(_1657_),
    .Z(net225));
 BUF_X8 clone136 (.A(_1320_),
    .Z(net226));
 BUF_X16 clone137 (.A(_0053_),
    .Z(net227));
 BUF_X16 clone138 (.A(_0901_),
    .Z(net228));
 BUF_X16 clone139 (.A(_1321_),
    .Z(net229));
 BUF_X4 rebuffer140 (.A(_1882_),
    .Z(net230));
 BUF_X2 rebuffer141 (.A(_2815_),
    .Z(net231));
 BUF_X2 rebuffer142 (.A(_4123_),
    .Z(net232));
 BUF_X1 rebuffer143 (.A(_1888_),
    .Z(net233));
 BUF_X1 rebuffer144 (.A(_4068_),
    .Z(net234));
 BUF_X4 rebuffer145 (.A(net154),
    .Z(net235));
 BUF_X1 rebuffer146 (.A(_2070_),
    .Z(net236));
 BUF_X1 rebuffer147 (.A(_2039_),
    .Z(net237));
 BUF_X1 rebuffer155 (.A(_4415_),
    .Z(net245));
 BUF_X1 rebuffer156 (.A(_4437_),
    .Z(net246));
 BUF_X4 rebuffer157 (.A(net204),
    .Z(net247));
 BUF_X1 rebuffer158 (.A(_2797_),
    .Z(net248));
 BUF_X4 rebuffer171 (.A(_2812_),
    .Z(net261));
 BUF_X1 rebuffer172 (.A(_2071_),
    .Z(net262));
 BUF_X1 rebuffer173 (.A(_2229_),
    .Z(net263));
 BUF_X1 rebuffer174 (.A(_2229_),
    .Z(net264));
 BUF_X2 rebuffer175 (.A(_4303_),
    .Z(net265));
 BUF_X1 rebuffer181 (.A(_2596_),
    .Z(net271));
 BUF_X1 rebuffer182 (.A(net271),
    .Z(net272));
 BUF_X1 rebuffer183 (.A(net272),
    .Z(net273));
 BUF_X2 rebuffer184 (.A(_4273_),
    .Z(net274));
 BUF_X1 rebuffer185 (.A(_2068_),
    .Z(net275));
 BUF_X4 clone186 (.A(_2012_),
    .Z(net276));
 BUF_X8 clone187 (.A(_1791_),
    .Z(net277));
 BUF_X1 rebuffer188 (.A(_4167_),
    .Z(net278));
 BUF_X1 rebuffer197 (.A(_2826_),
    .Z(net287));
 BUF_X1 rebuffer198 (.A(net287),
    .Z(net288));
 BUF_X2 rebuffer199 (.A(_4378_),
    .Z(net289));
 BUF_X4 rebuffer200 (.A(_2830_),
    .Z(net290));
 BUF_X1 rebuffer201 (.A(_2229_),
    .Z(net291));
 BUF_X2 rebuffer213 (.A(_3000_),
    .Z(net303));
 BUF_X1 rebuffer61 (.A(_4422_),
    .Z(net153));
 BUF_X4 rebuffer62 (.A(_2045_),
    .Z(net154));
 BUF_X1 rebuffer63 (.A(_2135_),
    .Z(net155));
 BUF_X1 rebuffer76 (.A(_2258_),
    .Z(net168));
 BUF_X1 rebuffer80 (.A(_2742_),
    .Z(net172));
 BUF_X1 rebuffer86 (.A(_2011_),
    .Z(net178));
 BUF_X1 rebuffer88 (.A(_2703_),
    .Z(net180));
 BUF_X1 rebuffer110 (.A(_2824_),
    .Z(net202));
 BUF_X1 rebuffer111 (.A(net202),
    .Z(net203));
 BUF_X4 rebuffer112 (.A(_2083_),
    .Z(net204));
 BUF_X1 rebuffer168 (.A(_4510_),
    .Z(net284));
 BUF_X4 rebuffer169 (.A(_2224_),
    .Z(net285));
 BUF_X1 rebuffer186 (.A(_4499_),
    .Z(net297));
 BUF_X1 rebuffer208 (.A(_4344_),
    .Z(net314));
 BUF_X1 rebuffer209 (.A(_4344_),
    .Z(net315));
 BUF_X1 rebuffer210 (.A(_4542_),
    .Z(net316));
 FILLCELL_X8 FILLER_0_1 ();
 FILLCELL_X4 FILLER_0_9 ();
 FILLCELL_X1 FILLER_0_13 ();
 FILLCELL_X1 FILLER_0_29 ();
 FILLCELL_X1 FILLER_0_33 ();
 FILLCELL_X1 FILLER_0_47 ();
 FILLCELL_X4 FILLER_0_51 ();
 FILLCELL_X2 FILLER_0_55 ();
 FILLCELL_X8 FILLER_0_75 ();
 FILLCELL_X2 FILLER_0_83 ();
 FILLCELL_X1 FILLER_0_85 ();
 FILLCELL_X2 FILLER_0_96 ();
 FILLCELL_X4 FILLER_0_106 ();
 FILLCELL_X2 FILLER_0_110 ();
 FILLCELL_X1 FILLER_0_112 ();
 FILLCELL_X4 FILLER_0_131 ();
 FILLCELL_X2 FILLER_0_135 ();
 FILLCELL_X1 FILLER_0_137 ();
 FILLCELL_X1 FILLER_0_140 ();
 FILLCELL_X1 FILLER_0_157 ();
 FILLCELL_X4 FILLER_0_170 ();
 FILLCELL_X2 FILLER_0_174 ();
 FILLCELL_X1 FILLER_0_176 ();
 FILLCELL_X1 FILLER_0_183 ();
 FILLCELL_X2 FILLER_0_197 ();
 FILLCELL_X1 FILLER_0_217 ();
 FILLCELL_X1 FILLER_0_221 ();
 FILLCELL_X2 FILLER_0_226 ();
 FILLCELL_X1 FILLER_0_235 ();
 FILLCELL_X1 FILLER_0_240 ();
 FILLCELL_X1 FILLER_0_249 ();
 FILLCELL_X1 FILLER_0_285 ();
 FILLCELL_X1 FILLER_0_365 ();
 FILLCELL_X1 FILLER_0_377 ();
 FILLCELL_X2 FILLER_0_394 ();
 FILLCELL_X2 FILLER_0_405 ();
 FILLCELL_X2 FILLER_0_436 ();
 FILLCELL_X2 FILLER_0_451 ();
 FILLCELL_X1 FILLER_0_462 ();
 FILLCELL_X1 FILLER_0_466 ();
 FILLCELL_X1 FILLER_0_478 ();
 FILLCELL_X1 FILLER_0_484 ();
 FILLCELL_X2 FILLER_0_534 ();
 FILLCELL_X8 FILLER_1_1 ();
 FILLCELL_X2 FILLER_1_9 ();
 FILLCELL_X1 FILLER_1_11 ();
 FILLCELL_X4 FILLER_1_32 ();
 FILLCELL_X4 FILLER_1_38 ();
 FILLCELL_X4 FILLER_1_54 ();
 FILLCELL_X2 FILLER_1_58 ();
 FILLCELL_X1 FILLER_1_60 ();
 FILLCELL_X8 FILLER_1_78 ();
 FILLCELL_X2 FILLER_1_98 ();
 FILLCELL_X1 FILLER_1_100 ();
 FILLCELL_X4 FILLER_1_111 ();
 FILLCELL_X2 FILLER_1_115 ();
 FILLCELL_X1 FILLER_1_117 ();
 FILLCELL_X2 FILLER_1_120 ();
 FILLCELL_X4 FILLER_1_132 ();
 FILLCELL_X1 FILLER_1_136 ();
 FILLCELL_X1 FILLER_1_147 ();
 FILLCELL_X2 FILLER_1_150 ();
 FILLCELL_X1 FILLER_1_152 ();
 FILLCELL_X4 FILLER_1_157 ();
 FILLCELL_X1 FILLER_1_161 ();
 FILLCELL_X2 FILLER_1_190 ();
 FILLCELL_X1 FILLER_1_370 ();
 FILLCELL_X1 FILLER_1_398 ();
 FILLCELL_X2 FILLER_1_445 ();
 FILLCELL_X1 FILLER_1_447 ();
 FILLCELL_X4 FILLER_1_451 ();
 FILLCELL_X2 FILLER_1_455 ();
 FILLCELL_X1 FILLER_1_457 ();
 FILLCELL_X1 FILLER_1_461 ();
 FILLCELL_X2 FILLER_1_534 ();
 FILLCELL_X4 FILLER_2_30 ();
 FILLCELL_X1 FILLER_2_34 ();
 FILLCELL_X4 FILLER_2_49 ();
 FILLCELL_X2 FILLER_2_53 ();
 FILLCELL_X1 FILLER_2_55 ();
 FILLCELL_X1 FILLER_2_69 ();
 FILLCELL_X1 FILLER_2_75 ();
 FILLCELL_X1 FILLER_2_83 ();
 FILLCELL_X2 FILLER_2_88 ();
 FILLCELL_X2 FILLER_2_95 ();
 FILLCELL_X8 FILLER_2_104 ();
 FILLCELL_X4 FILLER_2_112 ();
 FILLCELL_X4 FILLER_2_126 ();
 FILLCELL_X2 FILLER_2_130 ();
 FILLCELL_X8 FILLER_2_136 ();
 FILLCELL_X1 FILLER_2_144 ();
 FILLCELL_X4 FILLER_2_155 ();
 FILLCELL_X2 FILLER_2_159 ();
 FILLCELL_X8 FILLER_2_171 ();
 FILLCELL_X4 FILLER_2_179 ();
 FILLCELL_X1 FILLER_2_183 ();
 FILLCELL_X1 FILLER_2_195 ();
 FILLCELL_X1 FILLER_2_222 ();
 FILLCELL_X1 FILLER_2_226 ();
 FILLCELL_X2 FILLER_2_265 ();
 FILLCELL_X1 FILLER_2_278 ();
 FILLCELL_X1 FILLER_2_289 ();
 FILLCELL_X1 FILLER_2_309 ();
 FILLCELL_X1 FILLER_2_340 ();
 FILLCELL_X2 FILLER_2_357 ();
 FILLCELL_X8 FILLER_2_366 ();
 FILLCELL_X2 FILLER_2_374 ();
 FILLCELL_X1 FILLER_2_376 ();
 FILLCELL_X2 FILLER_2_390 ();
 FILLCELL_X1 FILLER_2_392 ();
 FILLCELL_X4 FILLER_2_404 ();
 FILLCELL_X2 FILLER_2_408 ();
 FILLCELL_X1 FILLER_2_410 ();
 FILLCELL_X2 FILLER_2_435 ();
 FILLCELL_X2 FILLER_2_449 ();
 FILLCELL_X1 FILLER_2_495 ();
 FILLCELL_X1 FILLER_2_502 ();
 FILLCELL_X1 FILLER_2_527 ();
 FILLCELL_X2 FILLER_2_533 ();
 FILLCELL_X1 FILLER_2_535 ();
 FILLCELL_X8 FILLER_3_4 ();
 FILLCELL_X4 FILLER_3_22 ();
 FILLCELL_X2 FILLER_3_26 ();
 FILLCELL_X4 FILLER_3_32 ();
 FILLCELL_X1 FILLER_3_36 ();
 FILLCELL_X4 FILLER_3_41 ();
 FILLCELL_X2 FILLER_3_45 ();
 FILLCELL_X1 FILLER_3_56 ();
 FILLCELL_X1 FILLER_3_64 ();
 FILLCELL_X2 FILLER_3_78 ();
 FILLCELL_X1 FILLER_3_80 ();
 FILLCELL_X1 FILLER_3_101 ();
 FILLCELL_X2 FILLER_3_108 ();
 FILLCELL_X4 FILLER_3_121 ();
 FILLCELL_X1 FILLER_3_125 ();
 FILLCELL_X4 FILLER_3_160 ();
 FILLCELL_X2 FILLER_3_164 ();
 FILLCELL_X1 FILLER_3_174 ();
 FILLCELL_X2 FILLER_3_189 ();
 FILLCELL_X2 FILLER_3_229 ();
 FILLCELL_X4 FILLER_3_237 ();
 FILLCELL_X1 FILLER_3_241 ();
 FILLCELL_X1 FILLER_3_296 ();
 FILLCELL_X8 FILLER_3_343 ();
 FILLCELL_X4 FILLER_3_351 ();
 FILLCELL_X2 FILLER_3_366 ();
 FILLCELL_X2 FILLER_3_387 ();
 FILLCELL_X1 FILLER_3_396 ();
 FILLCELL_X1 FILLER_3_423 ();
 FILLCELL_X1 FILLER_3_455 ();
 FILLCELL_X1 FILLER_3_494 ();
 FILLCELL_X1 FILLER_3_512 ();
 FILLCELL_X8 FILLER_4_1 ();
 FILLCELL_X4 FILLER_4_9 ();
 FILLCELL_X1 FILLER_4_13 ();
 FILLCELL_X4 FILLER_4_28 ();
 FILLCELL_X4 FILLER_4_39 ();
 FILLCELL_X2 FILLER_4_43 ();
 FILLCELL_X1 FILLER_4_45 ();
 FILLCELL_X1 FILLER_4_50 ();
 FILLCELL_X2 FILLER_4_54 ();
 FILLCELL_X1 FILLER_4_99 ();
 FILLCELL_X1 FILLER_4_118 ();
 FILLCELL_X2 FILLER_4_126 ();
 FILLCELL_X2 FILLER_4_139 ();
 FILLCELL_X2 FILLER_4_148 ();
 FILLCELL_X4 FILLER_4_175 ();
 FILLCELL_X2 FILLER_4_179 ();
 FILLCELL_X1 FILLER_4_181 ();
 FILLCELL_X8 FILLER_4_184 ();
 FILLCELL_X4 FILLER_4_192 ();
 FILLCELL_X2 FILLER_4_196 ();
 FILLCELL_X1 FILLER_4_198 ();
 FILLCELL_X2 FILLER_4_209 ();
 FILLCELL_X2 FILLER_4_215 ();
 FILLCELL_X2 FILLER_4_225 ();
 FILLCELL_X1 FILLER_4_227 ();
 FILLCELL_X2 FILLER_4_237 ();
 FILLCELL_X2 FILLER_4_265 ();
 FILLCELL_X1 FILLER_4_280 ();
 FILLCELL_X4 FILLER_4_358 ();
 FILLCELL_X1 FILLER_4_362 ();
 FILLCELL_X4 FILLER_4_369 ();
 FILLCELL_X2 FILLER_4_387 ();
 FILLCELL_X2 FILLER_4_391 ();
 FILLCELL_X1 FILLER_4_407 ();
 FILLCELL_X1 FILLER_4_421 ();
 FILLCELL_X1 FILLER_4_437 ();
 FILLCELL_X2 FILLER_4_466 ();
 FILLCELL_X1 FILLER_4_468 ();
 FILLCELL_X4 FILLER_4_483 ();
 FILLCELL_X2 FILLER_4_487 ();
 FILLCELL_X8 FILLER_4_495 ();
 FILLCELL_X2 FILLER_4_503 ();
 FILLCELL_X1 FILLER_4_505 ();
 FILLCELL_X4 FILLER_4_518 ();
 FILLCELL_X8 FILLER_5_1 ();
 FILLCELL_X4 FILLER_5_9 ();
 FILLCELL_X2 FILLER_5_13 ();
 FILLCELL_X2 FILLER_5_31 ();
 FILLCELL_X2 FILLER_5_51 ();
 FILLCELL_X2 FILLER_5_59 ();
 FILLCELL_X1 FILLER_5_66 ();
 FILLCELL_X2 FILLER_5_71 ();
 FILLCELL_X1 FILLER_5_73 ();
 FILLCELL_X8 FILLER_5_115 ();
 FILLCELL_X1 FILLER_5_123 ();
 FILLCELL_X4 FILLER_5_140 ();
 FILLCELL_X1 FILLER_5_144 ();
 FILLCELL_X2 FILLER_5_153 ();
 FILLCELL_X2 FILLER_5_162 ();
 FILLCELL_X1 FILLER_5_164 ();
 FILLCELL_X2 FILLER_5_168 ();
 FILLCELL_X1 FILLER_5_170 ();
 FILLCELL_X4 FILLER_5_190 ();
 FILLCELL_X2 FILLER_5_210 ();
 FILLCELL_X2 FILLER_5_218 ();
 FILLCELL_X2 FILLER_5_224 ();
 FILLCELL_X1 FILLER_5_226 ();
 FILLCELL_X1 FILLER_5_244 ();
 FILLCELL_X1 FILLER_5_258 ();
 FILLCELL_X1 FILLER_5_264 ();
 FILLCELL_X1 FILLER_5_285 ();
 FILLCELL_X1 FILLER_5_327 ();
 FILLCELL_X8 FILLER_5_347 ();
 FILLCELL_X4 FILLER_5_355 ();
 FILLCELL_X1 FILLER_5_359 ();
 FILLCELL_X2 FILLER_5_372 ();
 FILLCELL_X2 FILLER_5_384 ();
 FILLCELL_X2 FILLER_5_395 ();
 FILLCELL_X2 FILLER_5_401 ();
 FILLCELL_X1 FILLER_5_403 ();
 FILLCELL_X4 FILLER_5_444 ();
 FILLCELL_X2 FILLER_5_448 ();
 FILLCELL_X1 FILLER_5_450 ();
 FILLCELL_X1 FILLER_5_453 ();
 FILLCELL_X8 FILLER_5_461 ();
 FILLCELL_X4 FILLER_5_469 ();
 FILLCELL_X1 FILLER_5_473 ();
 FILLCELL_X1 FILLER_5_481 ();
 FILLCELL_X4 FILLER_5_495 ();
 FILLCELL_X16 FILLER_5_519 ();
 FILLCELL_X1 FILLER_5_535 ();
 FILLCELL_X1 FILLER_6_1 ();
 FILLCELL_X1 FILLER_6_5 ();
 FILLCELL_X1 FILLER_6_8 ();
 FILLCELL_X2 FILLER_6_19 ();
 FILLCELL_X2 FILLER_6_35 ();
 FILLCELL_X1 FILLER_6_47 ();
 FILLCELL_X2 FILLER_6_52 ();
 FILLCELL_X2 FILLER_6_64 ();
 FILLCELL_X4 FILLER_6_87 ();
 FILLCELL_X2 FILLER_6_91 ();
 FILLCELL_X8 FILLER_6_96 ();
 FILLCELL_X2 FILLER_6_104 ();
 FILLCELL_X4 FILLER_6_115 ();
 FILLCELL_X1 FILLER_6_119 ();
 FILLCELL_X2 FILLER_6_133 ();
 FILLCELL_X1 FILLER_6_157 ();
 FILLCELL_X4 FILLER_6_176 ();
 FILLCELL_X4 FILLER_6_225 ();
 FILLCELL_X4 FILLER_6_238 ();
 FILLCELL_X2 FILLER_6_242 ();
 FILLCELL_X1 FILLER_6_244 ();
 FILLCELL_X4 FILLER_6_248 ();
 FILLCELL_X2 FILLER_6_252 ();
 FILLCELL_X1 FILLER_6_256 ();
 FILLCELL_X8 FILLER_6_279 ();
 FILLCELL_X2 FILLER_6_287 ();
 FILLCELL_X1 FILLER_6_323 ();
 FILLCELL_X8 FILLER_6_341 ();
 FILLCELL_X1 FILLER_6_349 ();
 FILLCELL_X4 FILLER_6_370 ();
 FILLCELL_X4 FILLER_6_378 ();
 FILLCELL_X2 FILLER_6_424 ();
 FILLCELL_X1 FILLER_6_426 ();
 FILLCELL_X2 FILLER_6_440 ();
 FILLCELL_X1 FILLER_6_446 ();
 FILLCELL_X1 FILLER_6_452 ();
 FILLCELL_X2 FILLER_6_473 ();
 FILLCELL_X2 FILLER_6_485 ();
 FILLCELL_X1 FILLER_6_495 ();
 FILLCELL_X8 FILLER_6_505 ();
 FILLCELL_X2 FILLER_6_513 ();
 FILLCELL_X2 FILLER_6_520 ();
 FILLCELL_X4 FILLER_6_531 ();
 FILLCELL_X1 FILLER_6_535 ();
 FILLCELL_X1 FILLER_7_6 ();
 FILLCELL_X1 FILLER_7_17 ();
 FILLCELL_X1 FILLER_7_21 ();
 FILLCELL_X1 FILLER_7_26 ();
 FILLCELL_X1 FILLER_7_34 ();
 FILLCELL_X2 FILLER_7_39 ();
 FILLCELL_X2 FILLER_7_49 ();
 FILLCELL_X1 FILLER_7_51 ();
 FILLCELL_X2 FILLER_7_55 ();
 FILLCELL_X1 FILLER_7_57 ();
 FILLCELL_X1 FILLER_7_69 ();
 FILLCELL_X2 FILLER_7_84 ();
 FILLCELL_X1 FILLER_7_86 ();
 FILLCELL_X8 FILLER_7_109 ();
 FILLCELL_X1 FILLER_7_117 ();
 FILLCELL_X4 FILLER_7_138 ();
 FILLCELL_X4 FILLER_7_149 ();
 FILLCELL_X1 FILLER_7_156 ();
 FILLCELL_X1 FILLER_7_164 ();
 FILLCELL_X4 FILLER_7_167 ();
 FILLCELL_X4 FILLER_7_175 ();
 FILLCELL_X8 FILLER_7_189 ();
 FILLCELL_X2 FILLER_7_197 ();
 FILLCELL_X1 FILLER_7_199 ();
 FILLCELL_X1 FILLER_7_218 ();
 FILLCELL_X4 FILLER_7_228 ();
 FILLCELL_X2 FILLER_7_232 ();
 FILLCELL_X1 FILLER_7_234 ();
 FILLCELL_X1 FILLER_7_248 ();
 FILLCELL_X2 FILLER_7_256 ();
 FILLCELL_X4 FILLER_7_269 ();
 FILLCELL_X2 FILLER_7_273 ();
 FILLCELL_X1 FILLER_7_302 ();
 FILLCELL_X1 FILLER_7_339 ();
 FILLCELL_X32 FILLER_7_350 ();
 FILLCELL_X16 FILLER_7_382 ();
 FILLCELL_X8 FILLER_7_398 ();
 FILLCELL_X1 FILLER_7_415 ();
 FILLCELL_X4 FILLER_7_434 ();
 FILLCELL_X2 FILLER_7_438 ();
 FILLCELL_X1 FILLER_7_440 ();
 FILLCELL_X1 FILLER_7_474 ();
 FILLCELL_X1 FILLER_7_493 ();
 FILLCELL_X2 FILLER_7_500 ();
 FILLCELL_X2 FILLER_7_519 ();
 FILLCELL_X2 FILLER_7_534 ();
 FILLCELL_X1 FILLER_8_1 ();
 FILLCELL_X2 FILLER_8_22 ();
 FILLCELL_X1 FILLER_8_27 ();
 FILLCELL_X2 FILLER_8_40 ();
 FILLCELL_X4 FILLER_8_52 ();
 FILLCELL_X2 FILLER_8_97 ();
 FILLCELL_X2 FILLER_8_119 ();
 FILLCELL_X1 FILLER_8_137 ();
 FILLCELL_X4 FILLER_8_161 ();
 FILLCELL_X2 FILLER_8_177 ();
 FILLCELL_X1 FILLER_8_179 ();
 FILLCELL_X8 FILLER_8_187 ();
 FILLCELL_X4 FILLER_8_195 ();
 FILLCELL_X2 FILLER_8_199 ();
 FILLCELL_X1 FILLER_8_205 ();
 FILLCELL_X4 FILLER_8_216 ();
 FILLCELL_X2 FILLER_8_220 ();
 FILLCELL_X1 FILLER_8_222 ();
 FILLCELL_X2 FILLER_8_235 ();
 FILLCELL_X1 FILLER_8_237 ();
 FILLCELL_X2 FILLER_8_251 ();
 FILLCELL_X8 FILLER_8_267 ();
 FILLCELL_X2 FILLER_8_275 ();
 FILLCELL_X2 FILLER_8_287 ();
 FILLCELL_X1 FILLER_8_289 ();
 FILLCELL_X1 FILLER_8_292 ();
 FILLCELL_X1 FILLER_8_304 ();
 FILLCELL_X2 FILLER_8_317 ();
 FILLCELL_X1 FILLER_8_319 ();
 FILLCELL_X2 FILLER_8_332 ();
 FILLCELL_X4 FILLER_8_345 ();
 FILLCELL_X2 FILLER_8_349 ();
 FILLCELL_X16 FILLER_8_380 ();
 FILLCELL_X8 FILLER_8_396 ();
 FILLCELL_X4 FILLER_8_404 ();
 FILLCELL_X4 FILLER_8_411 ();
 FILLCELL_X2 FILLER_8_415 ();
 FILLCELL_X1 FILLER_8_417 ();
 FILLCELL_X8 FILLER_8_427 ();
 FILLCELL_X1 FILLER_8_446 ();
 FILLCELL_X4 FILLER_8_454 ();
 FILLCELL_X1 FILLER_8_458 ();
 FILLCELL_X8 FILLER_8_502 ();
 FILLCELL_X2 FILLER_8_510 ();
 FILLCELL_X4 FILLER_8_529 ();
 FILLCELL_X2 FILLER_8_533 ();
 FILLCELL_X1 FILLER_8_535 ();
 FILLCELL_X8 FILLER_9_1 ();
 FILLCELL_X1 FILLER_9_9 ();
 FILLCELL_X1 FILLER_9_12 ();
 FILLCELL_X1 FILLER_9_46 ();
 FILLCELL_X2 FILLER_9_53 ();
 FILLCELL_X2 FILLER_9_57 ();
 FILLCELL_X4 FILLER_9_63 ();
 FILLCELL_X1 FILLER_9_67 ();
 FILLCELL_X1 FILLER_9_70 ();
 FILLCELL_X1 FILLER_9_84 ();
 FILLCELL_X2 FILLER_9_89 ();
 FILLCELL_X1 FILLER_9_91 ();
 FILLCELL_X1 FILLER_9_100 ();
 FILLCELL_X4 FILLER_9_124 ();
 FILLCELL_X2 FILLER_9_128 ();
 FILLCELL_X1 FILLER_9_130 ();
 FILLCELL_X2 FILLER_9_135 ();
 FILLCELL_X1 FILLER_9_137 ();
 FILLCELL_X4 FILLER_9_145 ();
 FILLCELL_X2 FILLER_9_149 ();
 FILLCELL_X2 FILLER_9_154 ();
 FILLCELL_X1 FILLER_9_156 ();
 FILLCELL_X4 FILLER_9_160 ();
 FILLCELL_X1 FILLER_9_164 ();
 FILLCELL_X4 FILLER_9_174 ();
 FILLCELL_X1 FILLER_9_178 ();
 FILLCELL_X16 FILLER_9_196 ();
 FILLCELL_X8 FILLER_9_212 ();
 FILLCELL_X2 FILLER_9_220 ();
 FILLCELL_X1 FILLER_9_222 ();
 FILLCELL_X2 FILLER_9_233 ();
 FILLCELL_X2 FILLER_9_245 ();
 FILLCELL_X1 FILLER_9_247 ();
 FILLCELL_X2 FILLER_9_254 ();
 FILLCELL_X8 FILLER_9_266 ();
 FILLCELL_X4 FILLER_9_274 ();
 FILLCELL_X2 FILLER_9_278 ();
 FILLCELL_X8 FILLER_9_315 ();
 FILLCELL_X1 FILLER_9_323 ();
 FILLCELL_X2 FILLER_9_328 ();
 FILLCELL_X1 FILLER_9_330 ();
 FILLCELL_X2 FILLER_9_348 ();
 FILLCELL_X2 FILLER_9_367 ();
 FILLCELL_X1 FILLER_9_369 ();
 FILLCELL_X16 FILLER_9_382 ();
 FILLCELL_X4 FILLER_9_398 ();
 FILLCELL_X1 FILLER_9_402 ();
 FILLCELL_X4 FILLER_9_412 ();
 FILLCELL_X2 FILLER_9_416 ();
 FILLCELL_X32 FILLER_9_427 ();
 FILLCELL_X4 FILLER_9_462 ();
 FILLCELL_X1 FILLER_9_466 ();
 FILLCELL_X4 FILLER_9_478 ();
 FILLCELL_X2 FILLER_9_482 ();
 FILLCELL_X4 FILLER_9_486 ();
 FILLCELL_X1 FILLER_9_490 ();
 FILLCELL_X16 FILLER_9_498 ();
 FILLCELL_X4 FILLER_9_514 ();
 FILLCELL_X2 FILLER_9_518 ();
 FILLCELL_X8 FILLER_10_1 ();
 FILLCELL_X4 FILLER_10_9 ();
 FILLCELL_X1 FILLER_10_13 ();
 FILLCELL_X2 FILLER_10_21 ();
 FILLCELL_X4 FILLER_10_39 ();
 FILLCELL_X2 FILLER_10_43 ();
 FILLCELL_X2 FILLER_10_52 ();
 FILLCELL_X1 FILLER_10_58 ();
 FILLCELL_X2 FILLER_10_75 ();
 FILLCELL_X1 FILLER_10_77 ();
 FILLCELL_X8 FILLER_10_94 ();
 FILLCELL_X2 FILLER_10_102 ();
 FILLCELL_X1 FILLER_10_104 ();
 FILLCELL_X8 FILLER_10_114 ();
 FILLCELL_X2 FILLER_10_122 ();
 FILLCELL_X1 FILLER_10_139 ();
 FILLCELL_X1 FILLER_10_157 ();
 FILLCELL_X4 FILLER_10_176 ();
 FILLCELL_X4 FILLER_10_185 ();
 FILLCELL_X1 FILLER_10_189 ();
 FILLCELL_X8 FILLER_10_206 ();
 FILLCELL_X4 FILLER_10_214 ();
 FILLCELL_X2 FILLER_10_225 ();
 FILLCELL_X1 FILLER_10_227 ();
 FILLCELL_X4 FILLER_10_232 ();
 FILLCELL_X1 FILLER_10_236 ();
 FILLCELL_X8 FILLER_10_247 ();
 FILLCELL_X2 FILLER_10_255 ();
 FILLCELL_X16 FILLER_10_269 ();
 FILLCELL_X4 FILLER_10_316 ();
 FILLCELL_X4 FILLER_10_324 ();
 FILLCELL_X2 FILLER_10_328 ();
 FILLCELL_X8 FILLER_10_348 ();
 FILLCELL_X2 FILLER_10_356 ();
 FILLCELL_X1 FILLER_10_372 ();
 FILLCELL_X1 FILLER_10_422 ();
 FILLCELL_X16 FILLER_10_434 ();
 FILLCELL_X2 FILLER_10_471 ();
 FILLCELL_X2 FILLER_10_483 ();
 FILLCELL_X2 FILLER_10_494 ();
 FILLCELL_X1 FILLER_10_496 ();
 FILLCELL_X2 FILLER_10_521 ();
 FILLCELL_X4 FILLER_10_532 ();
 FILLCELL_X2 FILLER_11_11 ();
 FILLCELL_X1 FILLER_11_17 ();
 FILLCELL_X2 FILLER_11_26 ();
 FILLCELL_X1 FILLER_11_28 ();
 FILLCELL_X2 FILLER_11_36 ();
 FILLCELL_X4 FILLER_11_46 ();
 FILLCELL_X1 FILLER_11_50 ();
 FILLCELL_X8 FILLER_11_53 ();
 FILLCELL_X2 FILLER_11_64 ();
 FILLCELL_X1 FILLER_11_66 ();
 FILLCELL_X16 FILLER_11_74 ();
 FILLCELL_X4 FILLER_11_90 ();
 FILLCELL_X2 FILLER_11_94 ();
 FILLCELL_X1 FILLER_11_96 ();
 FILLCELL_X1 FILLER_11_107 ();
 FILLCELL_X2 FILLER_11_110 ();
 FILLCELL_X1 FILLER_11_112 ();
 FILLCELL_X1 FILLER_11_120 ();
 FILLCELL_X1 FILLER_11_125 ();
 FILLCELL_X1 FILLER_11_129 ();
 FILLCELL_X4 FILLER_11_153 ();
 FILLCELL_X1 FILLER_11_157 ();
 FILLCELL_X1 FILLER_11_160 ();
 FILLCELL_X2 FILLER_11_175 ();
 FILLCELL_X2 FILLER_11_190 ();
 FILLCELL_X4 FILLER_11_205 ();
 FILLCELL_X2 FILLER_11_227 ();
 FILLCELL_X2 FILLER_11_231 ();
 FILLCELL_X1 FILLER_11_233 ();
 FILLCELL_X8 FILLER_11_244 ();
 FILLCELL_X4 FILLER_11_252 ();
 FILLCELL_X1 FILLER_11_256 ();
 FILLCELL_X4 FILLER_11_267 ();
 FILLCELL_X2 FILLER_11_271 ();
 FILLCELL_X1 FILLER_11_273 ();
 FILLCELL_X1 FILLER_11_309 ();
 FILLCELL_X1 FILLER_11_322 ();
 FILLCELL_X4 FILLER_11_325 ();
 FILLCELL_X2 FILLER_11_329 ();
 FILLCELL_X1 FILLER_11_352 ();
 FILLCELL_X1 FILLER_11_406 ();
 FILLCELL_X4 FILLER_11_418 ();
 FILLCELL_X1 FILLER_11_422 ();
 FILLCELL_X2 FILLER_11_433 ();
 FILLCELL_X1 FILLER_11_435 ();
 FILLCELL_X4 FILLER_11_438 ();
 FILLCELL_X2 FILLER_11_442 ();
 FILLCELL_X2 FILLER_11_462 ();
 FILLCELL_X4 FILLER_11_491 ();
 FILLCELL_X2 FILLER_11_495 ();
 FILLCELL_X1 FILLER_11_497 ();
 FILLCELL_X2 FILLER_11_533 ();
 FILLCELL_X1 FILLER_11_535 ();
 FILLCELL_X2 FILLER_12_1 ();
 FILLCELL_X8 FILLER_12_5 ();
 FILLCELL_X4 FILLER_12_13 ();
 FILLCELL_X4 FILLER_12_42 ();
 FILLCELL_X1 FILLER_12_50 ();
 FILLCELL_X1 FILLER_12_64 ();
 FILLCELL_X8 FILLER_12_128 ();
 FILLCELL_X2 FILLER_12_136 ();
 FILLCELL_X1 FILLER_12_138 ();
 FILLCELL_X1 FILLER_12_146 ();
 FILLCELL_X1 FILLER_12_151 ();
 FILLCELL_X1 FILLER_12_203 ();
 FILLCELL_X2 FILLER_12_209 ();
 FILLCELL_X1 FILLER_12_211 ();
 FILLCELL_X1 FILLER_12_221 ();
 FILLCELL_X2 FILLER_12_235 ();
 FILLCELL_X16 FILLER_12_247 ();
 FILLCELL_X8 FILLER_12_263 ();
 FILLCELL_X2 FILLER_12_271 ();
 FILLCELL_X1 FILLER_12_273 ();
 FILLCELL_X1 FILLER_12_354 ();
 FILLCELL_X2 FILLER_12_374 ();
 FILLCELL_X1 FILLER_12_403 ();
 FILLCELL_X8 FILLER_12_421 ();
 FILLCELL_X4 FILLER_12_429 ();
 FILLCELL_X2 FILLER_12_433 ();
 FILLCELL_X2 FILLER_12_471 ();
 FILLCELL_X2 FILLER_12_498 ();
 FILLCELL_X1 FILLER_12_500 ();
 FILLCELL_X4 FILLER_12_516 ();
 FILLCELL_X2 FILLER_12_523 ();
 FILLCELL_X4 FILLER_12_529 ();
 FILLCELL_X2 FILLER_12_533 ();
 FILLCELL_X1 FILLER_12_535 ();
 FILLCELL_X4 FILLER_13_11 ();
 FILLCELL_X4 FILLER_13_22 ();
 FILLCELL_X1 FILLER_13_26 ();
 FILLCELL_X2 FILLER_13_40 ();
 FILLCELL_X2 FILLER_13_52 ();
 FILLCELL_X8 FILLER_13_57 ();
 FILLCELL_X2 FILLER_13_65 ();
 FILLCELL_X1 FILLER_13_67 ();
 FILLCELL_X8 FILLER_13_77 ();
 FILLCELL_X1 FILLER_13_85 ();
 FILLCELL_X8 FILLER_13_93 ();
 FILLCELL_X4 FILLER_13_106 ();
 FILLCELL_X2 FILLER_13_110 ();
 FILLCELL_X8 FILLER_13_119 ();
 FILLCELL_X2 FILLER_13_130 ();
 FILLCELL_X1 FILLER_13_132 ();
 FILLCELL_X4 FILLER_13_135 ();
 FILLCELL_X2 FILLER_13_139 ();
 FILLCELL_X1 FILLER_13_141 ();
 FILLCELL_X1 FILLER_13_150 ();
 FILLCELL_X1 FILLER_13_155 ();
 FILLCELL_X1 FILLER_13_171 ();
 FILLCELL_X2 FILLER_13_176 ();
 FILLCELL_X1 FILLER_13_178 ();
 FILLCELL_X4 FILLER_13_182 ();
 FILLCELL_X1 FILLER_13_186 ();
 FILLCELL_X2 FILLER_13_194 ();
 FILLCELL_X2 FILLER_13_200 ();
 FILLCELL_X1 FILLER_13_202 ();
 FILLCELL_X1 FILLER_13_243 ();
 FILLCELL_X16 FILLER_13_254 ();
 FILLCELL_X4 FILLER_13_270 ();
 FILLCELL_X2 FILLER_13_274 ();
 FILLCELL_X2 FILLER_13_314 ();
 FILLCELL_X1 FILLER_13_357 ();
 FILLCELL_X1 FILLER_13_364 ();
 FILLCELL_X1 FILLER_13_369 ();
 FILLCELL_X8 FILLER_13_374 ();
 FILLCELL_X2 FILLER_13_382 ();
 FILLCELL_X2 FILLER_13_433 ();
 FILLCELL_X1 FILLER_13_435 ();
 FILLCELL_X4 FILLER_13_438 ();
 FILLCELL_X1 FILLER_13_452 ();
 FILLCELL_X8 FILLER_13_470 ();
 FILLCELL_X2 FILLER_13_506 ();
 FILLCELL_X8 FILLER_13_512 ();
 FILLCELL_X2 FILLER_13_520 ();
 FILLCELL_X1 FILLER_13_522 ();
 FILLCELL_X2 FILLER_13_534 ();
 FILLCELL_X1 FILLER_14_4 ();
 FILLCELL_X8 FILLER_14_7 ();
 FILLCELL_X1 FILLER_14_15 ();
 FILLCELL_X8 FILLER_14_20 ();
 FILLCELL_X1 FILLER_14_28 ();
 FILLCELL_X1 FILLER_14_47 ();
 FILLCELL_X2 FILLER_14_52 ();
 FILLCELL_X1 FILLER_14_54 ();
 FILLCELL_X2 FILLER_14_98 ();
 FILLCELL_X8 FILLER_14_107 ();
 FILLCELL_X4 FILLER_14_115 ();
 FILLCELL_X1 FILLER_14_119 ();
 FILLCELL_X1 FILLER_14_123 ();
 FILLCELL_X4 FILLER_14_139 ();
 FILLCELL_X1 FILLER_14_143 ();
 FILLCELL_X1 FILLER_14_151 ();
 FILLCELL_X2 FILLER_14_155 ();
 FILLCELL_X1 FILLER_14_157 ();
 FILLCELL_X2 FILLER_14_160 ();
 FILLCELL_X1 FILLER_14_170 ();
 FILLCELL_X4 FILLER_14_180 ();
 FILLCELL_X4 FILLER_14_195 ();
 FILLCELL_X1 FILLER_14_199 ();
 FILLCELL_X4 FILLER_14_233 ();
 FILLCELL_X2 FILLER_14_237 ();
 FILLCELL_X16 FILLER_14_246 ();
 FILLCELL_X8 FILLER_14_272 ();
 FILLCELL_X2 FILLER_14_280 ();
 FILLCELL_X1 FILLER_14_282 ();
 FILLCELL_X1 FILLER_14_309 ();
 FILLCELL_X2 FILLER_14_364 ();
 FILLCELL_X4 FILLER_14_378 ();
 FILLCELL_X2 FILLER_14_402 ();
 FILLCELL_X1 FILLER_14_470 ();
 FILLCELL_X4 FILLER_14_476 ();
 FILLCELL_X1 FILLER_14_503 ();
 FILLCELL_X2 FILLER_14_518 ();
 FILLCELL_X2 FILLER_14_534 ();
 FILLCELL_X4 FILLER_15_20 ();
 FILLCELL_X1 FILLER_15_24 ();
 FILLCELL_X2 FILLER_15_30 ();
 FILLCELL_X1 FILLER_15_62 ();
 FILLCELL_X8 FILLER_15_70 ();
 FILLCELL_X2 FILLER_15_78 ();
 FILLCELL_X1 FILLER_15_80 ();
 FILLCELL_X2 FILLER_15_93 ();
 FILLCELL_X2 FILLER_15_117 ();
 FILLCELL_X1 FILLER_15_119 ();
 FILLCELL_X1 FILLER_15_176 ();
 FILLCELL_X4 FILLER_15_179 ();
 FILLCELL_X4 FILLER_15_186 ();
 FILLCELL_X1 FILLER_15_190 ();
 FILLCELL_X1 FILLER_15_204 ();
 FILLCELL_X1 FILLER_15_209 ();
 FILLCELL_X4 FILLER_15_221 ();
 FILLCELL_X2 FILLER_15_225 ();
 FILLCELL_X1 FILLER_15_227 ();
 FILLCELL_X2 FILLER_15_244 ();
 FILLCELL_X16 FILLER_15_262 ();
 FILLCELL_X8 FILLER_15_278 ();
 FILLCELL_X2 FILLER_15_298 ();
 FILLCELL_X1 FILLER_15_300 ();
 FILLCELL_X8 FILLER_15_303 ();
 FILLCELL_X4 FILLER_15_311 ();
 FILLCELL_X1 FILLER_15_315 ();
 FILLCELL_X4 FILLER_15_357 ();
 FILLCELL_X2 FILLER_15_361 ();
 FILLCELL_X1 FILLER_15_363 ();
 FILLCELL_X1 FILLER_15_370 ();
 FILLCELL_X2 FILLER_15_375 ();
 FILLCELL_X2 FILLER_15_389 ();
 FILLCELL_X1 FILLER_15_391 ();
 FILLCELL_X2 FILLER_15_403 ();
 FILLCELL_X1 FILLER_15_405 ();
 FILLCELL_X1 FILLER_15_410 ();
 FILLCELL_X4 FILLER_15_417 ();
 FILLCELL_X4 FILLER_15_431 ();
 FILLCELL_X1 FILLER_15_435 ();
 FILLCELL_X1 FILLER_15_446 ();
 FILLCELL_X1 FILLER_15_450 ();
 FILLCELL_X1 FILLER_15_458 ();
 FILLCELL_X2 FILLER_15_469 ();
 FILLCELL_X1 FILLER_15_471 ();
 FILLCELL_X2 FILLER_15_484 ();
 FILLCELL_X1 FILLER_15_504 ();
 FILLCELL_X16 FILLER_15_515 ();
 FILLCELL_X4 FILLER_15_531 ();
 FILLCELL_X1 FILLER_15_535 ();
 FILLCELL_X4 FILLER_16_4 ();
 FILLCELL_X1 FILLER_16_8 ();
 FILLCELL_X1 FILLER_16_22 ();
 FILLCELL_X2 FILLER_16_27 ();
 FILLCELL_X1 FILLER_16_29 ();
 FILLCELL_X2 FILLER_16_32 ();
 FILLCELL_X1 FILLER_16_34 ();
 FILLCELL_X1 FILLER_16_42 ();
 FILLCELL_X2 FILLER_16_50 ();
 FILLCELL_X2 FILLER_16_59 ();
 FILLCELL_X2 FILLER_16_66 ();
 FILLCELL_X1 FILLER_16_68 ();
 FILLCELL_X1 FILLER_16_78 ();
 FILLCELL_X2 FILLER_16_88 ();
 FILLCELL_X1 FILLER_16_90 ();
 FILLCELL_X16 FILLER_16_108 ();
 FILLCELL_X1 FILLER_16_124 ();
 FILLCELL_X2 FILLER_16_128 ();
 FILLCELL_X8 FILLER_16_137 ();
 FILLCELL_X1 FILLER_16_163 ();
 FILLCELL_X2 FILLER_16_170 ();
 FILLCELL_X1 FILLER_16_183 ();
 FILLCELL_X4 FILLER_16_191 ();
 FILLCELL_X1 FILLER_16_195 ();
 FILLCELL_X2 FILLER_16_207 ();
 FILLCELL_X1 FILLER_16_209 ();
 FILLCELL_X8 FILLER_16_220 ();
 FILLCELL_X1 FILLER_16_228 ();
 FILLCELL_X32 FILLER_16_245 ();
 FILLCELL_X8 FILLER_16_277 ();
 FILLCELL_X4 FILLER_16_285 ();
 FILLCELL_X4 FILLER_16_293 ();
 FILLCELL_X1 FILLER_16_297 ();
 FILLCELL_X1 FILLER_16_307 ();
 FILLCELL_X1 FILLER_16_337 ();
 FILLCELL_X1 FILLER_16_351 ();
 FILLCELL_X1 FILLER_16_359 ();
 FILLCELL_X2 FILLER_16_380 ();
 FILLCELL_X4 FILLER_16_392 ();
 FILLCELL_X4 FILLER_16_410 ();
 FILLCELL_X16 FILLER_16_418 ();
 FILLCELL_X1 FILLER_16_434 ();
 FILLCELL_X8 FILLER_16_437 ();
 FILLCELL_X4 FILLER_16_445 ();
 FILLCELL_X4 FILLER_16_451 ();
 FILLCELL_X2 FILLER_16_455 ();
 FILLCELL_X1 FILLER_16_466 ();
 FILLCELL_X8 FILLER_16_470 ();
 FILLCELL_X2 FILLER_16_481 ();
 FILLCELL_X16 FILLER_16_504 ();
 FILLCELL_X1 FILLER_16_520 ();
 FILLCELL_X8 FILLER_16_524 ();
 FILLCELL_X4 FILLER_16_532 ();
 FILLCELL_X2 FILLER_17_1 ();
 FILLCELL_X1 FILLER_17_16 ();
 FILLCELL_X4 FILLER_17_52 ();
 FILLCELL_X1 FILLER_17_56 ();
 FILLCELL_X8 FILLER_17_79 ();
 FILLCELL_X4 FILLER_17_87 ();
 FILLCELL_X1 FILLER_17_91 ();
 FILLCELL_X8 FILLER_17_135 ();
 FILLCELL_X4 FILLER_17_143 ();
 FILLCELL_X1 FILLER_17_150 ();
 FILLCELL_X1 FILLER_17_161 ();
 FILLCELL_X1 FILLER_17_169 ();
 FILLCELL_X2 FILLER_17_174 ();
 FILLCELL_X1 FILLER_17_185 ();
 FILLCELL_X16 FILLER_17_202 ();
 FILLCELL_X8 FILLER_17_218 ();
 FILLCELL_X4 FILLER_17_226 ();
 FILLCELL_X2 FILLER_17_230 ();
 FILLCELL_X1 FILLER_17_232 ();
 FILLCELL_X8 FILLER_17_237 ();
 FILLCELL_X2 FILLER_17_245 ();
 FILLCELL_X2 FILLER_17_260 ();
 FILLCELL_X4 FILLER_17_272 ();
 FILLCELL_X2 FILLER_17_295 ();
 FILLCELL_X4 FILLER_17_307 ();
 FILLCELL_X1 FILLER_17_321 ();
 FILLCELL_X1 FILLER_17_326 ();
 FILLCELL_X8 FILLER_17_349 ();
 FILLCELL_X2 FILLER_17_357 ();
 FILLCELL_X1 FILLER_17_359 ();
 FILLCELL_X4 FILLER_17_366 ();
 FILLCELL_X4 FILLER_17_378 ();
 FILLCELL_X2 FILLER_17_382 ();
 FILLCELL_X1 FILLER_17_384 ();
 FILLCELL_X2 FILLER_17_394 ();
 FILLCELL_X1 FILLER_17_396 ();
 FILLCELL_X2 FILLER_17_399 ();
 FILLCELL_X1 FILLER_17_401 ();
 FILLCELL_X1 FILLER_17_407 ();
 FILLCELL_X4 FILLER_17_422 ();
 FILLCELL_X16 FILLER_17_446 ();
 FILLCELL_X4 FILLER_17_462 ();
 FILLCELL_X1 FILLER_17_466 ();
 FILLCELL_X2 FILLER_17_486 ();
 FILLCELL_X1 FILLER_17_503 ();
 FILLCELL_X2 FILLER_17_533 ();
 FILLCELL_X1 FILLER_17_535 ();
 FILLCELL_X4 FILLER_18_1 ();
 FILLCELL_X1 FILLER_18_5 ();
 FILLCELL_X2 FILLER_18_18 ();
 FILLCELL_X1 FILLER_18_20 ();
 FILLCELL_X2 FILLER_18_34 ();
 FILLCELL_X1 FILLER_18_48 ();
 FILLCELL_X8 FILLER_18_101 ();
 FILLCELL_X4 FILLER_18_109 ();
 FILLCELL_X2 FILLER_18_113 ();
 FILLCELL_X4 FILLER_18_138 ();
 FILLCELL_X1 FILLER_18_142 ();
 FILLCELL_X4 FILLER_18_148 ();
 FILLCELL_X2 FILLER_18_152 ();
 FILLCELL_X8 FILLER_18_159 ();
 FILLCELL_X2 FILLER_18_167 ();
 FILLCELL_X1 FILLER_18_169 ();
 FILLCELL_X4 FILLER_18_180 ();
 FILLCELL_X2 FILLER_18_184 ();
 FILLCELL_X1 FILLER_18_186 ();
 FILLCELL_X1 FILLER_18_189 ();
 FILLCELL_X2 FILLER_18_193 ();
 FILLCELL_X16 FILLER_18_199 ();
 FILLCELL_X4 FILLER_18_215 ();
 FILLCELL_X1 FILLER_18_219 ();
 FILLCELL_X2 FILLER_18_230 ();
 FILLCELL_X1 FILLER_18_232 ();
 FILLCELL_X4 FILLER_18_243 ();
 FILLCELL_X1 FILLER_18_247 ();
 FILLCELL_X2 FILLER_18_250 ();
 FILLCELL_X1 FILLER_18_252 ();
 FILLCELL_X4 FILLER_18_267 ();
 FILLCELL_X8 FILLER_18_275 ();
 FILLCELL_X4 FILLER_18_299 ();
 FILLCELL_X2 FILLER_18_303 ();
 FILLCELL_X1 FILLER_18_305 ();
 FILLCELL_X1 FILLER_18_309 ();
 FILLCELL_X4 FILLER_18_312 ();
 FILLCELL_X1 FILLER_18_326 ();
 FILLCELL_X4 FILLER_18_341 ();
 FILLCELL_X2 FILLER_18_351 ();
 FILLCELL_X2 FILLER_18_371 ();
 FILLCELL_X1 FILLER_18_373 ();
 FILLCELL_X4 FILLER_18_397 ();
 FILLCELL_X2 FILLER_18_401 ();
 FILLCELL_X2 FILLER_18_416 ();
 FILLCELL_X1 FILLER_18_418 ();
 FILLCELL_X16 FILLER_18_428 ();
 FILLCELL_X8 FILLER_18_444 ();
 FILLCELL_X4 FILLER_18_452 ();
 FILLCELL_X2 FILLER_18_456 ();
 FILLCELL_X1 FILLER_18_458 ();
 FILLCELL_X1 FILLER_18_478 ();
 FILLCELL_X1 FILLER_18_523 ();
 FILLCELL_X2 FILLER_18_534 ();
 FILLCELL_X2 FILLER_19_1 ();
 FILLCELL_X2 FILLER_19_13 ();
 FILLCELL_X8 FILLER_19_63 ();
 FILLCELL_X4 FILLER_19_71 ();
 FILLCELL_X2 FILLER_19_75 ();
 FILLCELL_X2 FILLER_19_86 ();
 FILLCELL_X4 FILLER_19_101 ();
 FILLCELL_X2 FILLER_19_114 ();
 FILLCELL_X2 FILLER_19_123 ();
 FILLCELL_X2 FILLER_19_132 ();
 FILLCELL_X1 FILLER_19_134 ();
 FILLCELL_X1 FILLER_19_142 ();
 FILLCELL_X8 FILLER_19_154 ();
 FILLCELL_X1 FILLER_19_162 ();
 FILLCELL_X16 FILLER_19_192 ();
 FILLCELL_X4 FILLER_19_208 ();
 FILLCELL_X2 FILLER_19_212 ();
 FILLCELL_X1 FILLER_19_214 ();
 FILLCELL_X8 FILLER_19_229 ();
 FILLCELL_X2 FILLER_19_237 ();
 FILLCELL_X1 FILLER_19_239 ();
 FILLCELL_X2 FILLER_19_253 ();
 FILLCELL_X16 FILLER_19_271 ();
 FILLCELL_X1 FILLER_19_296 ();
 FILLCELL_X8 FILLER_19_334 ();
 FILLCELL_X2 FILLER_19_342 ();
 FILLCELL_X16 FILLER_19_370 ();
 FILLCELL_X1 FILLER_19_395 ();
 FILLCELL_X1 FILLER_19_398 ();
 FILLCELL_X4 FILLER_19_403 ();
 FILLCELL_X2 FILLER_19_407 ();
 FILLCELL_X1 FILLER_19_409 ();
 FILLCELL_X2 FILLER_19_414 ();
 FILLCELL_X1 FILLER_19_416 ();
 FILLCELL_X1 FILLER_19_425 ();
 FILLCELL_X1 FILLER_19_440 ();
 FILLCELL_X16 FILLER_19_458 ();
 FILLCELL_X1 FILLER_19_504 ();
 FILLCELL_X2 FILLER_19_511 ();
 FILLCELL_X1 FILLER_19_513 ();
 FILLCELL_X1 FILLER_20_4 ();
 FILLCELL_X1 FILLER_20_40 ();
 FILLCELL_X2 FILLER_20_70 ();
 FILLCELL_X1 FILLER_20_72 ();
 FILLCELL_X1 FILLER_20_77 ();
 FILLCELL_X8 FILLER_20_87 ();
 FILLCELL_X2 FILLER_20_95 ();
 FILLCELL_X4 FILLER_20_104 ();
 FILLCELL_X1 FILLER_20_108 ();
 FILLCELL_X8 FILLER_20_118 ();
 FILLCELL_X1 FILLER_20_126 ();
 FILLCELL_X8 FILLER_20_135 ();
 FILLCELL_X4 FILLER_20_143 ();
 FILLCELL_X1 FILLER_20_147 ();
 FILLCELL_X1 FILLER_20_156 ();
 FILLCELL_X1 FILLER_20_161 ();
 FILLCELL_X1 FILLER_20_188 ();
 FILLCELL_X1 FILLER_20_194 ();
 FILLCELL_X2 FILLER_20_211 ();
 FILLCELL_X4 FILLER_20_225 ();
 FILLCELL_X2 FILLER_20_239 ();
 FILLCELL_X1 FILLER_20_241 ();
 FILLCELL_X2 FILLER_20_257 ();
 FILLCELL_X16 FILLER_20_261 ();
 FILLCELL_X2 FILLER_20_277 ();
 FILLCELL_X1 FILLER_20_279 ();
 FILLCELL_X2 FILLER_20_282 ();
 FILLCELL_X1 FILLER_20_284 ();
 FILLCELL_X1 FILLER_20_292 ();
 FILLCELL_X16 FILLER_20_326 ();
 FILLCELL_X8 FILLER_20_342 ();
 FILLCELL_X2 FILLER_20_386 ();
 FILLCELL_X1 FILLER_20_388 ();
 FILLCELL_X1 FILLER_20_393 ();
 FILLCELL_X2 FILLER_20_404 ();
 FILLCELL_X1 FILLER_20_406 ();
 FILLCELL_X8 FILLER_20_411 ();
 FILLCELL_X1 FILLER_20_419 ();
 FILLCELL_X2 FILLER_20_422 ();
 FILLCELL_X4 FILLER_20_451 ();
 FILLCELL_X8 FILLER_20_462 ();
 FILLCELL_X2 FILLER_20_470 ();
 FILLCELL_X4 FILLER_20_481 ();
 FILLCELL_X1 FILLER_20_485 ();
 FILLCELL_X1 FILLER_20_510 ();
 FILLCELL_X2 FILLER_20_521 ();
 FILLCELL_X4 FILLER_21_1 ();
 FILLCELL_X2 FILLER_21_5 ();
 FILLCELL_X1 FILLER_21_7 ();
 FILLCELL_X2 FILLER_21_26 ();
 FILLCELL_X4 FILLER_21_46 ();
 FILLCELL_X2 FILLER_21_50 ();
 FILLCELL_X1 FILLER_21_52 ();
 FILLCELL_X8 FILLER_21_63 ();
 FILLCELL_X1 FILLER_21_71 ();
 FILLCELL_X16 FILLER_21_74 ();
 FILLCELL_X8 FILLER_21_90 ();
 FILLCELL_X4 FILLER_21_98 ();
 FILLCELL_X2 FILLER_21_102 ();
 FILLCELL_X1 FILLER_21_104 ();
 FILLCELL_X2 FILLER_21_107 ();
 FILLCELL_X1 FILLER_21_109 ();
 FILLCELL_X4 FILLER_21_127 ();
 FILLCELL_X2 FILLER_21_131 ();
 FILLCELL_X2 FILLER_21_137 ();
 FILLCELL_X1 FILLER_21_139 ();
 FILLCELL_X2 FILLER_21_158 ();
 FILLCELL_X4 FILLER_21_163 ();
 FILLCELL_X2 FILLER_21_193 ();
 FILLCELL_X1 FILLER_21_195 ();
 FILLCELL_X8 FILLER_21_206 ();
 FILLCELL_X4 FILLER_21_214 ();
 FILLCELL_X2 FILLER_21_218 ();
 FILLCELL_X1 FILLER_21_220 ();
 FILLCELL_X16 FILLER_21_251 ();
 FILLCELL_X8 FILLER_21_267 ();
 FILLCELL_X4 FILLER_21_275 ();
 FILLCELL_X2 FILLER_21_307 ();
 FILLCELL_X1 FILLER_21_309 ();
 FILLCELL_X8 FILLER_21_312 ();
 FILLCELL_X2 FILLER_21_320 ();
 FILLCELL_X8 FILLER_21_343 ();
 FILLCELL_X16 FILLER_21_363 ();
 FILLCELL_X4 FILLER_21_379 ();
 FILLCELL_X2 FILLER_21_397 ();
 FILLCELL_X1 FILLER_21_435 ();
 FILLCELL_X4 FILLER_21_455 ();
 FILLCELL_X16 FILLER_21_487 ();
 FILLCELL_X4 FILLER_21_503 ();
 FILLCELL_X4 FILLER_21_510 ();
 FILLCELL_X2 FILLER_21_514 ();
 FILLCELL_X1 FILLER_21_535 ();
 FILLCELL_X16 FILLER_22_1 ();
 FILLCELL_X4 FILLER_22_41 ();
 FILLCELL_X8 FILLER_22_49 ();
 FILLCELL_X4 FILLER_22_57 ();
 FILLCELL_X4 FILLER_22_70 ();
 FILLCELL_X8 FILLER_22_87 ();
 FILLCELL_X4 FILLER_22_95 ();
 FILLCELL_X2 FILLER_22_99 ();
 FILLCELL_X1 FILLER_22_101 ();
 FILLCELL_X2 FILLER_22_109 ();
 FILLCELL_X1 FILLER_22_111 ();
 FILLCELL_X4 FILLER_22_114 ();
 FILLCELL_X1 FILLER_22_118 ();
 FILLCELL_X8 FILLER_22_144 ();
 FILLCELL_X1 FILLER_22_152 ();
 FILLCELL_X2 FILLER_22_159 ();
 FILLCELL_X1 FILLER_22_161 ();
 FILLCELL_X2 FILLER_22_182 ();
 FILLCELL_X1 FILLER_22_184 ();
 FILLCELL_X4 FILLER_22_189 ();
 FILLCELL_X4 FILLER_22_206 ();
 FILLCELL_X1 FILLER_22_245 ();
 FILLCELL_X16 FILLER_22_261 ();
 FILLCELL_X4 FILLER_22_277 ();
 FILLCELL_X1 FILLER_22_287 ();
 FILLCELL_X8 FILLER_22_309 ();
 FILLCELL_X4 FILLER_22_317 ();
 FILLCELL_X2 FILLER_22_321 ();
 FILLCELL_X16 FILLER_22_325 ();
 FILLCELL_X2 FILLER_22_341 ();
 FILLCELL_X1 FILLER_22_343 ();
 FILLCELL_X2 FILLER_22_354 ();
 FILLCELL_X1 FILLER_22_356 ();
 FILLCELL_X8 FILLER_22_379 ();
 FILLCELL_X2 FILLER_22_387 ();
 FILLCELL_X4 FILLER_22_399 ();
 FILLCELL_X4 FILLER_22_505 ();
 FILLCELL_X2 FILLER_22_509 ();
 FILLCELL_X1 FILLER_23_1 ();
 FILLCELL_X4 FILLER_23_34 ();
 FILLCELL_X2 FILLER_23_38 ();
 FILLCELL_X4 FILLER_23_59 ();
 FILLCELL_X1 FILLER_23_70 ();
 FILLCELL_X8 FILLER_23_79 ();
 FILLCELL_X4 FILLER_23_87 ();
 FILLCELL_X1 FILLER_23_91 ();
 FILLCELL_X16 FILLER_23_101 ();
 FILLCELL_X2 FILLER_23_117 ();
 FILLCELL_X16 FILLER_23_123 ();
 FILLCELL_X4 FILLER_23_139 ();
 FILLCELL_X2 FILLER_23_143 ();
 FILLCELL_X2 FILLER_23_180 ();
 FILLCELL_X1 FILLER_23_186 ();
 FILLCELL_X4 FILLER_23_200 ();
 FILLCELL_X2 FILLER_23_239 ();
 FILLCELL_X8 FILLER_23_251 ();
 FILLCELL_X4 FILLER_23_259 ();
 FILLCELL_X2 FILLER_23_263 ();
 FILLCELL_X4 FILLER_23_275 ();
 FILLCELL_X4 FILLER_23_289 ();
 FILLCELL_X1 FILLER_23_293 ();
 FILLCELL_X1 FILLER_23_337 ();
 FILLCELL_X32 FILLER_23_340 ();
 FILLCELL_X2 FILLER_23_374 ();
 FILLCELL_X4 FILLER_23_386 ();
 FILLCELL_X1 FILLER_23_394 ();
 FILLCELL_X1 FILLER_23_469 ();
 FILLCELL_X8 FILLER_24_1 ();
 FILLCELL_X2 FILLER_24_9 ();
 FILLCELL_X1 FILLER_24_11 ();
 FILLCELL_X4 FILLER_24_16 ();
 FILLCELL_X4 FILLER_24_24 ();
 FILLCELL_X2 FILLER_24_28 ();
 FILLCELL_X2 FILLER_24_44 ();
 FILLCELL_X1 FILLER_24_46 ();
 FILLCELL_X4 FILLER_24_56 ();
 FILLCELL_X1 FILLER_24_60 ();
 FILLCELL_X4 FILLER_24_79 ();
 FILLCELL_X1 FILLER_24_83 ();
 FILLCELL_X2 FILLER_24_108 ();
 FILLCELL_X16 FILLER_24_122 ();
 FILLCELL_X4 FILLER_24_138 ();
 FILLCELL_X16 FILLER_24_157 ();
 FILLCELL_X4 FILLER_24_173 ();
 FILLCELL_X4 FILLER_24_187 ();
 FILLCELL_X2 FILLER_24_191 ();
 FILLCELL_X1 FILLER_24_205 ();
 FILLCELL_X1 FILLER_24_236 ();
 FILLCELL_X4 FILLER_24_240 ();
 FILLCELL_X1 FILLER_24_244 ();
 FILLCELL_X2 FILLER_24_270 ();
 FILLCELL_X16 FILLER_24_285 ();
 FILLCELL_X4 FILLER_24_301 ();
 FILLCELL_X2 FILLER_24_305 ();
 FILLCELL_X2 FILLER_24_315 ();
 FILLCELL_X8 FILLER_24_356 ();
 FILLCELL_X1 FILLER_24_364 ();
 FILLCELL_X2 FILLER_24_369 ();
 FILLCELL_X4 FILLER_24_375 ();
 FILLCELL_X2 FILLER_24_379 ();
 FILLCELL_X4 FILLER_24_448 ();
 FILLCELL_X1 FILLER_24_452 ();
 FILLCELL_X4 FILLER_24_466 ();
 FILLCELL_X2 FILLER_24_470 ();
 FILLCELL_X1 FILLER_24_472 ();
 FILLCELL_X1 FILLER_24_518 ();
 FILLCELL_X1 FILLER_24_535 ();
 FILLCELL_X1 FILLER_25_1 ();
 FILLCELL_X2 FILLER_25_8 ();
 FILLCELL_X1 FILLER_25_10 ();
 FILLCELL_X1 FILLER_25_32 ();
 FILLCELL_X1 FILLER_25_37 ();
 FILLCELL_X1 FILLER_25_49 ();
 FILLCELL_X1 FILLER_25_56 ();
 FILLCELL_X1 FILLER_25_60 ();
 FILLCELL_X1 FILLER_25_71 ();
 FILLCELL_X8 FILLER_25_76 ();
 FILLCELL_X2 FILLER_25_94 ();
 FILLCELL_X2 FILLER_25_114 ();
 FILLCELL_X1 FILLER_25_125 ();
 FILLCELL_X2 FILLER_25_141 ();
 FILLCELL_X1 FILLER_25_143 ();
 FILLCELL_X1 FILLER_25_233 ();
 FILLCELL_X8 FILLER_25_277 ();
 FILLCELL_X2 FILLER_25_325 ();
 FILLCELL_X1 FILLER_25_327 ();
 FILLCELL_X4 FILLER_25_344 ();
 FILLCELL_X1 FILLER_25_348 ();
 FILLCELL_X4 FILLER_25_360 ();
 FILLCELL_X1 FILLER_25_364 ();
 FILLCELL_X8 FILLER_25_375 ();
 FILLCELL_X4 FILLER_25_383 ();
 FILLCELL_X2 FILLER_25_387 ();
 FILLCELL_X1 FILLER_25_441 ();
 FILLCELL_X1 FILLER_25_459 ();
 FILLCELL_X8 FILLER_25_476 ();
 FILLCELL_X4 FILLER_25_484 ();
 FILLCELL_X2 FILLER_25_488 ();
 FILLCELL_X1 FILLER_25_490 ();
 FILLCELL_X2 FILLER_25_510 ();
 FILLCELL_X2 FILLER_25_518 ();
 FILLCELL_X4 FILLER_25_530 ();
 FILLCELL_X2 FILLER_25_534 ();
 FILLCELL_X8 FILLER_26_1 ();
 FILLCELL_X4 FILLER_26_9 ();
 FILLCELL_X1 FILLER_26_20 ();
 FILLCELL_X2 FILLER_26_30 ();
 FILLCELL_X2 FILLER_26_36 ();
 FILLCELL_X1 FILLER_26_49 ();
 FILLCELL_X2 FILLER_26_66 ();
 FILLCELL_X2 FILLER_26_71 ();
 FILLCELL_X2 FILLER_26_79 ();
 FILLCELL_X1 FILLER_26_90 ();
 FILLCELL_X2 FILLER_26_120 ();
 FILLCELL_X2 FILLER_26_128 ();
 FILLCELL_X4 FILLER_26_140 ();
 FILLCELL_X2 FILLER_26_144 ();
 FILLCELL_X2 FILLER_26_151 ();
 FILLCELL_X1 FILLER_26_153 ();
 FILLCELL_X2 FILLER_26_168 ();
 FILLCELL_X16 FILLER_26_172 ();
 FILLCELL_X8 FILLER_26_188 ();
 FILLCELL_X1 FILLER_26_196 ();
 FILLCELL_X1 FILLER_26_211 ();
 FILLCELL_X8 FILLER_26_219 ();
 FILLCELL_X1 FILLER_26_227 ();
 FILLCELL_X1 FILLER_26_234 ();
 FILLCELL_X2 FILLER_26_237 ();
 FILLCELL_X4 FILLER_26_248 ();
 FILLCELL_X1 FILLER_26_252 ();
 FILLCELL_X2 FILLER_26_285 ();
 FILLCELL_X1 FILLER_26_287 ();
 FILLCELL_X8 FILLER_26_297 ();
 FILLCELL_X1 FILLER_26_311 ();
 FILLCELL_X16 FILLER_26_316 ();
 FILLCELL_X1 FILLER_26_332 ();
 FILLCELL_X2 FILLER_26_355 ();
 FILLCELL_X1 FILLER_26_357 ();
 FILLCELL_X2 FILLER_26_373 ();
 FILLCELL_X1 FILLER_26_375 ();
 FILLCELL_X2 FILLER_26_390 ();
 FILLCELL_X1 FILLER_26_435 ();
 FILLCELL_X1 FILLER_26_454 ();
 FILLCELL_X8 FILLER_26_480 ();
 FILLCELL_X4 FILLER_26_488 ();
 FILLCELL_X2 FILLER_26_492 ();
 FILLCELL_X8 FILLER_26_513 ();
 FILLCELL_X8 FILLER_26_523 ();
 FILLCELL_X4 FILLER_26_531 ();
 FILLCELL_X1 FILLER_26_535 ();
 FILLCELL_X2 FILLER_27_1 ();
 FILLCELL_X2 FILLER_27_13 ();
 FILLCELL_X1 FILLER_27_30 ();
 FILLCELL_X2 FILLER_27_62 ();
 FILLCELL_X1 FILLER_27_64 ();
 FILLCELL_X8 FILLER_27_72 ();
 FILLCELL_X4 FILLER_27_80 ();
 FILLCELL_X2 FILLER_27_84 ();
 FILLCELL_X4 FILLER_27_96 ();
 FILLCELL_X1 FILLER_27_100 ();
 FILLCELL_X4 FILLER_27_122 ();
 FILLCELL_X1 FILLER_27_126 ();
 FILLCELL_X8 FILLER_27_136 ();
 FILLCELL_X2 FILLER_27_144 ();
 FILLCELL_X1 FILLER_27_146 ();
 FILLCELL_X4 FILLER_27_152 ();
 FILLCELL_X8 FILLER_27_163 ();
 FILLCELL_X4 FILLER_27_171 ();
 FILLCELL_X2 FILLER_27_175 ();
 FILLCELL_X16 FILLER_27_187 ();
 FILLCELL_X1 FILLER_27_209 ();
 FILLCELL_X4 FILLER_27_223 ();
 FILLCELL_X2 FILLER_27_227 ();
 FILLCELL_X8 FILLER_27_238 ();
 FILLCELL_X4 FILLER_27_246 ();
 FILLCELL_X2 FILLER_27_250 ();
 FILLCELL_X2 FILLER_27_258 ();
 FILLCELL_X2 FILLER_27_279 ();
 FILLCELL_X2 FILLER_27_289 ();
 FILLCELL_X1 FILLER_27_291 ();
 FILLCELL_X8 FILLER_27_344 ();
 FILLCELL_X4 FILLER_27_352 ();
 FILLCELL_X1 FILLER_27_370 ();
 FILLCELL_X16 FILLER_27_378 ();
 FILLCELL_X8 FILLER_27_394 ();
 FILLCELL_X4 FILLER_27_402 ();
 FILLCELL_X1 FILLER_27_406 ();
 FILLCELL_X4 FILLER_27_416 ();
 FILLCELL_X16 FILLER_27_473 ();
 FILLCELL_X4 FILLER_27_489 ();
 FILLCELL_X2 FILLER_27_493 ();
 FILLCELL_X2 FILLER_27_498 ();
 FILLCELL_X1 FILLER_27_507 ();
 FILLCELL_X2 FILLER_27_510 ();
 FILLCELL_X1 FILLER_27_512 ();
 FILLCELL_X8 FILLER_27_523 ();
 FILLCELL_X4 FILLER_27_531 ();
 FILLCELL_X1 FILLER_27_535 ();
 FILLCELL_X8 FILLER_28_1 ();
 FILLCELL_X2 FILLER_28_9 ();
 FILLCELL_X2 FILLER_28_18 ();
 FILLCELL_X1 FILLER_28_20 ();
 FILLCELL_X2 FILLER_28_38 ();
 FILLCELL_X1 FILLER_28_40 ();
 FILLCELL_X2 FILLER_28_44 ();
 FILLCELL_X1 FILLER_28_46 ();
 FILLCELL_X1 FILLER_28_52 ();
 FILLCELL_X8 FILLER_28_78 ();
 FILLCELL_X1 FILLER_28_94 ();
 FILLCELL_X2 FILLER_28_106 ();
 FILLCELL_X4 FILLER_28_112 ();
 FILLCELL_X1 FILLER_28_116 ();
 FILLCELL_X4 FILLER_28_127 ();
 FILLCELL_X2 FILLER_28_141 ();
 FILLCELL_X1 FILLER_28_143 ();
 FILLCELL_X16 FILLER_28_162 ();
 FILLCELL_X4 FILLER_28_181 ();
 FILLCELL_X1 FILLER_28_191 ();
 FILLCELL_X4 FILLER_28_196 ();
 FILLCELL_X8 FILLER_28_211 ();
 FILLCELL_X2 FILLER_28_219 ();
 FILLCELL_X1 FILLER_28_221 ();
 FILLCELL_X2 FILLER_28_226 ();
 FILLCELL_X2 FILLER_28_247 ();
 FILLCELL_X16 FILLER_28_265 ();
 FILLCELL_X4 FILLER_28_281 ();
 FILLCELL_X2 FILLER_28_289 ();
 FILLCELL_X4 FILLER_28_302 ();
 FILLCELL_X2 FILLER_28_306 ();
 FILLCELL_X1 FILLER_28_308 ();
 FILLCELL_X4 FILLER_28_311 ();
 FILLCELL_X2 FILLER_28_315 ();
 FILLCELL_X1 FILLER_28_319 ();
 FILLCELL_X8 FILLER_28_330 ();
 FILLCELL_X4 FILLER_28_338 ();
 FILLCELL_X8 FILLER_28_352 ();
 FILLCELL_X4 FILLER_28_372 ();
 FILLCELL_X2 FILLER_28_376 ();
 FILLCELL_X1 FILLER_28_378 ();
 FILLCELL_X16 FILLER_28_387 ();
 FILLCELL_X8 FILLER_28_403 ();
 FILLCELL_X4 FILLER_28_411 ();
 FILLCELL_X1 FILLER_28_418 ();
 FILLCELL_X4 FILLER_28_448 ();
 FILLCELL_X1 FILLER_28_452 ();
 FILLCELL_X1 FILLER_28_456 ();
 FILLCELL_X1 FILLER_28_477 ();
 FILLCELL_X1 FILLER_28_491 ();
 FILLCELL_X4 FILLER_28_531 ();
 FILLCELL_X1 FILLER_28_535 ();
 FILLCELL_X4 FILLER_29_1 ();
 FILLCELL_X1 FILLER_29_5 ();
 FILLCELL_X4 FILLER_29_26 ();
 FILLCELL_X1 FILLER_29_30 ();
 FILLCELL_X8 FILLER_29_43 ();
 FILLCELL_X2 FILLER_29_51 ();
 FILLCELL_X4 FILLER_29_67 ();
 FILLCELL_X1 FILLER_29_71 ();
 FILLCELL_X4 FILLER_29_112 ();
 FILLCELL_X2 FILLER_29_118 ();
 FILLCELL_X1 FILLER_29_120 ();
 FILLCELL_X4 FILLER_29_125 ();
 FILLCELL_X1 FILLER_29_129 ();
 FILLCELL_X4 FILLER_29_140 ();
 FILLCELL_X2 FILLER_29_154 ();
 FILLCELL_X1 FILLER_29_156 ();
 FILLCELL_X4 FILLER_29_174 ();
 FILLCELL_X2 FILLER_29_178 ();
 FILLCELL_X4 FILLER_29_198 ();
 FILLCELL_X1 FILLER_29_202 ();
 FILLCELL_X2 FILLER_29_207 ();
 FILLCELL_X2 FILLER_29_216 ();
 FILLCELL_X1 FILLER_29_224 ();
 FILLCELL_X16 FILLER_29_235 ();
 FILLCELL_X1 FILLER_29_263 ();
 FILLCELL_X16 FILLER_29_266 ();
 FILLCELL_X2 FILLER_29_282 ();
 FILLCELL_X4 FILLER_29_294 ();
 FILLCELL_X1 FILLER_29_308 ();
 FILLCELL_X2 FILLER_29_319 ();
 FILLCELL_X1 FILLER_29_321 ();
 FILLCELL_X4 FILLER_29_345 ();
 FILLCELL_X2 FILLER_29_349 ();
 FILLCELL_X1 FILLER_29_351 ();
 FILLCELL_X8 FILLER_29_362 ();
 FILLCELL_X2 FILLER_29_370 ();
 FILLCELL_X1 FILLER_29_372 ();
 FILLCELL_X1 FILLER_29_386 ();
 FILLCELL_X16 FILLER_29_397 ();
 FILLCELL_X2 FILLER_29_413 ();
 FILLCELL_X1 FILLER_29_415 ();
 FILLCELL_X16 FILLER_29_426 ();
 FILLCELL_X1 FILLER_29_442 ();
 FILLCELL_X1 FILLER_29_477 ();
 FILLCELL_X1 FILLER_29_509 ();
 FILLCELL_X4 FILLER_29_530 ();
 FILLCELL_X2 FILLER_29_534 ();
 FILLCELL_X8 FILLER_30_1 ();
 FILLCELL_X4 FILLER_30_9 ();
 FILLCELL_X1 FILLER_30_13 ();
 FILLCELL_X16 FILLER_30_18 ();
 FILLCELL_X2 FILLER_30_34 ();
 FILLCELL_X4 FILLER_30_50 ();
 FILLCELL_X1 FILLER_30_54 ();
 FILLCELL_X8 FILLER_30_63 ();
 FILLCELL_X8 FILLER_30_81 ();
 FILLCELL_X2 FILLER_30_89 ();
 FILLCELL_X1 FILLER_30_91 ();
 FILLCELL_X4 FILLER_30_96 ();
 FILLCELL_X4 FILLER_30_105 ();
 FILLCELL_X1 FILLER_30_113 ();
 FILLCELL_X1 FILLER_30_118 ();
 FILLCELL_X1 FILLER_30_121 ();
 FILLCELL_X4 FILLER_30_126 ();
 FILLCELL_X1 FILLER_30_130 ();
 FILLCELL_X2 FILLER_30_135 ();
 FILLCELL_X1 FILLER_30_137 ();
 FILLCELL_X1 FILLER_30_141 ();
 FILLCELL_X8 FILLER_30_144 ();
 FILLCELL_X1 FILLER_30_152 ();
 FILLCELL_X8 FILLER_30_163 ();
 FILLCELL_X4 FILLER_30_171 ();
 FILLCELL_X2 FILLER_30_175 ();
 FILLCELL_X1 FILLER_30_177 ();
 FILLCELL_X1 FILLER_30_199 ();
 FILLCELL_X1 FILLER_30_213 ();
 FILLCELL_X8 FILLER_30_228 ();
 FILLCELL_X4 FILLER_30_236 ();
 FILLCELL_X4 FILLER_30_250 ();
 FILLCELL_X2 FILLER_30_254 ();
 FILLCELL_X1 FILLER_30_256 ();
 FILLCELL_X1 FILLER_30_277 ();
 FILLCELL_X16 FILLER_30_280 ();
 FILLCELL_X2 FILLER_30_318 ();
 FILLCELL_X8 FILLER_30_329 ();
 FILLCELL_X4 FILLER_30_337 ();
 FILLCELL_X4 FILLER_30_368 ();
 FILLCELL_X1 FILLER_30_382 ();
 FILLCELL_X8 FILLER_30_385 ();
 FILLCELL_X4 FILLER_30_393 ();
 FILLCELL_X2 FILLER_30_397 ();
 FILLCELL_X1 FILLER_30_399 ();
 FILLCELL_X2 FILLER_30_414 ();
 FILLCELL_X2 FILLER_30_426 ();
 FILLCELL_X1 FILLER_30_428 ();
 FILLCELL_X2 FILLER_30_444 ();
 FILLCELL_X1 FILLER_30_446 ();
 FILLCELL_X2 FILLER_30_478 ();
 FILLCELL_X8 FILLER_30_487 ();
 FILLCELL_X1 FILLER_30_495 ();
 FILLCELL_X2 FILLER_30_500 ();
 FILLCELL_X1 FILLER_30_502 ();
 FILLCELL_X4 FILLER_30_506 ();
 FILLCELL_X2 FILLER_30_510 ();
 FILLCELL_X1 FILLER_30_512 ();
 FILLCELL_X1 FILLER_30_525 ();
 FILLCELL_X1 FILLER_30_535 ();
 FILLCELL_X2 FILLER_31_1 ();
 FILLCELL_X1 FILLER_31_3 ();
 FILLCELL_X2 FILLER_31_13 ();
 FILLCELL_X1 FILLER_31_24 ();
 FILLCELL_X2 FILLER_31_34 ();
 FILLCELL_X1 FILLER_31_49 ();
 FILLCELL_X16 FILLER_31_56 ();
 FILLCELL_X2 FILLER_31_72 ();
 FILLCELL_X1 FILLER_31_74 ();
 FILLCELL_X2 FILLER_31_81 ();
 FILLCELL_X1 FILLER_31_85 ();
 FILLCELL_X2 FILLER_31_108 ();
 FILLCELL_X1 FILLER_31_120 ();
 FILLCELL_X2 FILLER_31_135 ();
 FILLCELL_X2 FILLER_31_145 ();
 FILLCELL_X1 FILLER_31_147 ();
 FILLCELL_X4 FILLER_31_155 ();
 FILLCELL_X1 FILLER_31_159 ();
 FILLCELL_X4 FILLER_31_164 ();
 FILLCELL_X1 FILLER_31_168 ();
 FILLCELL_X4 FILLER_31_181 ();
 FILLCELL_X4 FILLER_31_194 ();
 FILLCELL_X2 FILLER_31_198 ();
 FILLCELL_X4 FILLER_31_209 ();
 FILLCELL_X1 FILLER_31_213 ();
 FILLCELL_X1 FILLER_31_220 ();
 FILLCELL_X8 FILLER_31_231 ();
 FILLCELL_X1 FILLER_31_239 ();
 FILLCELL_X1 FILLER_31_249 ();
 FILLCELL_X4 FILLER_31_267 ();
 FILLCELL_X4 FILLER_31_284 ();
 FILLCELL_X1 FILLER_31_291 ();
 FILLCELL_X1 FILLER_31_294 ();
 FILLCELL_X1 FILLER_31_305 ();
 FILLCELL_X1 FILLER_31_310 ();
 FILLCELL_X2 FILLER_31_353 ();
 FILLCELL_X1 FILLER_31_355 ();
 FILLCELL_X8 FILLER_31_365 ();
 FILLCELL_X2 FILLER_31_373 ();
 FILLCELL_X1 FILLER_31_375 ();
 FILLCELL_X8 FILLER_31_382 ();
 FILLCELL_X4 FILLER_31_390 ();
 FILLCELL_X1 FILLER_31_394 ();
 FILLCELL_X2 FILLER_31_427 ();
 FILLCELL_X4 FILLER_31_457 ();
 FILLCELL_X4 FILLER_31_483 ();
 FILLCELL_X2 FILLER_31_487 ();
 FILLCELL_X8 FILLER_31_499 ();
 FILLCELL_X2 FILLER_31_507 ();
 FILLCELL_X1 FILLER_31_509 ();
 FILLCELL_X1 FILLER_31_520 ();
 FILLCELL_X4 FILLER_32_1 ();
 FILLCELL_X1 FILLER_32_19 ();
 FILLCELL_X4 FILLER_32_24 ();
 FILLCELL_X1 FILLER_32_28 ();
 FILLCELL_X2 FILLER_32_46 ();
 FILLCELL_X2 FILLER_32_53 ();
 FILLCELL_X2 FILLER_32_67 ();
 FILLCELL_X1 FILLER_32_80 ();
 FILLCELL_X4 FILLER_32_90 ();
 FILLCELL_X4 FILLER_32_112 ();
 FILLCELL_X2 FILLER_32_116 ();
 FILLCELL_X1 FILLER_32_118 ();
 FILLCELL_X1 FILLER_32_146 ();
 FILLCELL_X8 FILLER_32_149 ();
 FILLCELL_X4 FILLER_32_157 ();
 FILLCELL_X2 FILLER_32_161 ();
 FILLCELL_X1 FILLER_32_163 ();
 FILLCELL_X2 FILLER_32_168 ();
 FILLCELL_X1 FILLER_32_170 ();
 FILLCELL_X1 FILLER_32_175 ();
 FILLCELL_X8 FILLER_32_180 ();
 FILLCELL_X8 FILLER_32_199 ();
 FILLCELL_X2 FILLER_32_207 ();
 FILLCELL_X2 FILLER_32_219 ();
 FILLCELL_X1 FILLER_32_221 ();
 FILLCELL_X4 FILLER_32_239 ();
 FILLCELL_X2 FILLER_32_271 ();
 FILLCELL_X1 FILLER_32_273 ();
 FILLCELL_X8 FILLER_32_283 ();
 FILLCELL_X2 FILLER_32_291 ();
 FILLCELL_X2 FILLER_32_300 ();
 FILLCELL_X1 FILLER_32_302 ();
 FILLCELL_X8 FILLER_32_315 ();
 FILLCELL_X4 FILLER_32_323 ();
 FILLCELL_X2 FILLER_32_327 ();
 FILLCELL_X8 FILLER_32_333 ();
 FILLCELL_X2 FILLER_32_341 ();
 FILLCELL_X4 FILLER_32_351 ();
 FILLCELL_X1 FILLER_32_355 ();
 FILLCELL_X8 FILLER_32_367 ();
 FILLCELL_X8 FILLER_32_389 ();
 FILLCELL_X4 FILLER_32_397 ();
 FILLCELL_X16 FILLER_32_428 ();
 FILLCELL_X2 FILLER_32_444 ();
 FILLCELL_X1 FILLER_32_446 ();
 FILLCELL_X4 FILLER_32_506 ();
 FILLCELL_X1 FILLER_32_520 ();
 FILLCELL_X1 FILLER_32_523 ();
 FILLCELL_X4 FILLER_32_529 ();
 FILLCELL_X2 FILLER_32_533 ();
 FILLCELL_X1 FILLER_32_535 ();
 FILLCELL_X8 FILLER_33_1 ();
 FILLCELL_X4 FILLER_33_9 ();
 FILLCELL_X4 FILLER_33_25 ();
 FILLCELL_X4 FILLER_33_47 ();
 FILLCELL_X2 FILLER_33_61 ();
 FILLCELL_X2 FILLER_33_84 ();
 FILLCELL_X2 FILLER_33_95 ();
 FILLCELL_X1 FILLER_33_103 ();
 FILLCELL_X2 FILLER_33_114 ();
 FILLCELL_X1 FILLER_33_116 ();
 FILLCELL_X4 FILLER_33_127 ();
 FILLCELL_X4 FILLER_33_135 ();
 FILLCELL_X2 FILLER_33_157 ();
 FILLCELL_X16 FILLER_33_175 ();
 FILLCELL_X4 FILLER_33_191 ();
 FILLCELL_X1 FILLER_33_205 ();
 FILLCELL_X1 FILLER_33_219 ();
 FILLCELL_X1 FILLER_33_229 ();
 FILLCELL_X8 FILLER_33_232 ();
 FILLCELL_X8 FILLER_33_244 ();
 FILLCELL_X2 FILLER_33_252 ();
 FILLCELL_X1 FILLER_33_254 ();
 FILLCELL_X8 FILLER_33_268 ();
 FILLCELL_X4 FILLER_33_276 ();
 FILLCELL_X1 FILLER_33_290 ();
 FILLCELL_X8 FILLER_33_313 ();
 FILLCELL_X1 FILLER_33_376 ();
 FILLCELL_X4 FILLER_33_388 ();
 FILLCELL_X1 FILLER_33_392 ();
 FILLCELL_X2 FILLER_33_422 ();
 FILLCELL_X8 FILLER_33_437 ();
 FILLCELL_X4 FILLER_33_445 ();
 FILLCELL_X1 FILLER_33_449 ();
 FILLCELL_X8 FILLER_33_478 ();
 FILLCELL_X1 FILLER_33_486 ();
 FILLCELL_X4 FILLER_33_494 ();
 FILLCELL_X8 FILLER_33_524 ();
 FILLCELL_X4 FILLER_33_532 ();
 FILLCELL_X4 FILLER_34_1 ();
 FILLCELL_X1 FILLER_34_5 ();
 FILLCELL_X1 FILLER_34_49 ();
 FILLCELL_X1 FILLER_34_60 ();
 FILLCELL_X1 FILLER_34_71 ();
 FILLCELL_X4 FILLER_34_76 ();
 FILLCELL_X4 FILLER_34_84 ();
 FILLCELL_X2 FILLER_34_88 ();
 FILLCELL_X1 FILLER_34_90 ();
 FILLCELL_X8 FILLER_34_101 ();
 FILLCELL_X1 FILLER_34_109 ();
 FILLCELL_X8 FILLER_34_120 ();
 FILLCELL_X1 FILLER_34_128 ();
 FILLCELL_X8 FILLER_34_136 ();
 FILLCELL_X2 FILLER_34_144 ();
 FILLCELL_X8 FILLER_34_158 ();
 FILLCELL_X4 FILLER_34_179 ();
 FILLCELL_X2 FILLER_34_183 ();
 FILLCELL_X1 FILLER_34_185 ();
 FILLCELL_X8 FILLER_34_199 ();
 FILLCELL_X4 FILLER_34_207 ();
 FILLCELL_X2 FILLER_34_211 ();
 FILLCELL_X1 FILLER_34_213 ();
 FILLCELL_X4 FILLER_34_224 ();
 FILLCELL_X2 FILLER_34_228 ();
 FILLCELL_X1 FILLER_34_240 ();
 FILLCELL_X8 FILLER_34_256 ();
 FILLCELL_X4 FILLER_34_264 ();
 FILLCELL_X2 FILLER_34_268 ();
 FILLCELL_X4 FILLER_34_287 ();
 FILLCELL_X2 FILLER_34_291 ();
 FILLCELL_X1 FILLER_34_293 ();
 FILLCELL_X1 FILLER_34_298 ();
 FILLCELL_X32 FILLER_34_307 ();
 FILLCELL_X4 FILLER_34_339 ();
 FILLCELL_X8 FILLER_34_367 ();
 FILLCELL_X2 FILLER_34_375 ();
 FILLCELL_X1 FILLER_34_377 ();
 FILLCELL_X8 FILLER_34_388 ();
 FILLCELL_X2 FILLER_34_396 ();
 FILLCELL_X4 FILLER_34_413 ();
 FILLCELL_X1 FILLER_34_417 ();
 FILLCELL_X8 FILLER_34_424 ();
 FILLCELL_X4 FILLER_34_487 ();
 FILLCELL_X1 FILLER_34_507 ();
 FILLCELL_X8 FILLER_34_527 ();
 FILLCELL_X1 FILLER_34_535 ();
 FILLCELL_X2 FILLER_35_1 ();
 FILLCELL_X1 FILLER_35_3 ();
 FILLCELL_X8 FILLER_35_11 ();
 FILLCELL_X2 FILLER_35_19 ();
 FILLCELL_X2 FILLER_35_31 ();
 FILLCELL_X1 FILLER_35_33 ();
 FILLCELL_X1 FILLER_35_60 ();
 FILLCELL_X16 FILLER_35_69 ();
 FILLCELL_X2 FILLER_35_85 ();
 FILLCELL_X1 FILLER_35_87 ();
 FILLCELL_X8 FILLER_35_95 ();
 FILLCELL_X4 FILLER_35_103 ();
 FILLCELL_X1 FILLER_35_107 ();
 FILLCELL_X8 FILLER_35_116 ();
 FILLCELL_X2 FILLER_35_124 ();
 FILLCELL_X1 FILLER_35_126 ();
 FILLCELL_X4 FILLER_35_134 ();
 FILLCELL_X4 FILLER_35_155 ();
 FILLCELL_X2 FILLER_35_169 ();
 FILLCELL_X1 FILLER_35_171 ();
 FILLCELL_X8 FILLER_35_174 ();
 FILLCELL_X2 FILLER_35_182 ();
 FILLCELL_X1 FILLER_35_184 ();
 FILLCELL_X1 FILLER_35_187 ();
 FILLCELL_X1 FILLER_35_191 ();
 FILLCELL_X4 FILLER_35_202 ();
 FILLCELL_X2 FILLER_35_206 ();
 FILLCELL_X1 FILLER_35_208 ();
 FILLCELL_X4 FILLER_35_221 ();
 FILLCELL_X2 FILLER_35_225 ();
 FILLCELL_X1 FILLER_35_227 ();
 FILLCELL_X8 FILLER_35_231 ();
 FILLCELL_X1 FILLER_35_241 ();
 FILLCELL_X16 FILLER_35_254 ();
 FILLCELL_X4 FILLER_35_270 ();
 FILLCELL_X2 FILLER_35_274 ();
 FILLCELL_X1 FILLER_35_276 ();
 FILLCELL_X1 FILLER_35_287 ();
 FILLCELL_X8 FILLER_35_309 ();
 FILLCELL_X2 FILLER_35_317 ();
 FILLCELL_X1 FILLER_35_319 ();
 FILLCELL_X2 FILLER_35_326 ();
 FILLCELL_X8 FILLER_35_348 ();
 FILLCELL_X4 FILLER_35_356 ();
 FILLCELL_X2 FILLER_35_360 ();
 FILLCELL_X2 FILLER_35_396 ();
 FILLCELL_X4 FILLER_35_449 ();
 FILLCELL_X1 FILLER_35_453 ();
 FILLCELL_X8 FILLER_35_487 ();
 FILLCELL_X2 FILLER_35_495 ();
 FILLCELL_X1 FILLER_35_497 ();
 FILLCELL_X16 FILLER_35_518 ();
 FILLCELL_X2 FILLER_35_534 ();
 FILLCELL_X4 FILLER_36_1 ();
 FILLCELL_X2 FILLER_36_5 ();
 FILLCELL_X1 FILLER_36_21 ();
 FILLCELL_X4 FILLER_36_47 ();
 FILLCELL_X2 FILLER_36_60 ();
 FILLCELL_X1 FILLER_36_62 ();
 FILLCELL_X1 FILLER_36_81 ();
 FILLCELL_X1 FILLER_36_102 ();
 FILLCELL_X2 FILLER_36_110 ();
 FILLCELL_X4 FILLER_36_124 ();
 FILLCELL_X2 FILLER_36_128 ();
 FILLCELL_X2 FILLER_36_137 ();
 FILLCELL_X4 FILLER_36_141 ();
 FILLCELL_X1 FILLER_36_145 ();
 FILLCELL_X8 FILLER_36_150 ();
 FILLCELL_X2 FILLER_36_158 ();
 FILLCELL_X1 FILLER_36_160 ();
 FILLCELL_X1 FILLER_36_170 ();
 FILLCELL_X4 FILLER_36_181 ();
 FILLCELL_X2 FILLER_36_203 ();
 FILLCELL_X4 FILLER_36_208 ();
 FILLCELL_X1 FILLER_36_212 ();
 FILLCELL_X8 FILLER_36_219 ();
 FILLCELL_X1 FILLER_36_241 ();
 FILLCELL_X2 FILLER_36_266 ();
 FILLCELL_X1 FILLER_36_268 ();
 FILLCELL_X2 FILLER_36_316 ();
 FILLCELL_X2 FILLER_36_323 ();
 FILLCELL_X1 FILLER_36_325 ();
 FILLCELL_X16 FILLER_36_328 ();
 FILLCELL_X2 FILLER_36_344 ();
 FILLCELL_X1 FILLER_36_346 ();
 FILLCELL_X4 FILLER_36_365 ();
 FILLCELL_X2 FILLER_36_371 ();
 FILLCELL_X2 FILLER_36_389 ();
 FILLCELL_X1 FILLER_36_391 ();
 FILLCELL_X4 FILLER_36_411 ();
 FILLCELL_X2 FILLER_36_415 ();
 FILLCELL_X1 FILLER_36_417 ();
 FILLCELL_X4 FILLER_36_445 ();
 FILLCELL_X2 FILLER_36_449 ();
 FILLCELL_X2 FILLER_36_455 ();
 FILLCELL_X1 FILLER_36_481 ();
 FILLCELL_X2 FILLER_36_488 ();
 FILLCELL_X8 FILLER_36_522 ();
 FILLCELL_X4 FILLER_36_530 ();
 FILLCELL_X2 FILLER_36_534 ();
 FILLCELL_X8 FILLER_37_1 ();
 FILLCELL_X4 FILLER_37_9 ();
 FILLCELL_X2 FILLER_37_16 ();
 FILLCELL_X1 FILLER_37_22 ();
 FILLCELL_X1 FILLER_37_27 ();
 FILLCELL_X2 FILLER_37_43 ();
 FILLCELL_X1 FILLER_37_55 ();
 FILLCELL_X2 FILLER_37_62 ();
 FILLCELL_X8 FILLER_37_71 ();
 FILLCELL_X1 FILLER_37_79 ();
 FILLCELL_X2 FILLER_37_91 ();
 FILLCELL_X4 FILLER_37_95 ();
 FILLCELL_X1 FILLER_37_99 ();
 FILLCELL_X2 FILLER_37_102 ();
 FILLCELL_X4 FILLER_37_111 ();
 FILLCELL_X1 FILLER_37_115 ();
 FILLCELL_X4 FILLER_37_120 ();
 FILLCELL_X1 FILLER_37_151 ();
 FILLCELL_X2 FILLER_37_154 ();
 FILLCELL_X8 FILLER_37_174 ();
 FILLCELL_X8 FILLER_37_217 ();
 FILLCELL_X2 FILLER_37_225 ();
 FILLCELL_X1 FILLER_37_239 ();
 FILLCELL_X1 FILLER_37_242 ();
 FILLCELL_X4 FILLER_37_250 ();
 FILLCELL_X1 FILLER_37_254 ();
 FILLCELL_X4 FILLER_37_261 ();
 FILLCELL_X2 FILLER_37_265 ();
 FILLCELL_X1 FILLER_37_279 ();
 FILLCELL_X1 FILLER_37_299 ();
 FILLCELL_X2 FILLER_37_306 ();
 FILLCELL_X8 FILLER_37_357 ();
 FILLCELL_X4 FILLER_37_365 ();
 FILLCELL_X2 FILLER_37_392 ();
 FILLCELL_X1 FILLER_37_394 ();
 FILLCELL_X4 FILLER_37_404 ();
 FILLCELL_X1 FILLER_37_408 ();
 FILLCELL_X4 FILLER_37_426 ();
 FILLCELL_X2 FILLER_37_430 ();
 FILLCELL_X1 FILLER_37_432 ();
 FILLCELL_X4 FILLER_37_443 ();
 FILLCELL_X1 FILLER_37_460 ();
 FILLCELL_X1 FILLER_37_473 ();
 FILLCELL_X4 FILLER_37_488 ();
 FILLCELL_X1 FILLER_37_492 ();
 FILLCELL_X1 FILLER_37_505 ();
 FILLCELL_X4 FILLER_37_532 ();
 FILLCELL_X2 FILLER_38_1 ();
 FILLCELL_X1 FILLER_38_16 ();
 FILLCELL_X8 FILLER_38_35 ();
 FILLCELL_X1 FILLER_38_43 ();
 FILLCELL_X4 FILLER_38_52 ();
 FILLCELL_X1 FILLER_38_56 ();
 FILLCELL_X8 FILLER_38_76 ();
 FILLCELL_X4 FILLER_38_84 ();
 FILLCELL_X2 FILLER_38_88 ();
 FILLCELL_X4 FILLER_38_110 ();
 FILLCELL_X2 FILLER_38_121 ();
 FILLCELL_X2 FILLER_38_125 ();
 FILLCELL_X16 FILLER_38_161 ();
 FILLCELL_X8 FILLER_38_177 ();
 FILLCELL_X2 FILLER_38_189 ();
 FILLCELL_X16 FILLER_38_195 ();
 FILLCELL_X4 FILLER_38_211 ();
 FILLCELL_X2 FILLER_38_215 ();
 FILLCELL_X4 FILLER_38_227 ();
 FILLCELL_X2 FILLER_38_231 ();
 FILLCELL_X1 FILLER_38_233 ();
 FILLCELL_X1 FILLER_38_238 ();
 FILLCELL_X8 FILLER_38_256 ();
 FILLCELL_X4 FILLER_38_264 ();
 FILLCELL_X2 FILLER_38_268 ();
 FILLCELL_X2 FILLER_38_280 ();
 FILLCELL_X1 FILLER_38_286 ();
 FILLCELL_X32 FILLER_38_291 ();
 FILLCELL_X1 FILLER_38_323 ();
 FILLCELL_X8 FILLER_38_337 ();
 FILLCELL_X1 FILLER_38_368 ();
 FILLCELL_X2 FILLER_38_385 ();
 FILLCELL_X1 FILLER_38_387 ();
 FILLCELL_X2 FILLER_38_401 ();
 FILLCELL_X1 FILLER_38_403 ();
 FILLCELL_X1 FILLER_38_430 ();
 FILLCELL_X2 FILLER_38_433 ();
 FILLCELL_X4 FILLER_38_451 ();
 FILLCELL_X1 FILLER_38_455 ();
 FILLCELL_X8 FILLER_38_459 ();
 FILLCELL_X1 FILLER_38_467 ();
 FILLCELL_X1 FILLER_38_474 ();
 FILLCELL_X16 FILLER_38_484 ();
 FILLCELL_X1 FILLER_38_535 ();
 FILLCELL_X8 FILLER_39_1 ();
 FILLCELL_X2 FILLER_39_9 ();
 FILLCELL_X1 FILLER_39_20 ();
 FILLCELL_X1 FILLER_39_31 ();
 FILLCELL_X1 FILLER_39_36 ();
 FILLCELL_X1 FILLER_39_67 ();
 FILLCELL_X16 FILLER_39_78 ();
 FILLCELL_X4 FILLER_39_94 ();
 FILLCELL_X2 FILLER_39_98 ();
 FILLCELL_X1 FILLER_39_100 ();
 FILLCELL_X2 FILLER_39_111 ();
 FILLCELL_X1 FILLER_39_123 ();
 FILLCELL_X2 FILLER_39_148 ();
 FILLCELL_X8 FILLER_39_152 ();
 FILLCELL_X4 FILLER_39_160 ();
 FILLCELL_X2 FILLER_39_164 ();
 FILLCELL_X1 FILLER_39_166 ();
 FILLCELL_X4 FILLER_39_177 ();
 FILLCELL_X1 FILLER_39_181 ();
 FILLCELL_X8 FILLER_39_205 ();
 FILLCELL_X4 FILLER_39_213 ();
 FILLCELL_X2 FILLER_39_217 ();
 FILLCELL_X2 FILLER_39_236 ();
 FILLCELL_X16 FILLER_39_249 ();
 FILLCELL_X4 FILLER_39_265 ();
 FILLCELL_X2 FILLER_39_269 ();
 FILLCELL_X1 FILLER_39_271 ();
 FILLCELL_X1 FILLER_39_278 ();
 FILLCELL_X8 FILLER_39_298 ();
 FILLCELL_X4 FILLER_39_312 ();
 FILLCELL_X2 FILLER_39_316 ();
 FILLCELL_X2 FILLER_39_347 ();
 FILLCELL_X1 FILLER_39_367 ();
 FILLCELL_X1 FILLER_39_377 ();
 FILLCELL_X2 FILLER_39_404 ();
 FILLCELL_X1 FILLER_39_416 ();
 FILLCELL_X1 FILLER_39_462 ();
 FILLCELL_X1 FILLER_39_465 ();
 FILLCELL_X8 FILLER_39_479 ();
 FILLCELL_X2 FILLER_39_487 ();
 FILLCELL_X1 FILLER_39_489 ();
 FILLCELL_X8 FILLER_39_515 ();
 FILLCELL_X1 FILLER_39_523 ();
 FILLCELL_X2 FILLER_39_534 ();
 FILLCELL_X16 FILLER_40_1 ();
 FILLCELL_X4 FILLER_40_17 ();
 FILLCELL_X2 FILLER_40_21 ();
 FILLCELL_X1 FILLER_40_23 ();
 FILLCELL_X4 FILLER_40_34 ();
 FILLCELL_X1 FILLER_40_38 ();
 FILLCELL_X4 FILLER_40_49 ();
 FILLCELL_X1 FILLER_40_57 ();
 FILLCELL_X2 FILLER_40_62 ();
 FILLCELL_X1 FILLER_40_64 ();
 FILLCELL_X1 FILLER_40_75 ();
 FILLCELL_X4 FILLER_40_92 ();
 FILLCELL_X2 FILLER_40_96 ();
 FILLCELL_X4 FILLER_40_101 ();
 FILLCELL_X1 FILLER_40_112 ();
 FILLCELL_X16 FILLER_40_116 ();
 FILLCELL_X1 FILLER_40_132 ();
 FILLCELL_X4 FILLER_40_135 ();
 FILLCELL_X2 FILLER_40_139 ();
 FILLCELL_X4 FILLER_40_162 ();
 FILLCELL_X4 FILLER_40_180 ();
 FILLCELL_X4 FILLER_40_190 ();
 FILLCELL_X8 FILLER_40_207 ();
 FILLCELL_X1 FILLER_40_215 ();
 FILLCELL_X1 FILLER_40_243 ();
 FILLCELL_X4 FILLER_40_250 ();
 FILLCELL_X2 FILLER_40_254 ();
 FILLCELL_X2 FILLER_40_266 ();
 FILLCELL_X1 FILLER_40_289 ();
 FILLCELL_X2 FILLER_40_300 ();
 FILLCELL_X1 FILLER_40_306 ();
 FILLCELL_X4 FILLER_40_327 ();
 FILLCELL_X2 FILLER_40_331 ();
 FILLCELL_X1 FILLER_40_371 ();
 FILLCELL_X4 FILLER_40_400 ();
 FILLCELL_X2 FILLER_40_404 ();
 FILLCELL_X1 FILLER_40_406 ();
 FILLCELL_X8 FILLER_40_412 ();
 FILLCELL_X4 FILLER_40_420 ();
 FILLCELL_X2 FILLER_40_460 ();
 FILLCELL_X16 FILLER_40_474 ();
 FILLCELL_X8 FILLER_40_501 ();
 FILLCELL_X2 FILLER_40_509 ();
 FILLCELL_X1 FILLER_40_511 ();
 FILLCELL_X1 FILLER_40_522 ();
 FILLCELL_X2 FILLER_40_533 ();
 FILLCELL_X1 FILLER_40_535 ();
 FILLCELL_X16 FILLER_41_1 ();
 FILLCELL_X2 FILLER_41_17 ();
 FILLCELL_X8 FILLER_41_32 ();
 FILLCELL_X8 FILLER_41_59 ();
 FILLCELL_X4 FILLER_41_67 ();
 FILLCELL_X2 FILLER_41_71 ();
 FILLCELL_X1 FILLER_41_73 ();
 FILLCELL_X2 FILLER_41_76 ();
 FILLCELL_X1 FILLER_41_78 ();
 FILLCELL_X1 FILLER_41_84 ();
 FILLCELL_X1 FILLER_41_102 ();
 FILLCELL_X4 FILLER_41_118 ();
 FILLCELL_X1 FILLER_41_122 ();
 FILLCELL_X2 FILLER_41_152 ();
 FILLCELL_X8 FILLER_41_156 ();
 FILLCELL_X2 FILLER_41_180 ();
 FILLCELL_X8 FILLER_41_196 ();
 FILLCELL_X4 FILLER_41_204 ();
 FILLCELL_X2 FILLER_41_208 ();
 FILLCELL_X1 FILLER_41_210 ();
 FILLCELL_X4 FILLER_41_246 ();
 FILLCELL_X2 FILLER_41_250 ();
 FILLCELL_X8 FILLER_41_262 ();
 FILLCELL_X4 FILLER_41_270 ();
 FILLCELL_X8 FILLER_41_280 ();
 FILLCELL_X4 FILLER_41_288 ();
 FILLCELL_X2 FILLER_41_292 ();
 FILLCELL_X1 FILLER_41_294 ();
 FILLCELL_X2 FILLER_41_304 ();
 FILLCELL_X1 FILLER_41_306 ();
 FILLCELL_X2 FILLER_41_339 ();
 FILLCELL_X1 FILLER_41_341 ();
 FILLCELL_X4 FILLER_41_352 ();
 FILLCELL_X2 FILLER_41_356 ();
 FILLCELL_X1 FILLER_41_358 ();
 FILLCELL_X2 FILLER_41_378 ();
 FILLCELL_X2 FILLER_41_409 ();
 FILLCELL_X4 FILLER_41_431 ();
 FILLCELL_X1 FILLER_41_435 ();
 FILLCELL_X4 FILLER_41_452 ();
 FILLCELL_X16 FILLER_41_475 ();
 FILLCELL_X2 FILLER_41_491 ();
 FILLCELL_X1 FILLER_41_493 ();
 FILLCELL_X16 FILLER_41_500 ();
 FILLCELL_X2 FILLER_41_516 ();
 FILLCELL_X1 FILLER_41_518 ();
 FILLCELL_X2 FILLER_42_29 ();
 FILLCELL_X2 FILLER_42_43 ();
 FILLCELL_X1 FILLER_42_45 ();
 FILLCELL_X1 FILLER_42_59 ();
 FILLCELL_X8 FILLER_42_63 ();
 FILLCELL_X1 FILLER_42_71 ();
 FILLCELL_X1 FILLER_42_77 ();
 FILLCELL_X2 FILLER_42_95 ();
 FILLCELL_X1 FILLER_42_97 ();
 FILLCELL_X4 FILLER_42_106 ();
 FILLCELL_X2 FILLER_42_110 ();
 FILLCELL_X8 FILLER_42_122 ();
 FILLCELL_X2 FILLER_42_130 ();
 FILLCELL_X1 FILLER_42_139 ();
 FILLCELL_X1 FILLER_42_143 ();
 FILLCELL_X1 FILLER_42_147 ();
 FILLCELL_X1 FILLER_42_154 ();
 FILLCELL_X1 FILLER_42_167 ();
 FILLCELL_X8 FILLER_42_178 ();
 FILLCELL_X2 FILLER_42_186 ();
 FILLCELL_X1 FILLER_42_188 ();
 FILLCELL_X1 FILLER_42_224 ();
 FILLCELL_X8 FILLER_42_241 ();
 FILLCELL_X2 FILLER_42_303 ();
 FILLCELL_X1 FILLER_42_305 ();
 FILLCELL_X4 FILLER_42_308 ();
 FILLCELL_X1 FILLER_42_312 ();
 FILLCELL_X4 FILLER_42_325 ();
 FILLCELL_X2 FILLER_42_329 ();
 FILLCELL_X1 FILLER_42_331 ();
 FILLCELL_X4 FILLER_42_341 ();
 FILLCELL_X2 FILLER_42_345 ();
 FILLCELL_X2 FILLER_42_357 ();
 FILLCELL_X16 FILLER_42_362 ();
 FILLCELL_X1 FILLER_42_385 ();
 FILLCELL_X2 FILLER_42_396 ();
 FILLCELL_X1 FILLER_42_398 ();
 FILLCELL_X8 FILLER_42_409 ();
 FILLCELL_X1 FILLER_42_417 ();
 FILLCELL_X2 FILLER_42_420 ();
 FILLCELL_X2 FILLER_42_429 ();
 FILLCELL_X2 FILLER_42_444 ();
 FILLCELL_X4 FILLER_42_461 ();
 FILLCELL_X2 FILLER_42_490 ();
 FILLCELL_X1 FILLER_42_492 ();
 FILLCELL_X2 FILLER_42_496 ();
 FILLCELL_X2 FILLER_42_504 ();
 FILLCELL_X4 FILLER_42_531 ();
 FILLCELL_X1 FILLER_42_535 ();
 FILLCELL_X16 FILLER_43_1 ();
 FILLCELL_X2 FILLER_43_17 ();
 FILLCELL_X2 FILLER_43_55 ();
 FILLCELL_X2 FILLER_43_66 ();
 FILLCELL_X4 FILLER_43_127 ();
 FILLCELL_X1 FILLER_43_131 ();
 FILLCELL_X4 FILLER_43_157 ();
 FILLCELL_X32 FILLER_43_170 ();
 FILLCELL_X8 FILLER_43_202 ();
 FILLCELL_X4 FILLER_43_210 ();
 FILLCELL_X2 FILLER_43_214 ();
 FILLCELL_X1 FILLER_43_216 ();
 FILLCELL_X8 FILLER_43_244 ();
 FILLCELL_X4 FILLER_43_252 ();
 FILLCELL_X1 FILLER_43_262 ();
 FILLCELL_X16 FILLER_43_309 ();
 FILLCELL_X8 FILLER_43_325 ();
 FILLCELL_X2 FILLER_43_333 ();
 FILLCELL_X1 FILLER_43_335 ();
 FILLCELL_X8 FILLER_43_352 ();
 FILLCELL_X8 FILLER_43_372 ();
 FILLCELL_X2 FILLER_43_380 ();
 FILLCELL_X1 FILLER_43_382 ();
 FILLCELL_X4 FILLER_43_398 ();
 FILLCELL_X1 FILLER_43_402 ();
 FILLCELL_X4 FILLER_43_421 ();
 FILLCELL_X2 FILLER_43_425 ();
 FILLCELL_X1 FILLER_43_427 ();
 FILLCELL_X1 FILLER_43_432 ();
 FILLCELL_X16 FILLER_43_443 ();
 FILLCELL_X1 FILLER_43_459 ();
 FILLCELL_X16 FILLER_43_463 ();
 FILLCELL_X4 FILLER_43_479 ();
 FILLCELL_X2 FILLER_43_496 ();
 FILLCELL_X2 FILLER_43_520 ();
 FILLCELL_X1 FILLER_43_524 ();
 FILLCELL_X8 FILLER_43_527 ();
 FILLCELL_X1 FILLER_43_535 ();
 FILLCELL_X8 FILLER_44_1 ();
 FILLCELL_X4 FILLER_44_9 ();
 FILLCELL_X2 FILLER_44_13 ();
 FILLCELL_X4 FILLER_44_41 ();
 FILLCELL_X2 FILLER_44_45 ();
 FILLCELL_X4 FILLER_44_61 ();
 FILLCELL_X2 FILLER_44_65 ();
 FILLCELL_X1 FILLER_44_67 ();
 FILLCELL_X2 FILLER_44_73 ();
 FILLCELL_X4 FILLER_44_84 ();
 FILLCELL_X2 FILLER_44_92 ();
 FILLCELL_X1 FILLER_44_97 ();
 FILLCELL_X1 FILLER_44_100 ();
 FILLCELL_X1 FILLER_44_111 ();
 FILLCELL_X2 FILLER_44_128 ();
 FILLCELL_X1 FILLER_44_130 ();
 FILLCELL_X16 FILLER_44_133 ();
 FILLCELL_X8 FILLER_44_149 ();
 FILLCELL_X4 FILLER_44_170 ();
 FILLCELL_X16 FILLER_44_176 ();
 FILLCELL_X8 FILLER_44_192 ();
 FILLCELL_X4 FILLER_44_200 ();
 FILLCELL_X2 FILLER_44_204 ();
 FILLCELL_X1 FILLER_44_206 ();
 FILLCELL_X4 FILLER_44_220 ();
 FILLCELL_X2 FILLER_44_224 ();
 FILLCELL_X1 FILLER_44_226 ();
 FILLCELL_X1 FILLER_44_235 ();
 FILLCELL_X1 FILLER_44_242 ();
 FILLCELL_X2 FILLER_44_253 ();
 FILLCELL_X16 FILLER_44_263 ();
 FILLCELL_X4 FILLER_44_279 ();
 FILLCELL_X2 FILLER_44_283 ();
 FILLCELL_X4 FILLER_44_287 ();
 FILLCELL_X1 FILLER_44_291 ();
 FILLCELL_X8 FILLER_44_320 ();
 FILLCELL_X2 FILLER_44_328 ();
 FILLCELL_X1 FILLER_44_330 ();
 FILLCELL_X8 FILLER_44_340 ();
 FILLCELL_X4 FILLER_44_348 ();
 FILLCELL_X2 FILLER_44_352 ();
 FILLCELL_X1 FILLER_44_354 ();
 FILLCELL_X4 FILLER_44_357 ();
 FILLCELL_X1 FILLER_44_361 ();
 FILLCELL_X2 FILLER_44_378 ();
 FILLCELL_X1 FILLER_44_392 ();
 FILLCELL_X4 FILLER_44_406 ();
 FILLCELL_X4 FILLER_44_421 ();
 FILLCELL_X1 FILLER_44_425 ();
 FILLCELL_X4 FILLER_44_432 ();
 FILLCELL_X2 FILLER_44_436 ();
 FILLCELL_X1 FILLER_44_453 ();
 FILLCELL_X1 FILLER_44_483 ();
 FILLCELL_X8 FILLER_44_501 ();
 FILLCELL_X4 FILLER_44_509 ();
 FILLCELL_X2 FILLER_44_513 ();
 FILLCELL_X1 FILLER_44_515 ();
 FILLCELL_X4 FILLER_44_519 ();
 FILLCELL_X16 FILLER_45_1 ();
 FILLCELL_X2 FILLER_45_17 ();
 FILLCELL_X1 FILLER_45_26 ();
 FILLCELL_X1 FILLER_45_36 ();
 FILLCELL_X4 FILLER_45_41 ();
 FILLCELL_X2 FILLER_45_45 ();
 FILLCELL_X1 FILLER_45_47 ();
 FILLCELL_X2 FILLER_45_64 ();
 FILLCELL_X1 FILLER_45_66 ();
 FILLCELL_X2 FILLER_45_86 ();
 FILLCELL_X4 FILLER_45_109 ();
 FILLCELL_X1 FILLER_45_113 ();
 FILLCELL_X1 FILLER_45_118 ();
 FILLCELL_X1 FILLER_45_126 ();
 FILLCELL_X4 FILLER_45_134 ();
 FILLCELL_X1 FILLER_45_138 ();
 FILLCELL_X8 FILLER_45_159 ();
 FILLCELL_X4 FILLER_45_194 ();
 FILLCELL_X2 FILLER_45_198 ();
 FILLCELL_X1 FILLER_45_210 ();
 FILLCELL_X2 FILLER_45_224 ();
 FILLCELL_X1 FILLER_45_226 ();
 FILLCELL_X16 FILLER_45_239 ();
 FILLCELL_X2 FILLER_45_255 ();
 FILLCELL_X4 FILLER_45_276 ();
 FILLCELL_X2 FILLER_45_290 ();
 FILLCELL_X2 FILLER_45_296 ();
 FILLCELL_X1 FILLER_45_331 ();
 FILLCELL_X4 FILLER_45_345 ();
 FILLCELL_X2 FILLER_45_349 ();
 FILLCELL_X8 FILLER_45_360 ();
 FILLCELL_X2 FILLER_45_368 ();
 FILLCELL_X1 FILLER_45_370 ();
 FILLCELL_X16 FILLER_45_373 ();
 FILLCELL_X2 FILLER_45_389 ();
 FILLCELL_X8 FILLER_45_398 ();
 FILLCELL_X2 FILLER_45_406 ();
 FILLCELL_X1 FILLER_45_408 ();
 FILLCELL_X4 FILLER_45_426 ();
 FILLCELL_X2 FILLER_45_430 ();
 FILLCELL_X1 FILLER_45_432 ();
 FILLCELL_X4 FILLER_45_459 ();
 FILLCELL_X1 FILLER_45_463 ();
 FILLCELL_X4 FILLER_45_494 ();
 FILLCELL_X2 FILLER_45_508 ();
 FILLCELL_X8 FILLER_45_526 ();
 FILLCELL_X2 FILLER_45_534 ();
 FILLCELL_X8 FILLER_46_1 ();
 FILLCELL_X2 FILLER_46_9 ();
 FILLCELL_X1 FILLER_46_11 ();
 FILLCELL_X1 FILLER_46_14 ();
 FILLCELL_X4 FILLER_46_23 ();
 FILLCELL_X16 FILLER_46_29 ();
 FILLCELL_X4 FILLER_46_71 ();
 FILLCELL_X2 FILLER_46_75 ();
 FILLCELL_X8 FILLER_46_81 ();
 FILLCELL_X1 FILLER_46_105 ();
 FILLCELL_X1 FILLER_46_108 ();
 FILLCELL_X4 FILLER_46_113 ();
 FILLCELL_X1 FILLER_46_117 ();
 FILLCELL_X1 FILLER_46_135 ();
 FILLCELL_X4 FILLER_46_146 ();
 FILLCELL_X1 FILLER_46_150 ();
 FILLCELL_X2 FILLER_46_162 ();
 FILLCELL_X1 FILLER_46_164 ();
 FILLCELL_X16 FILLER_46_177 ();
 FILLCELL_X1 FILLER_46_193 ();
 FILLCELL_X2 FILLER_46_204 ();
 FILLCELL_X1 FILLER_46_206 ();
 FILLCELL_X4 FILLER_46_217 ();
 FILLCELL_X2 FILLER_46_221 ();
 FILLCELL_X1 FILLER_46_223 ();
 FILLCELL_X1 FILLER_46_232 ();
 FILLCELL_X4 FILLER_46_238 ();
 FILLCELL_X2 FILLER_46_242 ();
 FILLCELL_X1 FILLER_46_244 ();
 FILLCELL_X1 FILLER_46_255 ();
 FILLCELL_X1 FILLER_46_283 ();
 FILLCELL_X4 FILLER_46_290 ();
 FILLCELL_X2 FILLER_46_304 ();
 FILLCELL_X1 FILLER_46_306 ();
 FILLCELL_X4 FILLER_46_319 ();
 FILLCELL_X1 FILLER_46_323 ();
 FILLCELL_X4 FILLER_46_328 ();
 FILLCELL_X1 FILLER_46_337 ();
 FILLCELL_X1 FILLER_46_364 ();
 FILLCELL_X8 FILLER_46_396 ();
 FILLCELL_X16 FILLER_46_424 ();
 FILLCELL_X8 FILLER_46_440 ();
 FILLCELL_X1 FILLER_46_448 ();
 FILLCELL_X2 FILLER_46_458 ();
 FILLCELL_X1 FILLER_46_460 ();
 FILLCELL_X1 FILLER_46_486 ();
 FILLCELL_X2 FILLER_46_500 ();
 FILLCELL_X1 FILLER_46_502 ();
 FILLCELL_X1 FILLER_46_509 ();
 FILLCELL_X4 FILLER_46_512 ();
 FILLCELL_X2 FILLER_46_533 ();
 FILLCELL_X1 FILLER_46_535 ();
 FILLCELL_X2 FILLER_47_1 ();
 FILLCELL_X1 FILLER_47_3 ();
 FILLCELL_X1 FILLER_47_37 ();
 FILLCELL_X4 FILLER_47_42 ();
 FILLCELL_X2 FILLER_47_50 ();
 FILLCELL_X4 FILLER_47_56 ();
 FILLCELL_X1 FILLER_47_60 ();
 FILLCELL_X8 FILLER_47_75 ();
 FILLCELL_X2 FILLER_47_83 ();
 FILLCELL_X1 FILLER_47_85 ();
 FILLCELL_X4 FILLER_47_116 ();
 FILLCELL_X1 FILLER_47_120 ();
 FILLCELL_X4 FILLER_47_131 ();
 FILLCELL_X1 FILLER_47_135 ();
 FILLCELL_X8 FILLER_47_140 ();
 FILLCELL_X2 FILLER_47_148 ();
 FILLCELL_X1 FILLER_47_161 ();
 FILLCELL_X4 FILLER_47_184 ();
 FILLCELL_X4 FILLER_47_200 ();
 FILLCELL_X1 FILLER_47_204 ();
 FILLCELL_X1 FILLER_47_212 ();
 FILLCELL_X2 FILLER_47_218 ();
 FILLCELL_X1 FILLER_47_220 ();
 FILLCELL_X2 FILLER_47_227 ();
 FILLCELL_X1 FILLER_47_234 ();
 FILLCELL_X4 FILLER_47_239 ();
 FILLCELL_X2 FILLER_47_243 ();
 FILLCELL_X1 FILLER_47_245 ();
 FILLCELL_X1 FILLER_47_256 ();
 FILLCELL_X2 FILLER_47_262 ();
 FILLCELL_X1 FILLER_47_264 ();
 FILLCELL_X1 FILLER_47_271 ();
 FILLCELL_X1 FILLER_47_295 ();
 FILLCELL_X2 FILLER_47_301 ();
 FILLCELL_X1 FILLER_47_303 ();
 FILLCELL_X2 FILLER_47_313 ();
 FILLCELL_X4 FILLER_47_335 ();
 FILLCELL_X1 FILLER_47_339 ();
 FILLCELL_X8 FILLER_47_352 ();
 FILLCELL_X1 FILLER_47_360 ();
 FILLCELL_X1 FILLER_47_389 ();
 FILLCELL_X1 FILLER_47_406 ();
 FILLCELL_X1 FILLER_47_423 ();
 FILLCELL_X1 FILLER_47_437 ();
 FILLCELL_X1 FILLER_47_440 ();
 FILLCELL_X4 FILLER_47_462 ();
 FILLCELL_X2 FILLER_47_466 ();
 FILLCELL_X1 FILLER_47_468 ();
 FILLCELL_X8 FILLER_47_490 ();
 FILLCELL_X2 FILLER_47_498 ();
 FILLCELL_X1 FILLER_47_533 ();
 FILLCELL_X4 FILLER_48_1 ();
 FILLCELL_X2 FILLER_48_5 ();
 FILLCELL_X1 FILLER_48_7 ();
 FILLCELL_X2 FILLER_48_17 ();
 FILLCELL_X1 FILLER_48_29 ();
 FILLCELL_X1 FILLER_48_32 ();
 FILLCELL_X4 FILLER_48_36 ();
 FILLCELL_X4 FILLER_48_65 ();
 FILLCELL_X1 FILLER_48_88 ();
 FILLCELL_X4 FILLER_48_126 ();
 FILLCELL_X1 FILLER_48_130 ();
 FILLCELL_X4 FILLER_48_143 ();
 FILLCELL_X2 FILLER_48_147 ();
 FILLCELL_X16 FILLER_48_159 ();
 FILLCELL_X8 FILLER_48_175 ();
 FILLCELL_X2 FILLER_48_183 ();
 FILLCELL_X1 FILLER_48_185 ();
 FILLCELL_X2 FILLER_48_188 ();
 FILLCELL_X2 FILLER_48_193 ();
 FILLCELL_X1 FILLER_48_195 ();
 FILLCELL_X2 FILLER_48_220 ();
 FILLCELL_X16 FILLER_48_232 ();
 FILLCELL_X4 FILLER_48_248 ();
 FILLCELL_X2 FILLER_48_252 ();
 FILLCELL_X1 FILLER_48_254 ();
 FILLCELL_X2 FILLER_48_257 ();
 FILLCELL_X1 FILLER_48_259 ();
 FILLCELL_X1 FILLER_48_263 ();
 FILLCELL_X1 FILLER_48_291 ();
 FILLCELL_X32 FILLER_48_319 ();
 FILLCELL_X4 FILLER_48_351 ();
 FILLCELL_X2 FILLER_48_355 ();
 FILLCELL_X8 FILLER_48_359 ();
 FILLCELL_X2 FILLER_48_367 ();
 FILLCELL_X1 FILLER_48_369 ();
 FILLCELL_X2 FILLER_48_384 ();
 FILLCELL_X2 FILLER_48_403 ();
 FILLCELL_X8 FILLER_48_469 ();
 FILLCELL_X1 FILLER_48_497 ();
 FILLCELL_X8 FILLER_48_508 ();
 FILLCELL_X2 FILLER_48_516 ();
 FILLCELL_X1 FILLER_48_535 ();
 FILLCELL_X8 FILLER_49_1 ();
 FILLCELL_X2 FILLER_49_9 ();
 FILLCELL_X1 FILLER_49_11 ();
 FILLCELL_X4 FILLER_49_25 ();
 FILLCELL_X2 FILLER_49_29 ();
 FILLCELL_X1 FILLER_49_37 ();
 FILLCELL_X2 FILLER_49_58 ();
 FILLCELL_X1 FILLER_49_60 ();
 FILLCELL_X8 FILLER_49_64 ();
 FILLCELL_X4 FILLER_49_72 ();
 FILLCELL_X1 FILLER_49_76 ();
 FILLCELL_X2 FILLER_49_105 ();
 FILLCELL_X2 FILLER_49_117 ();
 FILLCELL_X2 FILLER_49_124 ();
 FILLCELL_X1 FILLER_49_126 ();
 FILLCELL_X2 FILLER_49_134 ();
 FILLCELL_X1 FILLER_49_136 ();
 FILLCELL_X2 FILLER_49_150 ();
 FILLCELL_X1 FILLER_49_152 ();
 FILLCELL_X4 FILLER_49_163 ();
 FILLCELL_X2 FILLER_49_167 ();
 FILLCELL_X1 FILLER_49_200 ();
 FILLCELL_X32 FILLER_49_211 ();
 FILLCELL_X1 FILLER_49_243 ();
 FILLCELL_X8 FILLER_49_297 ();
 FILLCELL_X4 FILLER_49_305 ();
 FILLCELL_X1 FILLER_49_309 ();
 FILLCELL_X8 FILLER_49_326 ();
 FILLCELL_X4 FILLER_49_334 ();
 FILLCELL_X4 FILLER_49_354 ();
 FILLCELL_X2 FILLER_49_364 ();
 FILLCELL_X1 FILLER_49_366 ();
 FILLCELL_X1 FILLER_49_388 ();
 FILLCELL_X4 FILLER_49_408 ();
 FILLCELL_X4 FILLER_49_422 ();
 FILLCELL_X1 FILLER_49_426 ();
 FILLCELL_X2 FILLER_49_439 ();
 FILLCELL_X1 FILLER_49_441 ();
 FILLCELL_X1 FILLER_49_444 ();
 FILLCELL_X8 FILLER_49_455 ();
 FILLCELL_X4 FILLER_49_463 ();
 FILLCELL_X1 FILLER_49_467 ();
 FILLCELL_X4 FILLER_49_494 ();
 FILLCELL_X1 FILLER_49_498 ();
 FILLCELL_X1 FILLER_49_535 ();
 FILLCELL_X2 FILLER_50_1 ();
 FILLCELL_X2 FILLER_50_9 ();
 FILLCELL_X1 FILLER_50_11 ();
 FILLCELL_X2 FILLER_50_15 ();
 FILLCELL_X1 FILLER_50_17 ();
 FILLCELL_X16 FILLER_50_23 ();
 FILLCELL_X2 FILLER_50_43 ();
 FILLCELL_X1 FILLER_50_45 ();
 FILLCELL_X2 FILLER_50_49 ();
 FILLCELL_X1 FILLER_50_51 ();
 FILLCELL_X1 FILLER_50_54 ();
 FILLCELL_X8 FILLER_50_58 ();
 FILLCELL_X2 FILLER_50_66 ();
 FILLCELL_X1 FILLER_50_68 ();
 FILLCELL_X4 FILLER_50_82 ();
 FILLCELL_X2 FILLER_50_88 ();
 FILLCELL_X1 FILLER_50_90 ();
 FILLCELL_X1 FILLER_50_95 ();
 FILLCELL_X8 FILLER_50_102 ();
 FILLCELL_X1 FILLER_50_114 ();
 FILLCELL_X1 FILLER_50_127 ();
 FILLCELL_X4 FILLER_50_138 ();
 FILLCELL_X2 FILLER_50_142 ();
 FILLCELL_X8 FILLER_50_146 ();
 FILLCELL_X1 FILLER_50_154 ();
 FILLCELL_X4 FILLER_50_163 ();
 FILLCELL_X2 FILLER_50_177 ();
 FILLCELL_X4 FILLER_50_195 ();
 FILLCELL_X1 FILLER_50_199 ();
 FILLCELL_X8 FILLER_50_226 ();
 FILLCELL_X4 FILLER_50_234 ();
 FILLCELL_X1 FILLER_50_238 ();
 FILLCELL_X4 FILLER_50_249 ();
 FILLCELL_X2 FILLER_50_253 ();
 FILLCELL_X1 FILLER_50_265 ();
 FILLCELL_X1 FILLER_50_280 ();
 FILLCELL_X2 FILLER_50_283 ();
 FILLCELL_X1 FILLER_50_301 ();
 FILLCELL_X8 FILLER_50_322 ();
 FILLCELL_X2 FILLER_50_330 ();
 FILLCELL_X8 FILLER_50_346 ();
 FILLCELL_X4 FILLER_50_354 ();
 FILLCELL_X1 FILLER_50_358 ();
 FILLCELL_X4 FILLER_50_367 ();
 FILLCELL_X2 FILLER_50_384 ();
 FILLCELL_X1 FILLER_50_386 ();
 FILLCELL_X2 FILLER_50_449 ();
 FILLCELL_X1 FILLER_50_454 ();
 FILLCELL_X4 FILLER_50_472 ();
 FILLCELL_X2 FILLER_50_476 ();
 FILLCELL_X8 FILLER_50_485 ();
 FILLCELL_X1 FILLER_50_493 ();
 FILLCELL_X8 FILLER_50_511 ();
 FILLCELL_X2 FILLER_50_519 ();
 FILLCELL_X4 FILLER_51_1 ();
 FILLCELL_X2 FILLER_51_7 ();
 FILLCELL_X2 FILLER_51_26 ();
 FILLCELL_X1 FILLER_51_28 ();
 FILLCELL_X2 FILLER_51_39 ();
 FILLCELL_X2 FILLER_51_55 ();
 FILLCELL_X2 FILLER_51_81 ();
 FILLCELL_X1 FILLER_51_90 ();
 FILLCELL_X1 FILLER_51_123 ();
 FILLCELL_X4 FILLER_51_133 ();
 FILLCELL_X2 FILLER_51_137 ();
 FILLCELL_X1 FILLER_51_139 ();
 FILLCELL_X2 FILLER_51_168 ();
 FILLCELL_X8 FILLER_51_180 ();
 FILLCELL_X1 FILLER_51_188 ();
 FILLCELL_X8 FILLER_51_192 ();
 FILLCELL_X2 FILLER_51_200 ();
 FILLCELL_X1 FILLER_51_202 ();
 FILLCELL_X4 FILLER_51_207 ();
 FILLCELL_X8 FILLER_51_224 ();
 FILLCELL_X4 FILLER_51_232 ();
 FILLCELL_X2 FILLER_51_236 ();
 FILLCELL_X8 FILLER_51_256 ();
 FILLCELL_X4 FILLER_51_264 ();
 FILLCELL_X2 FILLER_51_268 ();
 FILLCELL_X1 FILLER_51_270 ();
 FILLCELL_X2 FILLER_51_283 ();
 FILLCELL_X1 FILLER_51_285 ();
 FILLCELL_X8 FILLER_51_292 ();
 FILLCELL_X4 FILLER_51_300 ();
 FILLCELL_X2 FILLER_51_304 ();
 FILLCELL_X1 FILLER_51_306 ();
 FILLCELL_X8 FILLER_51_322 ();
 FILLCELL_X2 FILLER_51_330 ();
 FILLCELL_X1 FILLER_51_332 ();
 FILLCELL_X1 FILLER_51_351 ();
 FILLCELL_X16 FILLER_51_366 ();
 FILLCELL_X8 FILLER_51_382 ();
 FILLCELL_X1 FILLER_51_390 ();
 FILLCELL_X2 FILLER_51_400 ();
 FILLCELL_X2 FILLER_51_415 ();
 FILLCELL_X1 FILLER_51_441 ();
 FILLCELL_X16 FILLER_51_460 ();
 FILLCELL_X2 FILLER_51_476 ();
 FILLCELL_X2 FILLER_51_492 ();
 FILLCELL_X1 FILLER_51_494 ();
 FILLCELL_X4 FILLER_51_506 ();
 FILLCELL_X16 FILLER_51_520 ();
 FILLCELL_X2 FILLER_52_1 ();
 FILLCELL_X8 FILLER_52_13 ();
 FILLCELL_X1 FILLER_52_21 ();
 FILLCELL_X2 FILLER_52_36 ();
 FILLCELL_X1 FILLER_52_38 ();
 FILLCELL_X1 FILLER_52_43 ();
 FILLCELL_X4 FILLER_52_47 ();
 FILLCELL_X2 FILLER_52_51 ();
 FILLCELL_X2 FILLER_52_56 ();
 FILLCELL_X1 FILLER_52_58 ();
 FILLCELL_X8 FILLER_52_82 ();
 FILLCELL_X2 FILLER_52_90 ();
 FILLCELL_X16 FILLER_52_126 ();
 FILLCELL_X2 FILLER_52_142 ();
 FILLCELL_X1 FILLER_52_144 ();
 FILLCELL_X2 FILLER_52_153 ();
 FILLCELL_X1 FILLER_52_155 ();
 FILLCELL_X2 FILLER_52_184 ();
 FILLCELL_X1 FILLER_52_186 ();
 FILLCELL_X2 FILLER_52_256 ();
 FILLCELL_X4 FILLER_52_268 ();
 FILLCELL_X2 FILLER_52_279 ();
 FILLCELL_X8 FILLER_52_293 ();
 FILLCELL_X1 FILLER_52_317 ();
 FILLCELL_X16 FILLER_52_335 ();
 FILLCELL_X8 FILLER_52_351 ();
 FILLCELL_X4 FILLER_52_359 ();
 FILLCELL_X2 FILLER_52_363 ();
 FILLCELL_X8 FILLER_52_373 ();
 FILLCELL_X2 FILLER_52_381 ();
 FILLCELL_X4 FILLER_52_393 ();
 FILLCELL_X4 FILLER_52_414 ();
 FILLCELL_X2 FILLER_52_418 ();
 FILLCELL_X1 FILLER_52_420 ();
 FILLCELL_X1 FILLER_52_430 ();
 FILLCELL_X8 FILLER_52_451 ();
 FILLCELL_X1 FILLER_52_459 ();
 FILLCELL_X4 FILLER_52_479 ();
 FILLCELL_X8 FILLER_52_493 ();
 FILLCELL_X4 FILLER_52_501 ();
 FILLCELL_X4 FILLER_52_508 ();
 FILLCELL_X2 FILLER_52_512 ();
 FILLCELL_X1 FILLER_52_520 ();
 FILLCELL_X4 FILLER_52_531 ();
 FILLCELL_X1 FILLER_52_535 ();
 FILLCELL_X4 FILLER_53_1 ();
 FILLCELL_X2 FILLER_53_5 ();
 FILLCELL_X4 FILLER_53_16 ();
 FILLCELL_X1 FILLER_53_34 ();
 FILLCELL_X2 FILLER_53_42 ();
 FILLCELL_X1 FILLER_53_53 ();
 FILLCELL_X2 FILLER_53_64 ();
 FILLCELL_X4 FILLER_53_70 ();
 FILLCELL_X8 FILLER_53_93 ();
 FILLCELL_X2 FILLER_53_101 ();
 FILLCELL_X1 FILLER_53_103 ();
 FILLCELL_X1 FILLER_53_106 ();
 FILLCELL_X1 FILLER_53_114 ();
 FILLCELL_X1 FILLER_53_117 ();
 FILLCELL_X2 FILLER_53_122 ();
 FILLCELL_X4 FILLER_53_129 ();
 FILLCELL_X2 FILLER_53_133 ();
 FILLCELL_X1 FILLER_53_135 ();
 FILLCELL_X4 FILLER_53_152 ();
 FILLCELL_X1 FILLER_53_161 ();
 FILLCELL_X16 FILLER_53_172 ();
 FILLCELL_X2 FILLER_53_188 ();
 FILLCELL_X2 FILLER_53_200 ();
 FILLCELL_X1 FILLER_53_202 ();
 FILLCELL_X1 FILLER_53_209 ();
 FILLCELL_X16 FILLER_53_216 ();
 FILLCELL_X2 FILLER_53_232 ();
 FILLCELL_X4 FILLER_53_236 ();
 FILLCELL_X2 FILLER_53_240 ();
 FILLCELL_X2 FILLER_53_246 ();
 FILLCELL_X8 FILLER_53_252 ();
 FILLCELL_X1 FILLER_53_260 ();
 FILLCELL_X8 FILLER_53_271 ();
 FILLCELL_X2 FILLER_53_279 ();
 FILLCELL_X8 FILLER_53_284 ();
 FILLCELL_X2 FILLER_53_292 ();
 FILLCELL_X16 FILLER_53_302 ();
 FILLCELL_X2 FILLER_53_318 ();
 FILLCELL_X2 FILLER_53_326 ();
 FILLCELL_X2 FILLER_53_337 ();
 FILLCELL_X1 FILLER_53_339 ();
 FILLCELL_X1 FILLER_53_350 ();
 FILLCELL_X1 FILLER_53_361 ();
 FILLCELL_X2 FILLER_53_375 ();
 FILLCELL_X8 FILLER_53_383 ();
 FILLCELL_X4 FILLER_53_391 ();
 FILLCELL_X2 FILLER_53_395 ();
 FILLCELL_X1 FILLER_53_397 ();
 FILLCELL_X4 FILLER_53_406 ();
 FILLCELL_X2 FILLER_53_410 ();
 FILLCELL_X4 FILLER_53_422 ();
 FILLCELL_X1 FILLER_53_426 ();
 FILLCELL_X16 FILLER_53_437 ();
 FILLCELL_X8 FILLER_53_453 ();
 FILLCELL_X4 FILLER_53_461 ();
 FILLCELL_X2 FILLER_53_465 ();
 FILLCELL_X2 FILLER_53_482 ();
 FILLCELL_X1 FILLER_53_484 ();
 FILLCELL_X2 FILLER_53_494 ();
 FILLCELL_X1 FILLER_53_503 ();
 FILLCELL_X16 FILLER_53_514 ();
 FILLCELL_X4 FILLER_53_530 ();
 FILLCELL_X2 FILLER_53_534 ();
 FILLCELL_X8 FILLER_54_1 ();
 FILLCELL_X4 FILLER_54_19 ();
 FILLCELL_X2 FILLER_54_23 ();
 FILLCELL_X1 FILLER_54_33 ();
 FILLCELL_X1 FILLER_54_38 ();
 FILLCELL_X1 FILLER_54_43 ();
 FILLCELL_X1 FILLER_54_54 ();
 FILLCELL_X4 FILLER_54_59 ();
 FILLCELL_X2 FILLER_54_70 ();
 FILLCELL_X1 FILLER_54_72 ();
 FILLCELL_X1 FILLER_54_75 ();
 FILLCELL_X2 FILLER_54_89 ();
 FILLCELL_X8 FILLER_54_113 ();
 FILLCELL_X1 FILLER_54_124 ();
 FILLCELL_X4 FILLER_54_140 ();
 FILLCELL_X1 FILLER_54_144 ();
 FILLCELL_X8 FILLER_54_157 ();
 FILLCELL_X1 FILLER_54_165 ();
 FILLCELL_X8 FILLER_54_187 ();
 FILLCELL_X4 FILLER_54_199 ();
 FILLCELL_X4 FILLER_54_212 ();
 FILLCELL_X2 FILLER_54_216 ();
 FILLCELL_X1 FILLER_54_218 ();
 FILLCELL_X1 FILLER_54_229 ();
 FILLCELL_X1 FILLER_54_240 ();
 FILLCELL_X4 FILLER_54_247 ();
 FILLCELL_X2 FILLER_54_251 ();
 FILLCELL_X1 FILLER_54_261 ();
 FILLCELL_X1 FILLER_54_269 ();
 FILLCELL_X8 FILLER_54_276 ();
 FILLCELL_X1 FILLER_54_288 ();
 FILLCELL_X1 FILLER_54_296 ();
 FILLCELL_X1 FILLER_54_301 ();
 FILLCELL_X2 FILLER_54_312 ();
 FILLCELL_X2 FILLER_54_356 ();
 FILLCELL_X1 FILLER_54_358 ();
 FILLCELL_X1 FILLER_54_369 ();
 FILLCELL_X2 FILLER_54_377 ();
 FILLCELL_X2 FILLER_54_410 ();
 FILLCELL_X2 FILLER_54_421 ();
 FILLCELL_X1 FILLER_54_423 ();
 FILLCELL_X4 FILLER_54_432 ();
 FILLCELL_X2 FILLER_54_436 ();
 FILLCELL_X2 FILLER_54_447 ();
 FILLCELL_X4 FILLER_54_452 ();
 FILLCELL_X1 FILLER_54_456 ();
 FILLCELL_X2 FILLER_54_469 ();
 FILLCELL_X1 FILLER_54_471 ();
 FILLCELL_X4 FILLER_54_485 ();
 FILLCELL_X8 FILLER_55_1 ();
 FILLCELL_X4 FILLER_55_9 ();
 FILLCELL_X8 FILLER_55_18 ();
 FILLCELL_X4 FILLER_55_26 ();
 FILLCELL_X4 FILLER_55_38 ();
 FILLCELL_X2 FILLER_55_42 ();
 FILLCELL_X1 FILLER_55_44 ();
 FILLCELL_X8 FILLER_55_49 ();
 FILLCELL_X1 FILLER_55_57 ();
 FILLCELL_X4 FILLER_55_88 ();
 FILLCELL_X1 FILLER_55_92 ();
 FILLCELL_X16 FILLER_55_98 ();
 FILLCELL_X4 FILLER_55_114 ();
 FILLCELL_X2 FILLER_55_118 ();
 FILLCELL_X1 FILLER_55_120 ();
 FILLCELL_X2 FILLER_55_125 ();
 FILLCELL_X8 FILLER_55_137 ();
 FILLCELL_X2 FILLER_55_154 ();
 FILLCELL_X4 FILLER_55_166 ();
 FILLCELL_X1 FILLER_55_170 ();
 FILLCELL_X1 FILLER_55_175 ();
 FILLCELL_X1 FILLER_55_178 ();
 FILLCELL_X2 FILLER_55_181 ();
 FILLCELL_X2 FILLER_55_193 ();
 FILLCELL_X2 FILLER_55_199 ();
 FILLCELL_X4 FILLER_55_211 ();
 FILLCELL_X2 FILLER_55_215 ();
 FILLCELL_X1 FILLER_55_217 ();
 FILLCELL_X16 FILLER_55_220 ();
 FILLCELL_X4 FILLER_55_236 ();
 FILLCELL_X2 FILLER_55_240 ();
 FILLCELL_X1 FILLER_55_242 ();
 FILLCELL_X2 FILLER_55_245 ();
 FILLCELL_X1 FILLER_55_257 ();
 FILLCELL_X2 FILLER_55_268 ();
 FILLCELL_X8 FILLER_55_289 ();
 FILLCELL_X8 FILLER_55_314 ();
 FILLCELL_X2 FILLER_55_322 ();
 FILLCELL_X1 FILLER_55_324 ();
 FILLCELL_X16 FILLER_55_327 ();
 FILLCELL_X4 FILLER_55_343 ();
 FILLCELL_X1 FILLER_55_347 ();
 FILLCELL_X1 FILLER_55_376 ();
 FILLCELL_X2 FILLER_55_383 ();
 FILLCELL_X1 FILLER_55_385 ();
 FILLCELL_X2 FILLER_55_398 ();
 FILLCELL_X8 FILLER_55_403 ();
 FILLCELL_X1 FILLER_55_417 ();
 FILLCELL_X1 FILLER_55_425 ();
 FILLCELL_X1 FILLER_55_429 ();
 FILLCELL_X2 FILLER_55_434 ();
 FILLCELL_X1 FILLER_55_459 ();
 FILLCELL_X2 FILLER_55_492 ();
 FILLCELL_X8 FILLER_55_504 ();
 FILLCELL_X1 FILLER_55_522 ();
 FILLCELL_X2 FILLER_56_1 ();
 FILLCELL_X1 FILLER_56_3 ();
 FILLCELL_X4 FILLER_56_9 ();
 FILLCELL_X4 FILLER_56_26 ();
 FILLCELL_X1 FILLER_56_72 ();
 FILLCELL_X8 FILLER_56_82 ();
 FILLCELL_X2 FILLER_56_90 ();
 FILLCELL_X1 FILLER_56_92 ();
 FILLCELL_X4 FILLER_56_112 ();
 FILLCELL_X2 FILLER_56_116 ();
 FILLCELL_X4 FILLER_56_149 ();
 FILLCELL_X1 FILLER_56_163 ();
 FILLCELL_X1 FILLER_56_175 ();
 FILLCELL_X1 FILLER_56_183 ();
 FILLCELL_X1 FILLER_56_196 ();
 FILLCELL_X4 FILLER_56_210 ();
 FILLCELL_X4 FILLER_56_233 ();
 FILLCELL_X1 FILLER_56_237 ();
 FILLCELL_X2 FILLER_56_310 ();
 FILLCELL_X1 FILLER_56_312 ();
 FILLCELL_X4 FILLER_56_332 ();
 FILLCELL_X1 FILLER_56_336 ();
 FILLCELL_X4 FILLER_56_339 ();
 FILLCELL_X2 FILLER_56_343 ();
 FILLCELL_X1 FILLER_56_345 ();
 FILLCELL_X1 FILLER_56_356 ();
 FILLCELL_X4 FILLER_56_361 ();
 FILLCELL_X1 FILLER_56_365 ();
 FILLCELL_X1 FILLER_56_376 ();
 FILLCELL_X1 FILLER_56_387 ();
 FILLCELL_X1 FILLER_56_395 ();
 FILLCELL_X4 FILLER_56_398 ();
 FILLCELL_X2 FILLER_56_402 ();
 FILLCELL_X8 FILLER_56_417 ();
 FILLCELL_X4 FILLER_56_425 ();
 FILLCELL_X1 FILLER_56_429 ();
 FILLCELL_X4 FILLER_56_436 ();
 FILLCELL_X1 FILLER_56_476 ();
 FILLCELL_X2 FILLER_56_505 ();
 FILLCELL_X2 FILLER_56_511 ();
 FILLCELL_X1 FILLER_56_535 ();
 FILLCELL_X4 FILLER_57_1 ();
 FILLCELL_X2 FILLER_57_5 ();
 FILLCELL_X4 FILLER_57_11 ();
 FILLCELL_X2 FILLER_57_15 ();
 FILLCELL_X4 FILLER_57_26 ();
 FILLCELL_X1 FILLER_57_37 ();
 FILLCELL_X1 FILLER_57_43 ();
 FILLCELL_X2 FILLER_57_56 ();
 FILLCELL_X1 FILLER_57_61 ();
 FILLCELL_X2 FILLER_57_69 ();
 FILLCELL_X32 FILLER_57_74 ();
 FILLCELL_X2 FILLER_57_106 ();
 FILLCELL_X1 FILLER_57_108 ();
 FILLCELL_X8 FILLER_57_118 ();
 FILLCELL_X4 FILLER_57_126 ();
 FILLCELL_X2 FILLER_57_130 ();
 FILLCELL_X2 FILLER_57_138 ();
 FILLCELL_X1 FILLER_57_149 ();
 FILLCELL_X2 FILLER_57_160 ();
 FILLCELL_X1 FILLER_57_162 ();
 FILLCELL_X2 FILLER_57_165 ();
 FILLCELL_X2 FILLER_57_174 ();
 FILLCELL_X1 FILLER_57_176 ();
 FILLCELL_X2 FILLER_57_187 ();
 FILLCELL_X1 FILLER_57_189 ();
 FILLCELL_X2 FILLER_57_194 ();
 FILLCELL_X32 FILLER_57_208 ();
 FILLCELL_X1 FILLER_57_240 ();
 FILLCELL_X2 FILLER_57_245 ();
 FILLCELL_X1 FILLER_57_250 ();
 FILLCELL_X2 FILLER_57_259 ();
 FILLCELL_X1 FILLER_57_271 ();
 FILLCELL_X1 FILLER_57_276 ();
 FILLCELL_X2 FILLER_57_287 ();
 FILLCELL_X1 FILLER_57_299 ();
 FILLCELL_X1 FILLER_57_306 ();
 FILLCELL_X1 FILLER_57_311 ();
 FILLCELL_X4 FILLER_57_319 ();
 FILLCELL_X2 FILLER_57_330 ();
 FILLCELL_X16 FILLER_57_376 ();
 FILLCELL_X8 FILLER_57_392 ();
 FILLCELL_X4 FILLER_57_400 ();
 FILLCELL_X2 FILLER_57_414 ();
 FILLCELL_X4 FILLER_57_476 ();
 FILLCELL_X2 FILLER_57_480 ();
 FILLCELL_X1 FILLER_57_482 ();
 FILLCELL_X8 FILLER_57_497 ();
 FILLCELL_X2 FILLER_57_512 ();
 FILLCELL_X1 FILLER_57_514 ();
 FILLCELL_X2 FILLER_57_525 ();
 FILLCELL_X4 FILLER_58_1 ();
 FILLCELL_X4 FILLER_58_9 ();
 FILLCELL_X2 FILLER_58_13 ();
 FILLCELL_X1 FILLER_58_15 ();
 FILLCELL_X4 FILLER_58_24 ();
 FILLCELL_X2 FILLER_58_37 ();
 FILLCELL_X1 FILLER_58_39 ();
 FILLCELL_X1 FILLER_58_52 ();
 FILLCELL_X4 FILLER_58_56 ();
 FILLCELL_X1 FILLER_58_69 ();
 FILLCELL_X4 FILLER_58_80 ();
 FILLCELL_X2 FILLER_58_84 ();
 FILLCELL_X2 FILLER_58_91 ();
 FILLCELL_X8 FILLER_58_97 ();
 FILLCELL_X2 FILLER_58_105 ();
 FILLCELL_X1 FILLER_58_113 ();
 FILLCELL_X2 FILLER_58_129 ();
 FILLCELL_X8 FILLER_58_147 ();
 FILLCELL_X2 FILLER_58_155 ();
 FILLCELL_X1 FILLER_58_157 ();
 FILLCELL_X2 FILLER_58_162 ();
 FILLCELL_X2 FILLER_58_166 ();
 FILLCELL_X4 FILLER_58_178 ();
 FILLCELL_X1 FILLER_58_192 ();
 FILLCELL_X4 FILLER_58_206 ();
 FILLCELL_X1 FILLER_58_210 ();
 FILLCELL_X1 FILLER_58_223 ();
 FILLCELL_X8 FILLER_58_227 ();
 FILLCELL_X2 FILLER_58_235 ();
 FILLCELL_X1 FILLER_58_237 ();
 FILLCELL_X1 FILLER_58_242 ();
 FILLCELL_X1 FILLER_58_245 ();
 FILLCELL_X8 FILLER_58_259 ();
 FILLCELL_X4 FILLER_58_267 ();
 FILLCELL_X16 FILLER_58_287 ();
 FILLCELL_X4 FILLER_58_303 ();
 FILLCELL_X2 FILLER_58_307 ();
 FILLCELL_X1 FILLER_58_309 ();
 FILLCELL_X2 FILLER_58_331 ();
 FILLCELL_X2 FILLER_58_340 ();
 FILLCELL_X2 FILLER_58_347 ();
 FILLCELL_X4 FILLER_58_352 ();
 FILLCELL_X2 FILLER_58_356 ();
 FILLCELL_X1 FILLER_58_358 ();
 FILLCELL_X8 FILLER_58_376 ();
 FILLCELL_X4 FILLER_58_384 ();
 FILLCELL_X1 FILLER_58_388 ();
 FILLCELL_X2 FILLER_58_424 ();
 FILLCELL_X1 FILLER_58_426 ();
 FILLCELL_X1 FILLER_58_452 ();
 FILLCELL_X1 FILLER_58_466 ();
 FILLCELL_X1 FILLER_58_478 ();
 FILLCELL_X2 FILLER_58_492 ();
 FILLCELL_X4 FILLER_58_511 ();
 FILLCELL_X1 FILLER_58_515 ();
 FILLCELL_X1 FILLER_59_1 ();
 FILLCELL_X4 FILLER_59_15 ();
 FILLCELL_X1 FILLER_59_19 ();
 FILLCELL_X2 FILLER_59_29 ();
 FILLCELL_X1 FILLER_59_31 ();
 FILLCELL_X2 FILLER_59_48 ();
 FILLCELL_X1 FILLER_59_50 ();
 FILLCELL_X8 FILLER_59_63 ();
 FILLCELL_X4 FILLER_59_71 ();
 FILLCELL_X2 FILLER_59_75 ();
 FILLCELL_X1 FILLER_59_90 ();
 FILLCELL_X8 FILLER_59_99 ();
 FILLCELL_X2 FILLER_59_107 ();
 FILLCELL_X1 FILLER_59_109 ();
 FILLCELL_X2 FILLER_59_116 ();
 FILLCELL_X4 FILLER_59_124 ();
 FILLCELL_X2 FILLER_59_128 ();
 FILLCELL_X1 FILLER_59_130 ();
 FILLCELL_X8 FILLER_59_136 ();
 FILLCELL_X4 FILLER_59_144 ();
 FILLCELL_X2 FILLER_59_148 ();
 FILLCELL_X1 FILLER_59_150 ();
 FILLCELL_X2 FILLER_59_162 ();
 FILLCELL_X2 FILLER_59_170 ();
 FILLCELL_X1 FILLER_59_172 ();
 FILLCELL_X2 FILLER_59_187 ();
 FILLCELL_X8 FILLER_59_206 ();
 FILLCELL_X1 FILLER_59_214 ();
 FILLCELL_X16 FILLER_59_229 ();
 FILLCELL_X2 FILLER_59_245 ();
 FILLCELL_X2 FILLER_59_250 ();
 FILLCELL_X1 FILLER_59_258 ();
 FILLCELL_X1 FILLER_59_275 ();
 FILLCELL_X4 FILLER_59_290 ();
 FILLCELL_X4 FILLER_59_321 ();
 FILLCELL_X8 FILLER_59_335 ();
 FILLCELL_X2 FILLER_59_345 ();
 FILLCELL_X1 FILLER_59_347 ();
 FILLCELL_X1 FILLER_59_367 ();
 FILLCELL_X1 FILLER_59_371 ();
 FILLCELL_X1 FILLER_59_395 ();
 FILLCELL_X2 FILLER_59_406 ();
 FILLCELL_X4 FILLER_59_414 ();
 FILLCELL_X1 FILLER_59_418 ();
 FILLCELL_X8 FILLER_59_453 ();
 FILLCELL_X1 FILLER_59_461 ();
 FILLCELL_X8 FILLER_59_476 ();
 FILLCELL_X2 FILLER_59_484 ();
 FILLCELL_X2 FILLER_59_489 ();
 FILLCELL_X1 FILLER_59_491 ();
 FILLCELL_X1 FILLER_59_502 ();
 FILLCELL_X1 FILLER_59_535 ();
 FILLCELL_X4 FILLER_60_1 ();
 FILLCELL_X1 FILLER_60_5 ();
 FILLCELL_X2 FILLER_60_24 ();
 FILLCELL_X16 FILLER_60_33 ();
 FILLCELL_X1 FILLER_60_49 ();
 FILLCELL_X2 FILLER_60_59 ();
 FILLCELL_X1 FILLER_60_61 ();
 FILLCELL_X4 FILLER_60_67 ();
 FILLCELL_X2 FILLER_60_71 ();
 FILLCELL_X4 FILLER_60_82 ();
 FILLCELL_X2 FILLER_60_86 ();
 FILLCELL_X1 FILLER_60_91 ();
 FILLCELL_X8 FILLER_60_96 ();
 FILLCELL_X4 FILLER_60_104 ();
 FILLCELL_X2 FILLER_60_110 ();
 FILLCELL_X1 FILLER_60_112 ();
 FILLCELL_X1 FILLER_60_116 ();
 FILLCELL_X1 FILLER_60_135 ();
 FILLCELL_X4 FILLER_60_177 ();
 FILLCELL_X2 FILLER_60_181 ();
 FILLCELL_X16 FILLER_60_198 ();
 FILLCELL_X1 FILLER_60_214 ();
 FILLCELL_X4 FILLER_60_219 ();
 FILLCELL_X2 FILLER_60_223 ();
 FILLCELL_X1 FILLER_60_225 ();
 FILLCELL_X2 FILLER_60_238 ();
 FILLCELL_X1 FILLER_60_243 ();
 FILLCELL_X1 FILLER_60_248 ();
 FILLCELL_X16 FILLER_60_260 ();
 FILLCELL_X2 FILLER_60_276 ();
 FILLCELL_X8 FILLER_60_286 ();
 FILLCELL_X2 FILLER_60_294 ();
 FILLCELL_X2 FILLER_60_300 ();
 FILLCELL_X1 FILLER_60_319 ();
 FILLCELL_X4 FILLER_60_322 ();
 FILLCELL_X4 FILLER_60_335 ();
 FILLCELL_X2 FILLER_60_339 ();
 FILLCELL_X1 FILLER_60_341 ();
 FILLCELL_X2 FILLER_60_346 ();
 FILLCELL_X1 FILLER_60_348 ();
 FILLCELL_X1 FILLER_60_374 ();
 FILLCELL_X1 FILLER_60_382 ();
 FILLCELL_X1 FILLER_60_397 ();
 FILLCELL_X8 FILLER_60_423 ();
 FILLCELL_X4 FILLER_60_431 ();
 FILLCELL_X2 FILLER_60_435 ();
 FILLCELL_X1 FILLER_60_440 ();
 FILLCELL_X1 FILLER_60_492 ();
 FILLCELL_X1 FILLER_60_522 ();
 FILLCELL_X4 FILLER_61_1 ();
 FILLCELL_X1 FILLER_61_14 ();
 FILLCELL_X4 FILLER_61_47 ();
 FILLCELL_X2 FILLER_61_51 ();
 FILLCELL_X1 FILLER_61_53 ();
 FILLCELL_X1 FILLER_61_64 ();
 FILLCELL_X4 FILLER_61_68 ();
 FILLCELL_X1 FILLER_61_79 ();
 FILLCELL_X4 FILLER_61_101 ();
 FILLCELL_X4 FILLER_61_108 ();
 FILLCELL_X1 FILLER_61_112 ();
 FILLCELL_X16 FILLER_61_122 ();
 FILLCELL_X4 FILLER_61_138 ();
 FILLCELL_X2 FILLER_61_142 ();
 FILLCELL_X4 FILLER_61_163 ();
 FILLCELL_X2 FILLER_61_167 ();
 FILLCELL_X1 FILLER_61_169 ();
 FILLCELL_X2 FILLER_61_180 ();
 FILLCELL_X2 FILLER_61_184 ();
 FILLCELL_X1 FILLER_61_186 ();
 FILLCELL_X16 FILLER_61_197 ();
 FILLCELL_X4 FILLER_61_213 ();
 FILLCELL_X1 FILLER_61_217 ();
 FILLCELL_X2 FILLER_61_221 ();
 FILLCELL_X1 FILLER_61_223 ();
 FILLCELL_X1 FILLER_61_251 ();
 FILLCELL_X4 FILLER_61_271 ();
 FILLCELL_X1 FILLER_61_275 ();
 FILLCELL_X4 FILLER_61_289 ();
 FILLCELL_X1 FILLER_61_293 ();
 FILLCELL_X1 FILLER_61_304 ();
 FILLCELL_X2 FILLER_61_313 ();
 FILLCELL_X4 FILLER_61_319 ();
 FILLCELL_X2 FILLER_61_323 ();
 FILLCELL_X8 FILLER_61_331 ();
 FILLCELL_X2 FILLER_61_352 ();
 FILLCELL_X1 FILLER_61_358 ();
 FILLCELL_X1 FILLER_61_361 ();
 FILLCELL_X1 FILLER_61_368 ();
 FILLCELL_X1 FILLER_61_393 ();
 FILLCELL_X2 FILLER_61_462 ();
 FILLCELL_X4 FILLER_61_489 ();
 FILLCELL_X2 FILLER_61_534 ();
 FILLCELL_X16 FILLER_62_1 ();
 FILLCELL_X8 FILLER_62_17 ();
 FILLCELL_X2 FILLER_62_48 ();
 FILLCELL_X1 FILLER_62_50 ();
 FILLCELL_X4 FILLER_62_74 ();
 FILLCELL_X1 FILLER_62_78 ();
 FILLCELL_X1 FILLER_62_85 ();
 FILLCELL_X2 FILLER_62_88 ();
 FILLCELL_X1 FILLER_62_90 ();
 FILLCELL_X4 FILLER_62_97 ();
 FILLCELL_X1 FILLER_62_101 ();
 FILLCELL_X1 FILLER_62_131 ();
 FILLCELL_X1 FILLER_62_134 ();
 FILLCELL_X4 FILLER_62_154 ();
 FILLCELL_X8 FILLER_62_172 ();
 FILLCELL_X4 FILLER_62_180 ();
 FILLCELL_X2 FILLER_62_184 ();
 FILLCELL_X8 FILLER_62_199 ();
 FILLCELL_X2 FILLER_62_207 ();
 FILLCELL_X1 FILLER_62_209 ();
 FILLCELL_X4 FILLER_62_216 ();
 FILLCELL_X1 FILLER_62_220 ();
 FILLCELL_X1 FILLER_62_224 ();
 FILLCELL_X2 FILLER_62_244 ();
 FILLCELL_X2 FILLER_62_255 ();
 FILLCELL_X2 FILLER_62_267 ();
 FILLCELL_X2 FILLER_62_284 ();
 FILLCELL_X16 FILLER_62_296 ();
 FILLCELL_X4 FILLER_62_312 ();
 FILLCELL_X1 FILLER_62_316 ();
 FILLCELL_X4 FILLER_62_332 ();
 FILLCELL_X16 FILLER_62_339 ();
 FILLCELL_X4 FILLER_62_355 ();
 FILLCELL_X8 FILLER_62_396 ();
 FILLCELL_X2 FILLER_62_404 ();
 FILLCELL_X8 FILLER_62_426 ();
 FILLCELL_X4 FILLER_62_434 ();
 FILLCELL_X2 FILLER_62_438 ();
 FILLCELL_X1 FILLER_62_440 ();
 FILLCELL_X8 FILLER_62_476 ();
 FILLCELL_X2 FILLER_62_484 ();
 FILLCELL_X2 FILLER_62_506 ();
 FILLCELL_X1 FILLER_62_508 ();
 FILLCELL_X8 FILLER_62_523 ();
 FILLCELL_X4 FILLER_62_531 ();
 FILLCELL_X1 FILLER_62_535 ();
 FILLCELL_X8 FILLER_63_1 ();
 FILLCELL_X4 FILLER_63_40 ();
 FILLCELL_X2 FILLER_63_44 ();
 FILLCELL_X1 FILLER_63_46 ();
 FILLCELL_X1 FILLER_63_64 ();
 FILLCELL_X4 FILLER_63_75 ();
 FILLCELL_X1 FILLER_63_88 ();
 FILLCELL_X8 FILLER_63_105 ();
 FILLCELL_X2 FILLER_63_121 ();
 FILLCELL_X1 FILLER_63_144 ();
 FILLCELL_X8 FILLER_63_155 ();
 FILLCELL_X4 FILLER_63_163 ();
 FILLCELL_X2 FILLER_63_167 ();
 FILLCELL_X1 FILLER_63_169 ();
 FILLCELL_X8 FILLER_63_202 ();
 FILLCELL_X4 FILLER_63_210 ();
 FILLCELL_X1 FILLER_63_218 ();
 FILLCELL_X2 FILLER_63_233 ();
 FILLCELL_X1 FILLER_63_235 ();
 FILLCELL_X2 FILLER_63_251 ();
 FILLCELL_X1 FILLER_63_255 ();
 FILLCELL_X1 FILLER_63_266 ();
 FILLCELL_X2 FILLER_63_292 ();
 FILLCELL_X1 FILLER_63_294 ();
 FILLCELL_X1 FILLER_63_316 ();
 FILLCELL_X2 FILLER_63_331 ();
 FILLCELL_X1 FILLER_63_354 ();
 FILLCELL_X16 FILLER_63_382 ();
 FILLCELL_X8 FILLER_63_427 ();
 FILLCELL_X4 FILLER_63_435 ();
 FILLCELL_X2 FILLER_63_439 ();
 FILLCELL_X1 FILLER_63_441 ();
 FILLCELL_X1 FILLER_63_461 ();
 FILLCELL_X4 FILLER_63_465 ();
 FILLCELL_X2 FILLER_63_469 ();
 FILLCELL_X8 FILLER_63_481 ();
 FILLCELL_X4 FILLER_63_489 ();
 FILLCELL_X2 FILLER_63_493 ();
 FILLCELL_X32 FILLER_63_499 ();
 FILLCELL_X4 FILLER_63_531 ();
 FILLCELL_X1 FILLER_63_535 ();
 FILLCELL_X8 FILLER_64_1 ();
 FILLCELL_X2 FILLER_64_9 ();
 FILLCELL_X1 FILLER_64_11 ();
 FILLCELL_X4 FILLER_64_22 ();
 FILLCELL_X8 FILLER_64_48 ();
 FILLCELL_X2 FILLER_64_56 ();
 FILLCELL_X1 FILLER_64_58 ();
 FILLCELL_X4 FILLER_64_63 ();
 FILLCELL_X2 FILLER_64_67 ();
 FILLCELL_X8 FILLER_64_92 ();
 FILLCELL_X1 FILLER_64_100 ();
 FILLCELL_X2 FILLER_64_111 ();
 FILLCELL_X1 FILLER_64_113 ();
 FILLCELL_X1 FILLER_64_130 ();
 FILLCELL_X1 FILLER_64_151 ();
 FILLCELL_X4 FILLER_64_162 ();
 FILLCELL_X1 FILLER_64_166 ();
 FILLCELL_X1 FILLER_64_169 ();
 FILLCELL_X4 FILLER_64_177 ();
 FILLCELL_X2 FILLER_64_181 ();
 FILLCELL_X4 FILLER_64_193 ();
 FILLCELL_X2 FILLER_64_197 ();
 FILLCELL_X4 FILLER_64_217 ();
 FILLCELL_X1 FILLER_64_221 ();
 FILLCELL_X4 FILLER_64_235 ();
 FILLCELL_X2 FILLER_64_239 ();
 FILLCELL_X1 FILLER_64_241 ();
 FILLCELL_X4 FILLER_64_249 ();
 FILLCELL_X1 FILLER_64_253 ();
 FILLCELL_X4 FILLER_64_258 ();
 FILLCELL_X4 FILLER_64_265 ();
 FILLCELL_X4 FILLER_64_285 ();
 FILLCELL_X8 FILLER_64_295 ();
 FILLCELL_X4 FILLER_64_303 ();
 FILLCELL_X2 FILLER_64_317 ();
 FILLCELL_X1 FILLER_64_319 ();
 FILLCELL_X16 FILLER_64_324 ();
 FILLCELL_X1 FILLER_64_388 ();
 FILLCELL_X4 FILLER_64_395 ();
 FILLCELL_X2 FILLER_64_399 ();
 FILLCELL_X1 FILLER_64_411 ();
 FILLCELL_X4 FILLER_64_434 ();
 FILLCELL_X4 FILLER_64_442 ();
 FILLCELL_X1 FILLER_64_456 ();
 FILLCELL_X16 FILLER_64_509 ();
 FILLCELL_X8 FILLER_64_525 ();
 FILLCELL_X2 FILLER_64_533 ();
 FILLCELL_X1 FILLER_64_535 ();
 FILLCELL_X4 FILLER_65_1 ();
 FILLCELL_X2 FILLER_65_5 ();
 FILLCELL_X1 FILLER_65_7 ();
 FILLCELL_X2 FILLER_65_31 ();
 FILLCELL_X1 FILLER_65_33 ();
 FILLCELL_X4 FILLER_65_67 ();
 FILLCELL_X2 FILLER_65_71 ();
 FILLCELL_X1 FILLER_65_73 ();
 FILLCELL_X8 FILLER_65_77 ();
 FILLCELL_X2 FILLER_65_85 ();
 FILLCELL_X4 FILLER_65_93 ();
 FILLCELL_X2 FILLER_65_110 ();
 FILLCELL_X1 FILLER_65_114 ();
 FILLCELL_X4 FILLER_65_125 ();
 FILLCELL_X4 FILLER_65_155 ();
 FILLCELL_X8 FILLER_65_181 ();
 FILLCELL_X4 FILLER_65_189 ();
 FILLCELL_X1 FILLER_65_193 ();
 FILLCELL_X2 FILLER_65_237 ();
 FILLCELL_X4 FILLER_65_248 ();
 FILLCELL_X2 FILLER_65_252 ();
 FILLCELL_X1 FILLER_65_254 ();
 FILLCELL_X2 FILLER_65_265 ();
 FILLCELL_X4 FILLER_65_279 ();
 FILLCELL_X4 FILLER_65_293 ();
 FILLCELL_X1 FILLER_65_297 ();
 FILLCELL_X2 FILLER_65_302 ();
 FILLCELL_X2 FILLER_65_306 ();
 FILLCELL_X1 FILLER_65_312 ();
 FILLCELL_X8 FILLER_65_322 ();
 FILLCELL_X2 FILLER_65_330 ();
 FILLCELL_X1 FILLER_65_390 ();
 FILLCELL_X4 FILLER_65_397 ();
 FILLCELL_X2 FILLER_65_401 ();
 FILLCELL_X1 FILLER_65_424 ();
 FILLCELL_X16 FILLER_65_442 ();
 FILLCELL_X4 FILLER_65_458 ();
 FILLCELL_X1 FILLER_65_462 ();
 FILLCELL_X2 FILLER_65_492 ();
 FILLCELL_X16 FILLER_65_505 ();
 FILLCELL_X8 FILLER_65_521 ();
 FILLCELL_X4 FILLER_65_529 ();
 FILLCELL_X2 FILLER_65_533 ();
 FILLCELL_X1 FILLER_65_535 ();
 FILLCELL_X8 FILLER_66_1 ();
 FILLCELL_X4 FILLER_66_9 ();
 FILLCELL_X2 FILLER_66_13 ();
 FILLCELL_X1 FILLER_66_15 ();
 FILLCELL_X2 FILLER_66_36 ();
 FILLCELL_X1 FILLER_66_38 ();
 FILLCELL_X1 FILLER_66_71 ();
 FILLCELL_X4 FILLER_66_78 ();
 FILLCELL_X1 FILLER_66_82 ();
 FILLCELL_X8 FILLER_66_93 ();
 FILLCELL_X4 FILLER_66_101 ();
 FILLCELL_X2 FILLER_66_123 ();
 FILLCELL_X1 FILLER_66_125 ();
 FILLCELL_X8 FILLER_66_146 ();
 FILLCELL_X2 FILLER_66_158 ();
 FILLCELL_X1 FILLER_66_160 ();
 FILLCELL_X2 FILLER_66_167 ();
 FILLCELL_X8 FILLER_66_178 ();
 FILLCELL_X1 FILLER_66_229 ();
 FILLCELL_X2 FILLER_66_243 ();
 FILLCELL_X8 FILLER_66_259 ();
 FILLCELL_X1 FILLER_66_267 ();
 FILLCELL_X2 FILLER_66_283 ();
 FILLCELL_X1 FILLER_66_285 ();
 FILLCELL_X32 FILLER_66_306 ();
 FILLCELL_X1 FILLER_66_338 ();
 FILLCELL_X2 FILLER_66_349 ();
 FILLCELL_X2 FILLER_66_382 ();
 FILLCELL_X1 FILLER_66_424 ();
 FILLCELL_X8 FILLER_66_442 ();
 FILLCELL_X8 FILLER_66_459 ();
 FILLCELL_X8 FILLER_66_477 ();
 FILLCELL_X2 FILLER_66_485 ();
 FILLCELL_X1 FILLER_66_491 ();
 FILLCELL_X32 FILLER_66_501 ();
 FILLCELL_X2 FILLER_66_533 ();
 FILLCELL_X1 FILLER_66_535 ();
 FILLCELL_X16 FILLER_67_1 ();
 FILLCELL_X2 FILLER_67_17 ();
 FILLCELL_X4 FILLER_67_30 ();
 FILLCELL_X1 FILLER_67_34 ();
 FILLCELL_X4 FILLER_67_49 ();
 FILLCELL_X1 FILLER_67_53 ();
 FILLCELL_X8 FILLER_67_78 ();
 FILLCELL_X1 FILLER_67_86 ();
 FILLCELL_X8 FILLER_67_134 ();
 FILLCELL_X4 FILLER_67_142 ();
 FILLCELL_X2 FILLER_67_146 ();
 FILLCELL_X1 FILLER_67_152 ();
 FILLCELL_X4 FILLER_67_159 ();
 FILLCELL_X2 FILLER_67_163 ();
 FILLCELL_X1 FILLER_67_165 ();
 FILLCELL_X8 FILLER_67_179 ();
 FILLCELL_X2 FILLER_67_187 ();
 FILLCELL_X1 FILLER_67_189 ();
 FILLCELL_X1 FILLER_67_224 ();
 FILLCELL_X1 FILLER_67_245 ();
 FILLCELL_X1 FILLER_67_249 ();
 FILLCELL_X2 FILLER_67_265 ();
 FILLCELL_X2 FILLER_67_273 ();
 FILLCELL_X1 FILLER_67_275 ();
 FILLCELL_X2 FILLER_67_289 ();
 FILLCELL_X4 FILLER_67_301 ();
 FILLCELL_X8 FILLER_67_334 ();
 FILLCELL_X1 FILLER_67_342 ();
 FILLCELL_X8 FILLER_67_410 ();
 FILLCELL_X1 FILLER_67_418 ();
 FILLCELL_X8 FILLER_67_421 ();
 FILLCELL_X1 FILLER_67_429 ();
 FILLCELL_X2 FILLER_67_441 ();
 FILLCELL_X2 FILLER_67_460 ();
 FILLCELL_X1 FILLER_67_462 ();
 FILLCELL_X2 FILLER_67_490 ();
 FILLCELL_X32 FILLER_67_503 ();
 FILLCELL_X1 FILLER_67_535 ();
 FILLCELL_X16 FILLER_68_1 ();
 FILLCELL_X2 FILLER_68_17 ();
 FILLCELL_X2 FILLER_68_37 ();
 FILLCELL_X1 FILLER_68_39 ();
 FILLCELL_X4 FILLER_68_57 ();
 FILLCELL_X2 FILLER_68_61 ();
 FILLCELL_X16 FILLER_68_97 ();
 FILLCELL_X4 FILLER_68_113 ();
 FILLCELL_X2 FILLER_68_117 ();
 FILLCELL_X1 FILLER_68_131 ();
 FILLCELL_X2 FILLER_68_146 ();
 FILLCELL_X4 FILLER_68_165 ();
 FILLCELL_X1 FILLER_68_169 ();
 FILLCELL_X1 FILLER_68_184 ();
 FILLCELL_X2 FILLER_68_206 ();
 FILLCELL_X1 FILLER_68_208 ();
 FILLCELL_X2 FILLER_68_245 ();
 FILLCELL_X4 FILLER_68_261 ();
 FILLCELL_X2 FILLER_68_265 ();
 FILLCELL_X1 FILLER_68_267 ();
 FILLCELL_X1 FILLER_68_289 ();
 FILLCELL_X1 FILLER_68_310 ();
 FILLCELL_X4 FILLER_68_321 ();
 FILLCELL_X1 FILLER_68_332 ();
 FILLCELL_X4 FILLER_68_343 ();
 FILLCELL_X2 FILLER_68_347 ();
 FILLCELL_X1 FILLER_68_370 ();
 FILLCELL_X1 FILLER_68_411 ();
 FILLCELL_X4 FILLER_68_425 ();
 FILLCELL_X2 FILLER_68_436 ();
 FILLCELL_X4 FILLER_68_449 ();
 FILLCELL_X2 FILLER_68_453 ();
 FILLCELL_X8 FILLER_68_462 ();
 FILLCELL_X2 FILLER_68_470 ();
 FILLCELL_X1 FILLER_68_472 ();
 FILLCELL_X1 FILLER_68_483 ();
 FILLCELL_X32 FILLER_68_498 ();
 FILLCELL_X4 FILLER_68_530 ();
 FILLCELL_X2 FILLER_68_534 ();
 FILLCELL_X16 FILLER_69_1 ();
 FILLCELL_X4 FILLER_69_17 ();
 FILLCELL_X2 FILLER_69_34 ();
 FILLCELL_X1 FILLER_69_36 ();
 FILLCELL_X2 FILLER_69_52 ();
 FILLCELL_X4 FILLER_69_67 ();
 FILLCELL_X2 FILLER_69_85 ();
 FILLCELL_X1 FILLER_69_127 ();
 FILLCELL_X8 FILLER_69_131 ();
 FILLCELL_X2 FILLER_69_139 ();
 FILLCELL_X1 FILLER_69_154 ();
 FILLCELL_X8 FILLER_69_169 ();
 FILLCELL_X4 FILLER_69_177 ();
 FILLCELL_X1 FILLER_69_218 ();
 FILLCELL_X1 FILLER_69_243 ();
 FILLCELL_X2 FILLER_69_254 ();
 FILLCELL_X1 FILLER_69_266 ();
 FILLCELL_X2 FILLER_69_269 ();
 FILLCELL_X8 FILLER_69_275 ();
 FILLCELL_X1 FILLER_69_283 ();
 FILLCELL_X8 FILLER_69_302 ();
 FILLCELL_X2 FILLER_69_321 ();
 FILLCELL_X8 FILLER_69_328 ();
 FILLCELL_X1 FILLER_69_336 ();
 FILLCELL_X16 FILLER_69_339 ();
 FILLCELL_X1 FILLER_69_385 ();
 FILLCELL_X2 FILLER_69_389 ();
 FILLCELL_X2 FILLER_69_404 ();
 FILLCELL_X2 FILLER_69_423 ();
 FILLCELL_X2 FILLER_69_429 ();
 FILLCELL_X16 FILLER_69_445 ();
 FILLCELL_X2 FILLER_69_461 ();
 FILLCELL_X2 FILLER_69_466 ();
 FILLCELL_X32 FILLER_69_501 ();
 FILLCELL_X2 FILLER_69_533 ();
 FILLCELL_X1 FILLER_69_535 ();
 FILLCELL_X32 FILLER_70_1 ();
 FILLCELL_X8 FILLER_70_33 ();
 FILLCELL_X1 FILLER_70_41 ();
 FILLCELL_X8 FILLER_70_48 ();
 FILLCELL_X1 FILLER_70_56 ();
 FILLCELL_X16 FILLER_70_63 ();
 FILLCELL_X4 FILLER_70_79 ();
 FILLCELL_X2 FILLER_70_100 ();
 FILLCELL_X1 FILLER_70_102 ();
 FILLCELL_X4 FILLER_70_113 ();
 FILLCELL_X16 FILLER_70_120 ();
 FILLCELL_X2 FILLER_70_140 ();
 FILLCELL_X1 FILLER_70_142 ();
 FILLCELL_X8 FILLER_70_157 ();
 FILLCELL_X4 FILLER_70_165 ();
 FILLCELL_X2 FILLER_70_169 ();
 FILLCELL_X4 FILLER_70_241 ();
 FILLCELL_X2 FILLER_70_248 ();
 FILLCELL_X1 FILLER_70_250 ();
 FILLCELL_X1 FILLER_70_264 ();
 FILLCELL_X2 FILLER_70_274 ();
 FILLCELL_X1 FILLER_70_276 ();
 FILLCELL_X4 FILLER_70_287 ();
 FILLCELL_X2 FILLER_70_291 ();
 FILLCELL_X2 FILLER_70_303 ();
 FILLCELL_X1 FILLER_70_305 ();
 FILLCELL_X8 FILLER_70_351 ();
 FILLCELL_X4 FILLER_70_359 ();
 FILLCELL_X1 FILLER_70_363 ();
 FILLCELL_X1 FILLER_70_379 ();
 FILLCELL_X1 FILLER_70_393 ();
 FILLCELL_X1 FILLER_70_414 ();
 FILLCELL_X2 FILLER_70_433 ();
 FILLCELL_X2 FILLER_70_442 ();
 FILLCELL_X1 FILLER_70_452 ();
 FILLCELL_X16 FILLER_70_457 ();
 FILLCELL_X4 FILLER_70_473 ();
 FILLCELL_X4 FILLER_70_484 ();
 FILLCELL_X1 FILLER_70_488 ();
 FILLCELL_X32 FILLER_70_498 ();
 FILLCELL_X4 FILLER_70_530 ();
 FILLCELL_X2 FILLER_70_534 ();
 FILLCELL_X32 FILLER_71_1 ();
 FILLCELL_X8 FILLER_71_33 ();
 FILLCELL_X1 FILLER_71_41 ();
 FILLCELL_X4 FILLER_71_51 ();
 FILLCELL_X2 FILLER_71_55 ();
 FILLCELL_X1 FILLER_71_57 ();
 FILLCELL_X32 FILLER_71_65 ();
 FILLCELL_X32 FILLER_71_97 ();
 FILLCELL_X4 FILLER_71_129 ();
 FILLCELL_X2 FILLER_71_133 ();
 FILLCELL_X1 FILLER_71_135 ();
 FILLCELL_X2 FILLER_71_144 ();
 FILLCELL_X32 FILLER_71_153 ();
 FILLCELL_X1 FILLER_71_185 ();
 FILLCELL_X8 FILLER_71_199 ();
 FILLCELL_X1 FILLER_71_207 ();
 FILLCELL_X8 FILLER_71_221 ();
 FILLCELL_X4 FILLER_71_229 ();
 FILLCELL_X4 FILLER_71_250 ();
 FILLCELL_X2 FILLER_71_254 ();
 FILLCELL_X2 FILLER_71_259 ();
 FILLCELL_X16 FILLER_71_274 ();
 FILLCELL_X4 FILLER_71_290 ();
 FILLCELL_X1 FILLER_71_294 ();
 FILLCELL_X4 FILLER_71_299 ();
 FILLCELL_X2 FILLER_71_303 ();
 FILLCELL_X8 FILLER_71_309 ();
 FILLCELL_X2 FILLER_71_317 ();
 FILLCELL_X1 FILLER_71_319 ();
 FILLCELL_X32 FILLER_71_346 ();
 FILLCELL_X2 FILLER_71_378 ();
 FILLCELL_X2 FILLER_71_389 ();
 FILLCELL_X8 FILLER_71_404 ();
 FILLCELL_X4 FILLER_71_412 ();
 FILLCELL_X2 FILLER_71_416 ();
 FILLCELL_X1 FILLER_71_418 ();
 FILLCELL_X16 FILLER_71_433 ();
 FILLCELL_X2 FILLER_71_449 ();
 FILLCELL_X16 FILLER_71_463 ();
 FILLCELL_X1 FILLER_71_479 ();
 FILLCELL_X32 FILLER_71_490 ();
 FILLCELL_X8 FILLER_71_522 ();
 FILLCELL_X4 FILLER_71_530 ();
 FILLCELL_X2 FILLER_71_534 ();
endmodule
